LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY encoderN128 IS
PORT( 
	in1                               :   IN    std_logic;
	in2                               :   IN    std_logic;
	in3                               :   IN    std_logic;
	in4                               :   IN    std_logic;
	in5                               :   IN    std_logic;
	in6                               :   IN    std_logic;
	in7                               :   IN    std_logic;
	in8                               :   IN    std_logic;
	in9                               :   IN    std_logic;
	in10                               :   IN    std_logic;
	in11                               :   IN    std_logic;
	in12                               :   IN    std_logic;
	in13                               :   IN    std_logic;
	in14                               :   IN    std_logic;
	in15                               :   IN    std_logic;
	in16                               :   IN    std_logic;
	in17                               :   IN    std_logic;
	in18                               :   IN    std_logic;
	in19                               :   IN    std_logic;
	in20                               :   IN    std_logic;
	in21                               :   IN    std_logic;
	in22                               :   IN    std_logic;
	in23                               :   IN    std_logic;
	in24                               :   IN    std_logic;
	in25                               :   IN    std_logic;
	in26                               :   IN    std_logic;
	in27                               :   IN    std_logic;
	in28                               :   IN    std_logic;
	in29                               :   IN    std_logic;
	in30                               :   IN    std_logic;
	in31                               :   IN    std_logic;
	in32                               :   IN    std_logic;
	in33                               :   IN    std_logic;
	in34                               :   IN    std_logic;
	in35                               :   IN    std_logic;
	in36                               :   IN    std_logic;
	in37                               :   IN    std_logic;
	in38                               :   IN    std_logic;
	in39                               :   IN    std_logic;
	in40                               :   IN    std_logic;
	in41                               :   IN    std_logic;
	in42                               :   IN    std_logic;
	in43                               :   IN    std_logic;
	in44                               :   IN    std_logic;
	in45                               :   IN    std_logic;
	in46                               :   IN    std_logic;
	in47                               :   IN    std_logic;
	in48                               :   IN    std_logic;
	in49                               :   IN    std_logic;
	in50                               :   IN    std_logic;
	in51                               :   IN    std_logic;
	in52                               :   IN    std_logic;
	in53                               :   IN    std_logic;
	in54                               :   IN    std_logic;
	in55                               :   IN    std_logic;
	in56                               :   IN    std_logic;
	in57                               :   IN    std_logic;
	in58                               :   IN    std_logic;
	in59                               :   IN    std_logic;
	in60                               :   IN    std_logic;
	in61                               :   IN    std_logic;
	in62                               :   IN    std_logic;
	in63                               :   IN    std_logic;
	in64                               :   IN    std_logic;
	in65                               :   IN    std_logic;
	in66                               :   IN    std_logic;
	in67                               :   IN    std_logic;
	in68                               :   IN    std_logic;
	in69                               :   IN    std_logic;
	in70                               :   IN    std_logic;
	in71                               :   IN    std_logic;
	in72                               :   IN    std_logic;
	in73                               :   IN    std_logic;
	in74                               :   IN    std_logic;
	in75                               :   IN    std_logic;
	in76                               :   IN    std_logic;
	in77                               :   IN    std_logic;
	in78                               :   IN    std_logic;
	in79                               :   IN    std_logic;
	in80                               :   IN    std_logic;
	in81                               :   IN    std_logic;
	in82                               :   IN    std_logic;
	in83                               :   IN    std_logic;
	in84                               :   IN    std_logic;
	in85                               :   IN    std_logic;
	in86                               :   IN    std_logic;
	in87                               :   IN    std_logic;
	in88                               :   IN    std_logic;
	in89                               :   IN    std_logic;
	in90                               :   IN    std_logic;
	in91                               :   IN    std_logic;
	in92                               :   IN    std_logic;
	in93                               :   IN    std_logic;
	in94                               :   IN    std_logic;
	in95                               :   IN    std_logic;
	in96                               :   IN    std_logic;
	in97                               :   IN    std_logic;
	in98                               :   IN    std_logic;
	in99                               :   IN    std_logic;
	in100                               :   IN    std_logic;
	in101                               :   IN    std_logic;
	in102                               :   IN    std_logic;
	in103                               :   IN    std_logic;
	in104                               :   IN    std_logic;
	in105                               :   IN    std_logic;
	in106                               :   IN    std_logic;
	in107                               :   IN    std_logic;
	in108                               :   IN    std_logic;
	in109                               :   IN    std_logic;
	in110                               :   IN    std_logic;
	in111                               :   IN    std_logic;
	in112                               :   IN    std_logic;
	in113                               :   IN    std_logic;
	in114                               :   IN    std_logic;
	in115                               :   IN    std_logic;
	in116                               :   IN    std_logic;
	in117                               :   IN    std_logic;
	in118                               :   IN    std_logic;
	in119                               :   IN    std_logic;
	in120                               :   IN    std_logic;
	in121                               :   IN    std_logic;
	in122                               :   IN    std_logic;
	in123                               :   IN    std_logic;
	in124                               :   IN    std_logic;
	in125                               :   IN    std_logic;
	in126                               :   IN    std_logic;
	in127                               :   IN    std_logic;
	in128                               :   IN    std_logic;
	out1                               :   OUT    std_logic;
	out2                               :   OUT    std_logic;
	out3                               :   OUT    std_logic;
	out4                               :   OUT    std_logic;
	out5                               :   OUT    std_logic;
	out6                               :   OUT    std_logic;
	out7                               :   OUT    std_logic;
	out8                               :   OUT    std_logic;
	out9                               :   OUT    std_logic;
	out10                               :   OUT    std_logic;
	out11                               :   OUT    std_logic;
	out12                               :   OUT    std_logic;
	out13                               :   OUT    std_logic;
	out14                               :   OUT    std_logic;
	out15                               :   OUT    std_logic;
	out16                               :   OUT    std_logic;
	out17                               :   OUT    std_logic;
	out18                               :   OUT    std_logic;
	out19                               :   OUT    std_logic;
	out20                               :   OUT    std_logic;
	out21                               :   OUT    std_logic;
	out22                               :   OUT    std_logic;
	out23                               :   OUT    std_logic;
	out24                               :   OUT    std_logic;
	out25                               :   OUT    std_logic;
	out26                               :   OUT    std_logic;
	out27                               :   OUT    std_logic;
	out28                               :   OUT    std_logic;
	out29                               :   OUT    std_logic;
	out30                               :   OUT    std_logic;
	out31                               :   OUT    std_logic;
	out32                               :   OUT    std_logic;
	out33                               :   OUT    std_logic;
	out34                               :   OUT    std_logic;
	out35                               :   OUT    std_logic;
	out36                               :   OUT    std_logic;
	out37                               :   OUT    std_logic;
	out38                               :   OUT    std_logic;
	out39                               :   OUT    std_logic;
	out40                               :   OUT    std_logic;
	out41                               :   OUT    std_logic;
	out42                               :   OUT    std_logic;
	out43                               :   OUT    std_logic;
	out44                               :   OUT    std_logic;
	out45                               :   OUT    std_logic;
	out46                               :   OUT    std_logic;
	out47                               :   OUT    std_logic;
	out48                               :   OUT    std_logic;
	out49                               :   OUT    std_logic;
	out50                               :   OUT    std_logic;
	out51                               :   OUT    std_logic;
	out52                               :   OUT    std_logic;
	out53                               :   OUT    std_logic;
	out54                               :   OUT    std_logic;
	out55                               :   OUT    std_logic;
	out56                               :   OUT    std_logic;
	out57                               :   OUT    std_logic;
	out58                               :   OUT    std_logic;
	out59                               :   OUT    std_logic;
	out60                               :   OUT    std_logic;
	out61                               :   OUT    std_logic;
	out62                               :   OUT    std_logic;
	out63                               :   OUT    std_logic;
	out64                               :   OUT    std_logic;
	out65                               :   OUT    std_logic;
	out66                               :   OUT    std_logic;
	out67                               :   OUT    std_logic;
	out68                               :   OUT    std_logic;
	out69                               :   OUT    std_logic;
	out70                               :   OUT    std_logic;
	out71                               :   OUT    std_logic;
	out72                               :   OUT    std_logic;
	out73                               :   OUT    std_logic;
	out74                               :   OUT    std_logic;
	out75                               :   OUT    std_logic;
	out76                               :   OUT    std_logic;
	out77                               :   OUT    std_logic;
	out78                               :   OUT    std_logic;
	out79                               :   OUT    std_logic;
	out80                               :   OUT    std_logic;
	out81                               :   OUT    std_logic;
	out82                               :   OUT    std_logic;
	out83                               :   OUT    std_logic;
	out84                               :   OUT    std_logic;
	out85                               :   OUT    std_logic;
	out86                               :   OUT    std_logic;
	out87                               :   OUT    std_logic;
	out88                               :   OUT    std_logic;
	out89                               :   OUT    std_logic;
	out90                               :   OUT    std_logic;
	out91                               :   OUT    std_logic;
	out92                               :   OUT    std_logic;
	out93                               :   OUT    std_logic;
	out94                               :   OUT    std_logic;
	out95                               :   OUT    std_logic;
	out96                               :   OUT    std_logic;
	out97                               :   OUT    std_logic;
	out98                               :   OUT    std_logic;
	out99                               :   OUT    std_logic;
	out100                               :   OUT    std_logic;
	out101                               :   OUT    std_logic;
	out102                               :   OUT    std_logic;
	out103                               :   OUT    std_logic;
	out104                               :   OUT    std_logic;
	out105                               :   OUT    std_logic;
	out106                               :   OUT    std_logic;
	out107                               :   OUT    std_logic;
	out108                               :   OUT    std_logic;
	out109                               :   OUT    std_logic;
	out110                               :   OUT    std_logic;
	out111                               :   OUT    std_logic;
	out112                               :   OUT    std_logic;
	out113                               :   OUT    std_logic;
	out114                               :   OUT    std_logic;
	out115                               :   OUT    std_logic;
	out116                               :   OUT    std_logic;
	out117                               :   OUT    std_logic;
	out118                               :   OUT    std_logic;
	out119                               :   OUT    std_logic;
	out120                               :   OUT    std_logic;
	out121                               :   OUT    std_logic;
	out122                               :   OUT    std_logic;
	out123                               :   OUT    std_logic;
	out124                               :   OUT    std_logic;
	out125                               :   OUT    std_logic;
	out126                               :   OUT    std_logic;
	out127                               :   OUT    std_logic;
	out128                               :   OUT    std_logic
	);
END encoderN128;

ARCHITECTURE rtl OF encoderN128 IS

  SIGNAL Logical_Operator_out1_out1            : std_logic;
  SIGNAL Logical_Operator_out2_out1            : std_logic;
  SIGNAL Logical_Operator_out3_out1            : std_logic;
  SIGNAL Logical_Operator_out4_out1            : std_logic;
  SIGNAL Logical_Operator_out5_out1            : std_logic;
  SIGNAL Logical_Operator_out6_out1            : std_logic;
  SIGNAL Logical_Operator_out7_out1            : std_logic;
  SIGNAL Logical_Operator_out8_out1            : std_logic;
  SIGNAL Logical_Operator_out9_out1            : std_logic;
  SIGNAL Logical_Operator_out10_out1            : std_logic;
  SIGNAL Logical_Operator_out11_out1            : std_logic;
  SIGNAL Logical_Operator_out12_out1            : std_logic;
  SIGNAL Logical_Operator_out13_out1            : std_logic;
  SIGNAL Logical_Operator_out14_out1            : std_logic;
  SIGNAL Logical_Operator_out15_out1            : std_logic;
  SIGNAL Logical_Operator_out16_out1            : std_logic;
  SIGNAL Logical_Operator_out17_out1            : std_logic;
  SIGNAL Logical_Operator_out18_out1            : std_logic;
  SIGNAL Logical_Operator_out19_out1            : std_logic;
  SIGNAL Logical_Operator_out20_out1            : std_logic;
  SIGNAL Logical_Operator_out21_out1            : std_logic;
  SIGNAL Logical_Operator_out22_out1            : std_logic;
  SIGNAL Logical_Operator_out23_out1            : std_logic;
  SIGNAL Logical_Operator_out24_out1            : std_logic;
  SIGNAL Logical_Operator_out25_out1            : std_logic;
  SIGNAL Logical_Operator_out26_out1            : std_logic;
  SIGNAL Logical_Operator_out27_out1            : std_logic;
  SIGNAL Logical_Operator_out28_out1            : std_logic;
  SIGNAL Logical_Operator_out29_out1            : std_logic;
  SIGNAL Logical_Operator_out30_out1            : std_logic;
  SIGNAL Logical_Operator_out31_out1            : std_logic;
  SIGNAL Logical_Operator_out32_out1            : std_logic;
  SIGNAL Logical_Operator_out33_out1            : std_logic;
  SIGNAL Logical_Operator_out34_out1            : std_logic;
  SIGNAL Logical_Operator_out35_out1            : std_logic;
  SIGNAL Logical_Operator_out36_out1            : std_logic;
  SIGNAL Logical_Operator_out37_out1            : std_logic;
  SIGNAL Logical_Operator_out38_out1            : std_logic;
  SIGNAL Logical_Operator_out39_out1            : std_logic;
  SIGNAL Logical_Operator_out40_out1            : std_logic;
  SIGNAL Logical_Operator_out41_out1            : std_logic;
  SIGNAL Logical_Operator_out42_out1            : std_logic;
  SIGNAL Logical_Operator_out43_out1            : std_logic;
  SIGNAL Logical_Operator_out44_out1            : std_logic;
  SIGNAL Logical_Operator_out45_out1            : std_logic;
  SIGNAL Logical_Operator_out46_out1            : std_logic;
  SIGNAL Logical_Operator_out47_out1            : std_logic;
  SIGNAL Logical_Operator_out48_out1            : std_logic;
  SIGNAL Logical_Operator_out49_out1            : std_logic;
  SIGNAL Logical_Operator_out50_out1            : std_logic;
  SIGNAL Logical_Operator_out51_out1            : std_logic;
  SIGNAL Logical_Operator_out52_out1            : std_logic;
  SIGNAL Logical_Operator_out53_out1            : std_logic;
  SIGNAL Logical_Operator_out54_out1            : std_logic;
  SIGNAL Logical_Operator_out55_out1            : std_logic;
  SIGNAL Logical_Operator_out56_out1            : std_logic;
  SIGNAL Logical_Operator_out57_out1            : std_logic;
  SIGNAL Logical_Operator_out58_out1            : std_logic;
  SIGNAL Logical_Operator_out59_out1            : std_logic;
  SIGNAL Logical_Operator_out60_out1            : std_logic;
  SIGNAL Logical_Operator_out61_out1            : std_logic;
  SIGNAL Logical_Operator_out62_out1            : std_logic;
  SIGNAL Logical_Operator_out63_out1            : std_logic;
  SIGNAL Logical_Operator_out64_out1            : std_logic;
  SIGNAL Logical_Operator_out65_out1            : std_logic;
  SIGNAL Logical_Operator_out66_out1            : std_logic;
  SIGNAL Logical_Operator_out67_out1            : std_logic;
  SIGNAL Logical_Operator_out68_out1            : std_logic;
  SIGNAL Logical_Operator_out69_out1            : std_logic;
  SIGNAL Logical_Operator_out70_out1            : std_logic;
  SIGNAL Logical_Operator_out71_out1            : std_logic;
  SIGNAL Logical_Operator_out72_out1            : std_logic;
  SIGNAL Logical_Operator_out73_out1            : std_logic;
  SIGNAL Logical_Operator_out74_out1            : std_logic;
  SIGNAL Logical_Operator_out75_out1            : std_logic;
  SIGNAL Logical_Operator_out76_out1            : std_logic;
  SIGNAL Logical_Operator_out77_out1            : std_logic;
  SIGNAL Logical_Operator_out78_out1            : std_logic;
  SIGNAL Logical_Operator_out79_out1            : std_logic;
  SIGNAL Logical_Operator_out80_out1            : std_logic;
  SIGNAL Logical_Operator_out81_out1            : std_logic;
  SIGNAL Logical_Operator_out82_out1            : std_logic;
  SIGNAL Logical_Operator_out83_out1            : std_logic;
  SIGNAL Logical_Operator_out84_out1            : std_logic;
  SIGNAL Logical_Operator_out85_out1            : std_logic;
  SIGNAL Logical_Operator_out86_out1            : std_logic;
  SIGNAL Logical_Operator_out87_out1            : std_logic;
  SIGNAL Logical_Operator_out88_out1            : std_logic;
  SIGNAL Logical_Operator_out89_out1            : std_logic;
  SIGNAL Logical_Operator_out90_out1            : std_logic;
  SIGNAL Logical_Operator_out91_out1            : std_logic;
  SIGNAL Logical_Operator_out92_out1            : std_logic;
  SIGNAL Logical_Operator_out93_out1            : std_logic;
  SIGNAL Logical_Operator_out94_out1            : std_logic;
  SIGNAL Logical_Operator_out95_out1            : std_logic;
  SIGNAL Logical_Operator_out96_out1            : std_logic;
  SIGNAL Logical_Operator_out97_out1            : std_logic;
  SIGNAL Logical_Operator_out98_out1            : std_logic;
  SIGNAL Logical_Operator_out99_out1            : std_logic;
  SIGNAL Logical_Operator_out100_out1            : std_logic;
  SIGNAL Logical_Operator_out101_out1            : std_logic;
  SIGNAL Logical_Operator_out102_out1            : std_logic;
  SIGNAL Logical_Operator_out103_out1            : std_logic;
  SIGNAL Logical_Operator_out104_out1            : std_logic;
  SIGNAL Logical_Operator_out105_out1            : std_logic;
  SIGNAL Logical_Operator_out106_out1            : std_logic;
  SIGNAL Logical_Operator_out107_out1            : std_logic;
  SIGNAL Logical_Operator_out108_out1            : std_logic;
  SIGNAL Logical_Operator_out109_out1            : std_logic;
  SIGNAL Logical_Operator_out110_out1            : std_logic;
  SIGNAL Logical_Operator_out111_out1            : std_logic;
  SIGNAL Logical_Operator_out112_out1            : std_logic;
  SIGNAL Logical_Operator_out113_out1            : std_logic;
  SIGNAL Logical_Operator_out114_out1            : std_logic;
  SIGNAL Logical_Operator_out115_out1            : std_logic;
  SIGNAL Logical_Operator_out116_out1            : std_logic;
  SIGNAL Logical_Operator_out117_out1            : std_logic;
  SIGNAL Logical_Operator_out118_out1            : std_logic;
  SIGNAL Logical_Operator_out119_out1            : std_logic;
  SIGNAL Logical_Operator_out120_out1            : std_logic;
  SIGNAL Logical_Operator_out121_out1            : std_logic;
  SIGNAL Logical_Operator_out122_out1            : std_logic;
  SIGNAL Logical_Operator_out123_out1            : std_logic;
  SIGNAL Logical_Operator_out124_out1            : std_logic;
  SIGNAL Logical_Operator_out125_out1            : std_logic;
  SIGNAL Logical_Operator_out126_out1            : std_logic;
  SIGNAL Logical_Operator_out127_out1            : std_logic;
  SIGNAL Logical_Operator_out128_out1            : std_logic;
  SIGNAL Logical_Operator_out129_out1            : std_logic;
  SIGNAL Logical_Operator_out130_out1            : std_logic;
  SIGNAL Logical_Operator_out131_out1            : std_logic;
  SIGNAL Logical_Operator_out132_out1            : std_logic;
  SIGNAL Logical_Operator_out133_out1            : std_logic;
  SIGNAL Logical_Operator_out134_out1            : std_logic;
  SIGNAL Logical_Operator_out135_out1            : std_logic;
  SIGNAL Logical_Operator_out136_out1            : std_logic;
  SIGNAL Logical_Operator_out137_out1            : std_logic;
  SIGNAL Logical_Operator_out138_out1            : std_logic;
  SIGNAL Logical_Operator_out139_out1            : std_logic;
  SIGNAL Logical_Operator_out140_out1            : std_logic;
  SIGNAL Logical_Operator_out141_out1            : std_logic;
  SIGNAL Logical_Operator_out142_out1            : std_logic;
  SIGNAL Logical_Operator_out143_out1            : std_logic;
  SIGNAL Logical_Operator_out144_out1            : std_logic;
  SIGNAL Logical_Operator_out145_out1            : std_logic;
  SIGNAL Logical_Operator_out146_out1            : std_logic;
  SIGNAL Logical_Operator_out147_out1            : std_logic;
  SIGNAL Logical_Operator_out148_out1            : std_logic;
  SIGNAL Logical_Operator_out149_out1            : std_logic;
  SIGNAL Logical_Operator_out150_out1            : std_logic;
  SIGNAL Logical_Operator_out151_out1            : std_logic;
  SIGNAL Logical_Operator_out152_out1            : std_logic;
  SIGNAL Logical_Operator_out153_out1            : std_logic;
  SIGNAL Logical_Operator_out154_out1            : std_logic;
  SIGNAL Logical_Operator_out155_out1            : std_logic;
  SIGNAL Logical_Operator_out156_out1            : std_logic;
  SIGNAL Logical_Operator_out157_out1            : std_logic;
  SIGNAL Logical_Operator_out158_out1            : std_logic;
  SIGNAL Logical_Operator_out159_out1            : std_logic;
  SIGNAL Logical_Operator_out160_out1            : std_logic;
  SIGNAL Logical_Operator_out161_out1            : std_logic;
  SIGNAL Logical_Operator_out162_out1            : std_logic;
  SIGNAL Logical_Operator_out163_out1            : std_logic;
  SIGNAL Logical_Operator_out164_out1            : std_logic;
  SIGNAL Logical_Operator_out165_out1            : std_logic;
  SIGNAL Logical_Operator_out166_out1            : std_logic;
  SIGNAL Logical_Operator_out167_out1            : std_logic;
  SIGNAL Logical_Operator_out168_out1            : std_logic;
  SIGNAL Logical_Operator_out169_out1            : std_logic;
  SIGNAL Logical_Operator_out170_out1            : std_logic;
  SIGNAL Logical_Operator_out171_out1            : std_logic;
  SIGNAL Logical_Operator_out172_out1            : std_logic;
  SIGNAL Logical_Operator_out173_out1            : std_logic;
  SIGNAL Logical_Operator_out174_out1            : std_logic;
  SIGNAL Logical_Operator_out175_out1            : std_logic;
  SIGNAL Logical_Operator_out176_out1            : std_logic;
  SIGNAL Logical_Operator_out177_out1            : std_logic;
  SIGNAL Logical_Operator_out178_out1            : std_logic;
  SIGNAL Logical_Operator_out179_out1            : std_logic;
  SIGNAL Logical_Operator_out180_out1            : std_logic;
  SIGNAL Logical_Operator_out181_out1            : std_logic;
  SIGNAL Logical_Operator_out182_out1            : std_logic;
  SIGNAL Logical_Operator_out183_out1            : std_logic;
  SIGNAL Logical_Operator_out184_out1            : std_logic;
  SIGNAL Logical_Operator_out185_out1            : std_logic;
  SIGNAL Logical_Operator_out186_out1            : std_logic;
  SIGNAL Logical_Operator_out187_out1            : std_logic;
  SIGNAL Logical_Operator_out188_out1            : std_logic;
  SIGNAL Logical_Operator_out189_out1            : std_logic;
  SIGNAL Logical_Operator_out190_out1            : std_logic;
  SIGNAL Logical_Operator_out191_out1            : std_logic;
  SIGNAL Logical_Operator_out192_out1            : std_logic;
  SIGNAL Logical_Operator_out193_out1            : std_logic;
  SIGNAL Logical_Operator_out194_out1            : std_logic;
  SIGNAL Logical_Operator_out195_out1            : std_logic;
  SIGNAL Logical_Operator_out196_out1            : std_logic;
  SIGNAL Logical_Operator_out197_out1            : std_logic;
  SIGNAL Logical_Operator_out198_out1            : std_logic;
  SIGNAL Logical_Operator_out199_out1            : std_logic;
  SIGNAL Logical_Operator_out200_out1            : std_logic;
  SIGNAL Logical_Operator_out201_out1            : std_logic;
  SIGNAL Logical_Operator_out202_out1            : std_logic;
  SIGNAL Logical_Operator_out203_out1            : std_logic;
  SIGNAL Logical_Operator_out204_out1            : std_logic;
  SIGNAL Logical_Operator_out205_out1            : std_logic;
  SIGNAL Logical_Operator_out206_out1            : std_logic;
  SIGNAL Logical_Operator_out207_out1            : std_logic;
  SIGNAL Logical_Operator_out208_out1            : std_logic;
  SIGNAL Logical_Operator_out209_out1            : std_logic;
  SIGNAL Logical_Operator_out210_out1            : std_logic;
  SIGNAL Logical_Operator_out211_out1            : std_logic;
  SIGNAL Logical_Operator_out212_out1            : std_logic;
  SIGNAL Logical_Operator_out213_out1            : std_logic;
  SIGNAL Logical_Operator_out214_out1            : std_logic;
  SIGNAL Logical_Operator_out215_out1            : std_logic;
  SIGNAL Logical_Operator_out216_out1            : std_logic;
  SIGNAL Logical_Operator_out217_out1            : std_logic;
  SIGNAL Logical_Operator_out218_out1            : std_logic;
  SIGNAL Logical_Operator_out219_out1            : std_logic;
  SIGNAL Logical_Operator_out220_out1            : std_logic;
  SIGNAL Logical_Operator_out221_out1            : std_logic;
  SIGNAL Logical_Operator_out222_out1            : std_logic;
  SIGNAL Logical_Operator_out223_out1            : std_logic;
  SIGNAL Logical_Operator_out224_out1            : std_logic;
  SIGNAL Logical_Operator_out225_out1            : std_logic;
  SIGNAL Logical_Operator_out226_out1            : std_logic;
  SIGNAL Logical_Operator_out227_out1            : std_logic;
  SIGNAL Logical_Operator_out228_out1            : std_logic;
  SIGNAL Logical_Operator_out229_out1            : std_logic;
  SIGNAL Logical_Operator_out230_out1            : std_logic;
  SIGNAL Logical_Operator_out231_out1            : std_logic;
  SIGNAL Logical_Operator_out232_out1            : std_logic;
  SIGNAL Logical_Operator_out233_out1            : std_logic;
  SIGNAL Logical_Operator_out234_out1            : std_logic;
  SIGNAL Logical_Operator_out235_out1            : std_logic;
  SIGNAL Logical_Operator_out236_out1            : std_logic;
  SIGNAL Logical_Operator_out237_out1            : std_logic;
  SIGNAL Logical_Operator_out238_out1            : std_logic;
  SIGNAL Logical_Operator_out239_out1            : std_logic;
  SIGNAL Logical_Operator_out240_out1            : std_logic;
  SIGNAL Logical_Operator_out241_out1            : std_logic;
  SIGNAL Logical_Operator_out242_out1            : std_logic;
  SIGNAL Logical_Operator_out243_out1            : std_logic;
  SIGNAL Logical_Operator_out244_out1            : std_logic;
  SIGNAL Logical_Operator_out245_out1            : std_logic;
  SIGNAL Logical_Operator_out246_out1            : std_logic;
  SIGNAL Logical_Operator_out247_out1            : std_logic;
  SIGNAL Logical_Operator_out248_out1            : std_logic;
  SIGNAL Logical_Operator_out249_out1            : std_logic;
  SIGNAL Logical_Operator_out250_out1            : std_logic;
  SIGNAL Logical_Operator_out251_out1            : std_logic;
  SIGNAL Logical_Operator_out252_out1            : std_logic;
  SIGNAL Logical_Operator_out253_out1            : std_logic;
  SIGNAL Logical_Operator_out254_out1            : std_logic;
  SIGNAL Logical_Operator_out255_out1            : std_logic;
  SIGNAL Logical_Operator_out256_out1            : std_logic;
  SIGNAL Logical_Operator_out257_out1            : std_logic;
  SIGNAL Logical_Operator_out258_out1            : std_logic;
  SIGNAL Logical_Operator_out259_out1            : std_logic;
  SIGNAL Logical_Operator_out260_out1            : std_logic;
  SIGNAL Logical_Operator_out261_out1            : std_logic;
  SIGNAL Logical_Operator_out262_out1            : std_logic;
  SIGNAL Logical_Operator_out263_out1            : std_logic;
  SIGNAL Logical_Operator_out264_out1            : std_logic;
  SIGNAL Logical_Operator_out265_out1            : std_logic;
  SIGNAL Logical_Operator_out266_out1            : std_logic;
  SIGNAL Logical_Operator_out267_out1            : std_logic;
  SIGNAL Logical_Operator_out268_out1            : std_logic;
  SIGNAL Logical_Operator_out269_out1            : std_logic;
  SIGNAL Logical_Operator_out270_out1            : std_logic;
  SIGNAL Logical_Operator_out271_out1            : std_logic;
  SIGNAL Logical_Operator_out272_out1            : std_logic;
  SIGNAL Logical_Operator_out273_out1            : std_logic;
  SIGNAL Logical_Operator_out274_out1            : std_logic;
  SIGNAL Logical_Operator_out275_out1            : std_logic;
  SIGNAL Logical_Operator_out276_out1            : std_logic;
  SIGNAL Logical_Operator_out277_out1            : std_logic;
  SIGNAL Logical_Operator_out278_out1            : std_logic;
  SIGNAL Logical_Operator_out279_out1            : std_logic;
  SIGNAL Logical_Operator_out280_out1            : std_logic;
  SIGNAL Logical_Operator_out281_out1            : std_logic;
  SIGNAL Logical_Operator_out282_out1            : std_logic;
  SIGNAL Logical_Operator_out283_out1            : std_logic;
  SIGNAL Logical_Operator_out284_out1            : std_logic;
  SIGNAL Logical_Operator_out285_out1            : std_logic;
  SIGNAL Logical_Operator_out286_out1            : std_logic;
  SIGNAL Logical_Operator_out287_out1            : std_logic;
  SIGNAL Logical_Operator_out288_out1            : std_logic;
  SIGNAL Logical_Operator_out289_out1            : std_logic;
  SIGNAL Logical_Operator_out290_out1            : std_logic;
  SIGNAL Logical_Operator_out291_out1            : std_logic;
  SIGNAL Logical_Operator_out292_out1            : std_logic;
  SIGNAL Logical_Operator_out293_out1            : std_logic;
  SIGNAL Logical_Operator_out294_out1            : std_logic;
  SIGNAL Logical_Operator_out295_out1            : std_logic;
  SIGNAL Logical_Operator_out296_out1            : std_logic;
  SIGNAL Logical_Operator_out297_out1            : std_logic;
  SIGNAL Logical_Operator_out298_out1            : std_logic;
  SIGNAL Logical_Operator_out299_out1            : std_logic;
  SIGNAL Logical_Operator_out300_out1            : std_logic;
  SIGNAL Logical_Operator_out301_out1            : std_logic;
  SIGNAL Logical_Operator_out302_out1            : std_logic;
  SIGNAL Logical_Operator_out303_out1            : std_logic;
  SIGNAL Logical_Operator_out304_out1            : std_logic;
  SIGNAL Logical_Operator_out305_out1            : std_logic;
  SIGNAL Logical_Operator_out306_out1            : std_logic;
  SIGNAL Logical_Operator_out307_out1            : std_logic;
  SIGNAL Logical_Operator_out308_out1            : std_logic;
  SIGNAL Logical_Operator_out309_out1            : std_logic;
  SIGNAL Logical_Operator_out310_out1            : std_logic;
  SIGNAL Logical_Operator_out311_out1            : std_logic;
  SIGNAL Logical_Operator_out312_out1            : std_logic;
  SIGNAL Logical_Operator_out313_out1            : std_logic;
  SIGNAL Logical_Operator_out314_out1            : std_logic;
  SIGNAL Logical_Operator_out315_out1            : std_logic;
  SIGNAL Logical_Operator_out316_out1            : std_logic;
  SIGNAL Logical_Operator_out317_out1            : std_logic;
  SIGNAL Logical_Operator_out318_out1            : std_logic;
  SIGNAL Logical_Operator_out319_out1            : std_logic;
  SIGNAL Logical_Operator_out320_out1            : std_logic;
  SIGNAL Logical_Operator_out321_out1            : std_logic;
  SIGNAL Logical_Operator_out322_out1            : std_logic;
  SIGNAL Logical_Operator_out323_out1            : std_logic;
  SIGNAL Logical_Operator_out324_out1            : std_logic;
  SIGNAL Logical_Operator_out325_out1            : std_logic;
  SIGNAL Logical_Operator_out326_out1            : std_logic;
  SIGNAL Logical_Operator_out327_out1            : std_logic;
  SIGNAL Logical_Operator_out328_out1            : std_logic;
  SIGNAL Logical_Operator_out329_out1            : std_logic;
  SIGNAL Logical_Operator_out330_out1            : std_logic;
  SIGNAL Logical_Operator_out331_out1            : std_logic;
  SIGNAL Logical_Operator_out332_out1            : std_logic;
  SIGNAL Logical_Operator_out333_out1            : std_logic;
  SIGNAL Logical_Operator_out334_out1            : std_logic;
  SIGNAL Logical_Operator_out335_out1            : std_logic;
  SIGNAL Logical_Operator_out336_out1            : std_logic;
  SIGNAL Logical_Operator_out337_out1            : std_logic;
  SIGNAL Logical_Operator_out338_out1            : std_logic;
  SIGNAL Logical_Operator_out339_out1            : std_logic;
  SIGNAL Logical_Operator_out340_out1            : std_logic;
  SIGNAL Logical_Operator_out341_out1            : std_logic;
  SIGNAL Logical_Operator_out342_out1            : std_logic;
  SIGNAL Logical_Operator_out343_out1            : std_logic;
  SIGNAL Logical_Operator_out344_out1            : std_logic;
  SIGNAL Logical_Operator_out345_out1            : std_logic;
  SIGNAL Logical_Operator_out346_out1            : std_logic;
  SIGNAL Logical_Operator_out347_out1            : std_logic;
  SIGNAL Logical_Operator_out348_out1            : std_logic;
  SIGNAL Logical_Operator_out349_out1            : std_logic;
  SIGNAL Logical_Operator_out350_out1            : std_logic;
  SIGNAL Logical_Operator_out351_out1            : std_logic;
  SIGNAL Logical_Operator_out352_out1            : std_logic;
  SIGNAL Logical_Operator_out353_out1            : std_logic;
  SIGNAL Logical_Operator_out354_out1            : std_logic;
  SIGNAL Logical_Operator_out355_out1            : std_logic;
  SIGNAL Logical_Operator_out356_out1            : std_logic;
  SIGNAL Logical_Operator_out357_out1            : std_logic;
  SIGNAL Logical_Operator_out358_out1            : std_logic;
  SIGNAL Logical_Operator_out359_out1            : std_logic;
  SIGNAL Logical_Operator_out360_out1            : std_logic;
  SIGNAL Logical_Operator_out361_out1            : std_logic;
  SIGNAL Logical_Operator_out362_out1            : std_logic;
  SIGNAL Logical_Operator_out363_out1            : std_logic;
  SIGNAL Logical_Operator_out364_out1            : std_logic;
  SIGNAL Logical_Operator_out365_out1            : std_logic;
  SIGNAL Logical_Operator_out366_out1            : std_logic;
  SIGNAL Logical_Operator_out367_out1            : std_logic;
  SIGNAL Logical_Operator_out368_out1            : std_logic;
  SIGNAL Logical_Operator_out369_out1            : std_logic;
  SIGNAL Logical_Operator_out370_out1            : std_logic;
  SIGNAL Logical_Operator_out371_out1            : std_logic;
  SIGNAL Logical_Operator_out372_out1            : std_logic;
  SIGNAL Logical_Operator_out373_out1            : std_logic;
  SIGNAL Logical_Operator_out374_out1            : std_logic;
  SIGNAL Logical_Operator_out375_out1            : std_logic;
  SIGNAL Logical_Operator_out376_out1            : std_logic;
  SIGNAL Logical_Operator_out377_out1            : std_logic;
  SIGNAL Logical_Operator_out378_out1            : std_logic;
  SIGNAL Logical_Operator_out379_out1            : std_logic;
  SIGNAL Logical_Operator_out380_out1            : std_logic;
  SIGNAL Logical_Operator_out381_out1            : std_logic;
  SIGNAL Logical_Operator_out382_out1            : std_logic;
  SIGNAL Logical_Operator_out383_out1            : std_logic;
  SIGNAL Logical_Operator_out384_out1            : std_logic;
  SIGNAL Logical_Operator_out385_out1            : std_logic;
  SIGNAL Logical_Operator_out386_out1            : std_logic;
  SIGNAL Logical_Operator_out387_out1            : std_logic;
  SIGNAL Logical_Operator_out388_out1            : std_logic;
  SIGNAL Logical_Operator_out389_out1            : std_logic;
  SIGNAL Logical_Operator_out390_out1            : std_logic;
  SIGNAL Logical_Operator_out391_out1            : std_logic;
  SIGNAL Logical_Operator_out392_out1            : std_logic;
  SIGNAL Logical_Operator_out393_out1            : std_logic;
  SIGNAL Logical_Operator_out394_out1            : std_logic;
  SIGNAL Logical_Operator_out395_out1            : std_logic;
  SIGNAL Logical_Operator_out396_out1            : std_logic;
  SIGNAL Logical_Operator_out397_out1            : std_logic;
  SIGNAL Logical_Operator_out398_out1            : std_logic;
  SIGNAL Logical_Operator_out399_out1            : std_logic;
  SIGNAL Logical_Operator_out400_out1            : std_logic;
  SIGNAL Logical_Operator_out401_out1            : std_logic;
  SIGNAL Logical_Operator_out402_out1            : std_logic;
  SIGNAL Logical_Operator_out403_out1            : std_logic;
  SIGNAL Logical_Operator_out404_out1            : std_logic;
  SIGNAL Logical_Operator_out405_out1            : std_logic;
  SIGNAL Logical_Operator_out406_out1            : std_logic;
  SIGNAL Logical_Operator_out407_out1            : std_logic;
  SIGNAL Logical_Operator_out408_out1            : std_logic;
  SIGNAL Logical_Operator_out409_out1            : std_logic;
  SIGNAL Logical_Operator_out410_out1            : std_logic;
  SIGNAL Logical_Operator_out411_out1            : std_logic;
  SIGNAL Logical_Operator_out412_out1            : std_logic;
  SIGNAL Logical_Operator_out413_out1            : std_logic;
  SIGNAL Logical_Operator_out414_out1            : std_logic;
  SIGNAL Logical_Operator_out415_out1            : std_logic;
  SIGNAL Logical_Operator_out416_out1            : std_logic;
  SIGNAL Logical_Operator_out417_out1            : std_logic;
  SIGNAL Logical_Operator_out418_out1            : std_logic;
  SIGNAL Logical_Operator_out419_out1            : std_logic;
  SIGNAL Logical_Operator_out420_out1            : std_logic;
  SIGNAL Logical_Operator_out421_out1            : std_logic;
  SIGNAL Logical_Operator_out422_out1            : std_logic;
  SIGNAL Logical_Operator_out423_out1            : std_logic;
  SIGNAL Logical_Operator_out424_out1            : std_logic;
  SIGNAL Logical_Operator_out425_out1            : std_logic;
  SIGNAL Logical_Operator_out426_out1            : std_logic;
  SIGNAL Logical_Operator_out427_out1            : std_logic;
  SIGNAL Logical_Operator_out428_out1            : std_logic;
  SIGNAL Logical_Operator_out429_out1            : std_logic;
  SIGNAL Logical_Operator_out430_out1            : std_logic;
  SIGNAL Logical_Operator_out431_out1            : std_logic;
  SIGNAL Logical_Operator_out432_out1            : std_logic;
  SIGNAL Logical_Operator_out433_out1            : std_logic;
  SIGNAL Logical_Operator_out434_out1            : std_logic;
  SIGNAL Logical_Operator_out435_out1            : std_logic;
  SIGNAL Logical_Operator_out436_out1            : std_logic;
  SIGNAL Logical_Operator_out437_out1            : std_logic;
  SIGNAL Logical_Operator_out438_out1            : std_logic;
  SIGNAL Logical_Operator_out439_out1            : std_logic;
  SIGNAL Logical_Operator_out440_out1            : std_logic;
  SIGNAL Logical_Operator_out441_out1            : std_logic;
  SIGNAL Logical_Operator_out442_out1            : std_logic;
  SIGNAL Logical_Operator_out443_out1            : std_logic;
  SIGNAL Logical_Operator_out444_out1            : std_logic;
  SIGNAL Logical_Operator_out445_out1            : std_logic;
  SIGNAL Logical_Operator_out446_out1            : std_logic;
  SIGNAL Logical_Operator_out447_out1            : std_logic;
  SIGNAL Logical_Operator_out448_out1            : std_logic;

BEGIN

  Logical_Operator_out1_out1 <= in1 XOR in2;

  Logical_Operator_out2_out1 <= in3 XOR in4;

  Logical_Operator_out3_out1 <= in5 XOR in6;

  Logical_Operator_out4_out1 <= in7 XOR in8;

  Logical_Operator_out5_out1 <= in9 XOR in10;

  Logical_Operator_out6_out1 <= in11 XOR in12;

  Logical_Operator_out7_out1 <= in13 XOR in14;

  Logical_Operator_out8_out1 <= in15 XOR in16;

  Logical_Operator_out9_out1 <= in17 XOR in18;

  Logical_Operator_out10_out1 <= in19 XOR in20;

  Logical_Operator_out11_out1 <= in21 XOR in22;

  Logical_Operator_out12_out1 <= in23 XOR in24;

  Logical_Operator_out13_out1 <= in25 XOR in26;

  Logical_Operator_out14_out1 <= in27 XOR in28;

  Logical_Operator_out15_out1 <= in29 XOR in30;

  Logical_Operator_out16_out1 <= in31 XOR in32;

  Logical_Operator_out17_out1 <= in33 XOR in34;

  Logical_Operator_out18_out1 <= in35 XOR in36;

  Logical_Operator_out19_out1 <= in37 XOR in38;

  Logical_Operator_out20_out1 <= in39 XOR in40;

  Logical_Operator_out21_out1 <= in41 XOR in42;

  Logical_Operator_out22_out1 <= in43 XOR in44;

  Logical_Operator_out23_out1 <= in45 XOR in46;

  Logical_Operator_out24_out1 <= in47 XOR in48;

  Logical_Operator_out25_out1 <= in49 XOR in50;

  Logical_Operator_out26_out1 <= in51 XOR in52;

  Logical_Operator_out27_out1 <= in53 XOR in54;

  Logical_Operator_out28_out1 <= in55 XOR in56;

  Logical_Operator_out29_out1 <= in57 XOR in58;

  Logical_Operator_out30_out1 <= in59 XOR in60;

  Logical_Operator_out31_out1 <= in61 XOR in62;

  Logical_Operator_out32_out1 <= in63 XOR in64;

  Logical_Operator_out33_out1 <= in65 XOR in66;

  Logical_Operator_out34_out1 <= in67 XOR in68;

  Logical_Operator_out35_out1 <= in69 XOR in70;

  Logical_Operator_out36_out1 <= in71 XOR in72;

  Logical_Operator_out37_out1 <= in73 XOR in74;

  Logical_Operator_out38_out1 <= in75 XOR in76;

  Logical_Operator_out39_out1 <= in77 XOR in78;

  Logical_Operator_out40_out1 <= in79 XOR in80;

  Logical_Operator_out41_out1 <= in81 XOR in82;

  Logical_Operator_out42_out1 <= in83 XOR in84;

  Logical_Operator_out43_out1 <= in85 XOR in86;

  Logical_Operator_out44_out1 <= in87 XOR in88;

  Logical_Operator_out45_out1 <= in89 XOR in90;

  Logical_Operator_out46_out1 <= in91 XOR in92;

  Logical_Operator_out47_out1 <= in93 XOR in94;

  Logical_Operator_out48_out1 <= in95 XOR in96;

  Logical_Operator_out49_out1 <= in97 XOR in98;

  Logical_Operator_out50_out1 <= in99 XOR in100;

  Logical_Operator_out51_out1 <= in101 XOR in102;

  Logical_Operator_out52_out1 <= in103 XOR in104;

  Logical_Operator_out53_out1 <= in105 XOR in106;

  Logical_Operator_out54_out1 <= in107 XOR in108;

  Logical_Operator_out55_out1 <= in109 XOR in110;

  Logical_Operator_out56_out1 <= in111 XOR in112;

  Logical_Operator_out57_out1 <= in113 XOR in114;

  Logical_Operator_out58_out1 <= in115 XOR in116;

  Logical_Operator_out59_out1 <= in117 XOR in118;

  Logical_Operator_out60_out1 <= in119 XOR in120;

  Logical_Operator_out61_out1 <= in121 XOR in122;

  Logical_Operator_out62_out1 <= in123 XOR in124;

  Logical_Operator_out63_out1 <= in125 XOR in126;

  Logical_Operator_out64_out1 <= in127 XOR in128;

  Logical_Operator_out65_out1 <= Logical_Operator_out1_out1 XOR Logical_Operator_out2_out1;

  Logical_Operator_out66_out1 <= in2 XOR in4;

  Logical_Operator_out67_out1 <= Logical_Operator_out3_out1 XOR Logical_Operator_out4_out1;

  Logical_Operator_out68_out1 <= in6 XOR in8;

  Logical_Operator_out69_out1 <= Logical_Operator_out5_out1 XOR Logical_Operator_out6_out1;

  Logical_Operator_out70_out1 <= in10 XOR in12;

  Logical_Operator_out71_out1 <= Logical_Operator_out7_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out72_out1 <= in14 XOR in16;

  Logical_Operator_out73_out1 <= Logical_Operator_out9_out1 XOR Logical_Operator_out10_out1;

  Logical_Operator_out74_out1 <= in18 XOR in20;

  Logical_Operator_out75_out1 <= Logical_Operator_out11_out1 XOR Logical_Operator_out12_out1;

  Logical_Operator_out76_out1 <= in22 XOR in24;

  Logical_Operator_out77_out1 <= Logical_Operator_out13_out1 XOR Logical_Operator_out14_out1;

  Logical_Operator_out78_out1 <= in26 XOR in28;

  Logical_Operator_out79_out1 <= Logical_Operator_out15_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out80_out1 <= in30 XOR in32;

  Logical_Operator_out81_out1 <= Logical_Operator_out17_out1 XOR Logical_Operator_out18_out1;

  Logical_Operator_out82_out1 <= in34 XOR in36;

  Logical_Operator_out83_out1 <= Logical_Operator_out19_out1 XOR Logical_Operator_out20_out1;

  Logical_Operator_out84_out1 <= in38 XOR in40;

  Logical_Operator_out85_out1 <= Logical_Operator_out21_out1 XOR Logical_Operator_out22_out1;

  Logical_Operator_out86_out1 <= in42 XOR in44;

  Logical_Operator_out87_out1 <= Logical_Operator_out23_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out88_out1 <= in46 XOR in48;

  Logical_Operator_out89_out1 <= Logical_Operator_out25_out1 XOR Logical_Operator_out26_out1;

  Logical_Operator_out90_out1 <= in50 XOR in52;

  Logical_Operator_out91_out1 <= Logical_Operator_out27_out1 XOR Logical_Operator_out28_out1;

  Logical_Operator_out92_out1 <= in54 XOR in56;

  Logical_Operator_out93_out1 <= Logical_Operator_out29_out1 XOR Logical_Operator_out30_out1;

  Logical_Operator_out94_out1 <= in58 XOR in60;

  Logical_Operator_out95_out1 <= Logical_Operator_out31_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out96_out1 <= in62 XOR in64;

  Logical_Operator_out97_out1 <= Logical_Operator_out33_out1 XOR Logical_Operator_out34_out1;

  Logical_Operator_out98_out1 <= in66 XOR in68;

  Logical_Operator_out99_out1 <= Logical_Operator_out35_out1 XOR Logical_Operator_out36_out1;

  Logical_Operator_out100_out1 <= in70 XOR in72;

  Logical_Operator_out101_out1 <= Logical_Operator_out37_out1 XOR Logical_Operator_out38_out1;

  Logical_Operator_out102_out1 <= in74 XOR in76;

  Logical_Operator_out103_out1 <= Logical_Operator_out39_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out104_out1 <= in78 XOR in80;

  Logical_Operator_out105_out1 <= Logical_Operator_out41_out1 XOR Logical_Operator_out42_out1;

  Logical_Operator_out106_out1 <= in82 XOR in84;

  Logical_Operator_out107_out1 <= Logical_Operator_out43_out1 XOR Logical_Operator_out44_out1;

  Logical_Operator_out108_out1 <= in86 XOR in88;

  Logical_Operator_out109_out1 <= Logical_Operator_out45_out1 XOR Logical_Operator_out46_out1;

  Logical_Operator_out110_out1 <= in90 XOR in92;

  Logical_Operator_out111_out1 <= Logical_Operator_out47_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out112_out1 <= in94 XOR in96;

  Logical_Operator_out113_out1 <= Logical_Operator_out49_out1 XOR Logical_Operator_out50_out1;

  Logical_Operator_out114_out1 <= in98 XOR in100;

  Logical_Operator_out115_out1 <= Logical_Operator_out51_out1 XOR Logical_Operator_out52_out1;

  Logical_Operator_out116_out1 <= in102 XOR in104;

  Logical_Operator_out117_out1 <= Logical_Operator_out53_out1 XOR Logical_Operator_out54_out1;

  Logical_Operator_out118_out1 <= in106 XOR in108;

  Logical_Operator_out119_out1 <= Logical_Operator_out55_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out120_out1 <= in110 XOR in112;

  Logical_Operator_out121_out1 <= Logical_Operator_out57_out1 XOR Logical_Operator_out58_out1;

  Logical_Operator_out122_out1 <= in114 XOR in116;

  Logical_Operator_out123_out1 <= Logical_Operator_out59_out1 XOR Logical_Operator_out60_out1;

  Logical_Operator_out124_out1 <= in118 XOR in120;

  Logical_Operator_out125_out1 <= Logical_Operator_out61_out1 XOR Logical_Operator_out62_out1;

  Logical_Operator_out126_out1 <= in122 XOR in124;

  Logical_Operator_out127_out1 <= Logical_Operator_out63_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out128_out1 <= in126 XOR in128;

  Logical_Operator_out129_out1 <= Logical_Operator_out65_out1 XOR Logical_Operator_out67_out1;

  Logical_Operator_out130_out1 <= Logical_Operator_out66_out1 XOR Logical_Operator_out68_out1;

  Logical_Operator_out131_out1 <= Logical_Operator_out2_out1 XOR Logical_Operator_out4_out1;

  Logical_Operator_out132_out1 <= in4 XOR in8;

  Logical_Operator_out133_out1 <= Logical_Operator_out69_out1 XOR Logical_Operator_out71_out1;

  Logical_Operator_out134_out1 <= Logical_Operator_out70_out1 XOR Logical_Operator_out72_out1;

  Logical_Operator_out135_out1 <= Logical_Operator_out6_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out136_out1 <= in12 XOR in16;

  Logical_Operator_out137_out1 <= Logical_Operator_out73_out1 XOR Logical_Operator_out75_out1;

  Logical_Operator_out138_out1 <= Logical_Operator_out74_out1 XOR Logical_Operator_out76_out1;

  Logical_Operator_out139_out1 <= Logical_Operator_out10_out1 XOR Logical_Operator_out12_out1;

  Logical_Operator_out140_out1 <= in20 XOR in24;

  Logical_Operator_out141_out1 <= Logical_Operator_out77_out1 XOR Logical_Operator_out79_out1;

  Logical_Operator_out142_out1 <= Logical_Operator_out78_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out143_out1 <= Logical_Operator_out14_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out144_out1 <= in28 XOR in32;

  Logical_Operator_out145_out1 <= Logical_Operator_out81_out1 XOR Logical_Operator_out83_out1;

  Logical_Operator_out146_out1 <= Logical_Operator_out82_out1 XOR Logical_Operator_out84_out1;

  Logical_Operator_out147_out1 <= Logical_Operator_out18_out1 XOR Logical_Operator_out20_out1;

  Logical_Operator_out148_out1 <= in36 XOR in40;

  Logical_Operator_out149_out1 <= Logical_Operator_out85_out1 XOR Logical_Operator_out87_out1;

  Logical_Operator_out150_out1 <= Logical_Operator_out86_out1 XOR Logical_Operator_out88_out1;

  Logical_Operator_out151_out1 <= Logical_Operator_out22_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out152_out1 <= in44 XOR in48;

  Logical_Operator_out153_out1 <= Logical_Operator_out89_out1 XOR Logical_Operator_out91_out1;

  Logical_Operator_out154_out1 <= Logical_Operator_out90_out1 XOR Logical_Operator_out92_out1;

  Logical_Operator_out155_out1 <= Logical_Operator_out26_out1 XOR Logical_Operator_out28_out1;

  Logical_Operator_out156_out1 <= in52 XOR in56;

  Logical_Operator_out157_out1 <= Logical_Operator_out93_out1 XOR Logical_Operator_out95_out1;

  Logical_Operator_out158_out1 <= Logical_Operator_out94_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out159_out1 <= Logical_Operator_out30_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out160_out1 <= in60 XOR in64;

  Logical_Operator_out161_out1 <= Logical_Operator_out97_out1 XOR Logical_Operator_out99_out1;

  Logical_Operator_out162_out1 <= Logical_Operator_out98_out1 XOR Logical_Operator_out100_out1;

  Logical_Operator_out163_out1 <= Logical_Operator_out34_out1 XOR Logical_Operator_out36_out1;

  Logical_Operator_out164_out1 <= in68 XOR in72;

  Logical_Operator_out165_out1 <= Logical_Operator_out101_out1 XOR Logical_Operator_out103_out1;

  Logical_Operator_out166_out1 <= Logical_Operator_out102_out1 XOR Logical_Operator_out104_out1;

  Logical_Operator_out167_out1 <= Logical_Operator_out38_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out168_out1 <= in76 XOR in80;

  Logical_Operator_out169_out1 <= Logical_Operator_out105_out1 XOR Logical_Operator_out107_out1;

  Logical_Operator_out170_out1 <= Logical_Operator_out106_out1 XOR Logical_Operator_out108_out1;

  Logical_Operator_out171_out1 <= Logical_Operator_out42_out1 XOR Logical_Operator_out44_out1;

  Logical_Operator_out172_out1 <= in84 XOR in88;

  Logical_Operator_out173_out1 <= Logical_Operator_out109_out1 XOR Logical_Operator_out111_out1;

  Logical_Operator_out174_out1 <= Logical_Operator_out110_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out175_out1 <= Logical_Operator_out46_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out176_out1 <= in92 XOR in96;

  Logical_Operator_out177_out1 <= Logical_Operator_out113_out1 XOR Logical_Operator_out115_out1;

  Logical_Operator_out178_out1 <= Logical_Operator_out114_out1 XOR Logical_Operator_out116_out1;

  Logical_Operator_out179_out1 <= Logical_Operator_out50_out1 XOR Logical_Operator_out52_out1;

  Logical_Operator_out180_out1 <= in100 XOR in104;

  Logical_Operator_out181_out1 <= Logical_Operator_out117_out1 XOR Logical_Operator_out119_out1;

  Logical_Operator_out182_out1 <= Logical_Operator_out118_out1 XOR Logical_Operator_out120_out1;

  Logical_Operator_out183_out1 <= Logical_Operator_out54_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out184_out1 <= in108 XOR in112;

  Logical_Operator_out185_out1 <= Logical_Operator_out121_out1 XOR Logical_Operator_out123_out1;

  Logical_Operator_out186_out1 <= Logical_Operator_out122_out1 XOR Logical_Operator_out124_out1;

  Logical_Operator_out187_out1 <= Logical_Operator_out58_out1 XOR Logical_Operator_out60_out1;

  Logical_Operator_out188_out1 <= in116 XOR in120;

  Logical_Operator_out189_out1 <= Logical_Operator_out125_out1 XOR Logical_Operator_out127_out1;

  Logical_Operator_out190_out1 <= Logical_Operator_out126_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out191_out1 <= Logical_Operator_out62_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out192_out1 <= in124 XOR in128;

  Logical_Operator_out193_out1 <= Logical_Operator_out129_out1 XOR Logical_Operator_out133_out1;

  Logical_Operator_out194_out1 <= Logical_Operator_out130_out1 XOR Logical_Operator_out134_out1;

  Logical_Operator_out195_out1 <= Logical_Operator_out131_out1 XOR Logical_Operator_out135_out1;

  Logical_Operator_out196_out1 <= Logical_Operator_out132_out1 XOR Logical_Operator_out136_out1;

  Logical_Operator_out197_out1 <= Logical_Operator_out67_out1 XOR Logical_Operator_out71_out1;

  Logical_Operator_out198_out1 <= Logical_Operator_out68_out1 XOR Logical_Operator_out72_out1;

  Logical_Operator_out199_out1 <= Logical_Operator_out4_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out200_out1 <= in8 XOR in16;

  Logical_Operator_out201_out1 <= Logical_Operator_out137_out1 XOR Logical_Operator_out141_out1;

  Logical_Operator_out202_out1 <= Logical_Operator_out138_out1 XOR Logical_Operator_out142_out1;

  Logical_Operator_out203_out1 <= Logical_Operator_out139_out1 XOR Logical_Operator_out143_out1;

  Logical_Operator_out204_out1 <= Logical_Operator_out140_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out205_out1 <= Logical_Operator_out75_out1 XOR Logical_Operator_out79_out1;

  Logical_Operator_out206_out1 <= Logical_Operator_out76_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out207_out1 <= Logical_Operator_out12_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out208_out1 <= in24 XOR in32;

  Logical_Operator_out209_out1 <= Logical_Operator_out145_out1 XOR Logical_Operator_out149_out1;

  Logical_Operator_out210_out1 <= Logical_Operator_out146_out1 XOR Logical_Operator_out150_out1;

  Logical_Operator_out211_out1 <= Logical_Operator_out147_out1 XOR Logical_Operator_out151_out1;

  Logical_Operator_out212_out1 <= Logical_Operator_out148_out1 XOR Logical_Operator_out152_out1;

  Logical_Operator_out213_out1 <= Logical_Operator_out83_out1 XOR Logical_Operator_out87_out1;

  Logical_Operator_out214_out1 <= Logical_Operator_out84_out1 XOR Logical_Operator_out88_out1;

  Logical_Operator_out215_out1 <= Logical_Operator_out20_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out216_out1 <= in40 XOR in48;

  Logical_Operator_out217_out1 <= Logical_Operator_out153_out1 XOR Logical_Operator_out157_out1;

  Logical_Operator_out218_out1 <= Logical_Operator_out154_out1 XOR Logical_Operator_out158_out1;

  Logical_Operator_out219_out1 <= Logical_Operator_out155_out1 XOR Logical_Operator_out159_out1;

  Logical_Operator_out220_out1 <= Logical_Operator_out156_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out221_out1 <= Logical_Operator_out91_out1 XOR Logical_Operator_out95_out1;

  Logical_Operator_out222_out1 <= Logical_Operator_out92_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out223_out1 <= Logical_Operator_out28_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out224_out1 <= in56 XOR in64;

  Logical_Operator_out225_out1 <= Logical_Operator_out161_out1 XOR Logical_Operator_out165_out1;

  Logical_Operator_out226_out1 <= Logical_Operator_out162_out1 XOR Logical_Operator_out166_out1;

  Logical_Operator_out227_out1 <= Logical_Operator_out163_out1 XOR Logical_Operator_out167_out1;

  Logical_Operator_out228_out1 <= Logical_Operator_out164_out1 XOR Logical_Operator_out168_out1;

  Logical_Operator_out229_out1 <= Logical_Operator_out99_out1 XOR Logical_Operator_out103_out1;

  Logical_Operator_out230_out1 <= Logical_Operator_out100_out1 XOR Logical_Operator_out104_out1;

  Logical_Operator_out231_out1 <= Logical_Operator_out36_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out232_out1 <= in72 XOR in80;

  Logical_Operator_out233_out1 <= Logical_Operator_out169_out1 XOR Logical_Operator_out173_out1;

  Logical_Operator_out234_out1 <= Logical_Operator_out170_out1 XOR Logical_Operator_out174_out1;

  Logical_Operator_out235_out1 <= Logical_Operator_out171_out1 XOR Logical_Operator_out175_out1;

  Logical_Operator_out236_out1 <= Logical_Operator_out172_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out237_out1 <= Logical_Operator_out107_out1 XOR Logical_Operator_out111_out1;

  Logical_Operator_out238_out1 <= Logical_Operator_out108_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out239_out1 <= Logical_Operator_out44_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out240_out1 <= in88 XOR in96;

  Logical_Operator_out241_out1 <= Logical_Operator_out177_out1 XOR Logical_Operator_out181_out1;

  Logical_Operator_out242_out1 <= Logical_Operator_out178_out1 XOR Logical_Operator_out182_out1;

  Logical_Operator_out243_out1 <= Logical_Operator_out179_out1 XOR Logical_Operator_out183_out1;

  Logical_Operator_out244_out1 <= Logical_Operator_out180_out1 XOR Logical_Operator_out184_out1;

  Logical_Operator_out245_out1 <= Logical_Operator_out115_out1 XOR Logical_Operator_out119_out1;

  Logical_Operator_out246_out1 <= Logical_Operator_out116_out1 XOR Logical_Operator_out120_out1;

  Logical_Operator_out247_out1 <= Logical_Operator_out52_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out248_out1 <= in104 XOR in112;

  Logical_Operator_out249_out1 <= Logical_Operator_out185_out1 XOR Logical_Operator_out189_out1;

  Logical_Operator_out250_out1 <= Logical_Operator_out186_out1 XOR Logical_Operator_out190_out1;

  Logical_Operator_out251_out1 <= Logical_Operator_out187_out1 XOR Logical_Operator_out191_out1;

  Logical_Operator_out252_out1 <= Logical_Operator_out188_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out253_out1 <= Logical_Operator_out123_out1 XOR Logical_Operator_out127_out1;

  Logical_Operator_out254_out1 <= Logical_Operator_out124_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out255_out1 <= Logical_Operator_out60_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out256_out1 <= in120 XOR in128;

  Logical_Operator_out257_out1 <= Logical_Operator_out193_out1 XOR Logical_Operator_out201_out1;

  Logical_Operator_out258_out1 <= Logical_Operator_out194_out1 XOR Logical_Operator_out202_out1;

  Logical_Operator_out259_out1 <= Logical_Operator_out195_out1 XOR Logical_Operator_out203_out1;

  Logical_Operator_out260_out1 <= Logical_Operator_out196_out1 XOR Logical_Operator_out204_out1;

  Logical_Operator_out261_out1 <= Logical_Operator_out197_out1 XOR Logical_Operator_out205_out1;

  Logical_Operator_out262_out1 <= Logical_Operator_out198_out1 XOR Logical_Operator_out206_out1;

  Logical_Operator_out263_out1 <= Logical_Operator_out199_out1 XOR Logical_Operator_out207_out1;

  Logical_Operator_out264_out1 <= Logical_Operator_out200_out1 XOR Logical_Operator_out208_out1;

  Logical_Operator_out265_out1 <= Logical_Operator_out133_out1 XOR Logical_Operator_out141_out1;

  Logical_Operator_out266_out1 <= Logical_Operator_out134_out1 XOR Logical_Operator_out142_out1;

  Logical_Operator_out267_out1 <= Logical_Operator_out135_out1 XOR Logical_Operator_out143_out1;

  Logical_Operator_out268_out1 <= Logical_Operator_out136_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out269_out1 <= Logical_Operator_out71_out1 XOR Logical_Operator_out79_out1;

  Logical_Operator_out270_out1 <= Logical_Operator_out72_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out271_out1 <= Logical_Operator_out8_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out272_out1 <= in16 XOR in32;

  Logical_Operator_out273_out1 <= Logical_Operator_out209_out1 XOR Logical_Operator_out217_out1;

  Logical_Operator_out274_out1 <= Logical_Operator_out210_out1 XOR Logical_Operator_out218_out1;

  Logical_Operator_out275_out1 <= Logical_Operator_out211_out1 XOR Logical_Operator_out219_out1;

  Logical_Operator_out276_out1 <= Logical_Operator_out212_out1 XOR Logical_Operator_out220_out1;

  Logical_Operator_out277_out1 <= Logical_Operator_out213_out1 XOR Logical_Operator_out221_out1;

  Logical_Operator_out278_out1 <= Logical_Operator_out214_out1 XOR Logical_Operator_out222_out1;

  Logical_Operator_out279_out1 <= Logical_Operator_out215_out1 XOR Logical_Operator_out223_out1;

  Logical_Operator_out280_out1 <= Logical_Operator_out216_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out281_out1 <= Logical_Operator_out149_out1 XOR Logical_Operator_out157_out1;

  Logical_Operator_out282_out1 <= Logical_Operator_out150_out1 XOR Logical_Operator_out158_out1;

  Logical_Operator_out283_out1 <= Logical_Operator_out151_out1 XOR Logical_Operator_out159_out1;

  Logical_Operator_out284_out1 <= Logical_Operator_out152_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out285_out1 <= Logical_Operator_out87_out1 XOR Logical_Operator_out95_out1;

  Logical_Operator_out286_out1 <= Logical_Operator_out88_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out287_out1 <= Logical_Operator_out24_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out288_out1 <= in48 XOR in64;

  Logical_Operator_out289_out1 <= Logical_Operator_out225_out1 XOR Logical_Operator_out233_out1;

  Logical_Operator_out290_out1 <= Logical_Operator_out226_out1 XOR Logical_Operator_out234_out1;

  Logical_Operator_out291_out1 <= Logical_Operator_out227_out1 XOR Logical_Operator_out235_out1;

  Logical_Operator_out292_out1 <= Logical_Operator_out228_out1 XOR Logical_Operator_out236_out1;

  Logical_Operator_out293_out1 <= Logical_Operator_out229_out1 XOR Logical_Operator_out237_out1;

  Logical_Operator_out294_out1 <= Logical_Operator_out230_out1 XOR Logical_Operator_out238_out1;

  Logical_Operator_out295_out1 <= Logical_Operator_out231_out1 XOR Logical_Operator_out239_out1;

  Logical_Operator_out296_out1 <= Logical_Operator_out232_out1 XOR Logical_Operator_out240_out1;

  Logical_Operator_out297_out1 <= Logical_Operator_out165_out1 XOR Logical_Operator_out173_out1;

  Logical_Operator_out298_out1 <= Logical_Operator_out166_out1 XOR Logical_Operator_out174_out1;

  Logical_Operator_out299_out1 <= Logical_Operator_out167_out1 XOR Logical_Operator_out175_out1;

  Logical_Operator_out300_out1 <= Logical_Operator_out168_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out301_out1 <= Logical_Operator_out103_out1 XOR Logical_Operator_out111_out1;

  Logical_Operator_out302_out1 <= Logical_Operator_out104_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out303_out1 <= Logical_Operator_out40_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out304_out1 <= in80 XOR in96;

  Logical_Operator_out305_out1 <= Logical_Operator_out241_out1 XOR Logical_Operator_out249_out1;

  Logical_Operator_out306_out1 <= Logical_Operator_out242_out1 XOR Logical_Operator_out250_out1;

  Logical_Operator_out307_out1 <= Logical_Operator_out243_out1 XOR Logical_Operator_out251_out1;

  Logical_Operator_out308_out1 <= Logical_Operator_out244_out1 XOR Logical_Operator_out252_out1;

  Logical_Operator_out309_out1 <= Logical_Operator_out245_out1 XOR Logical_Operator_out253_out1;

  Logical_Operator_out310_out1 <= Logical_Operator_out246_out1 XOR Logical_Operator_out254_out1;

  Logical_Operator_out311_out1 <= Logical_Operator_out247_out1 XOR Logical_Operator_out255_out1;

  Logical_Operator_out312_out1 <= Logical_Operator_out248_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out313_out1 <= Logical_Operator_out181_out1 XOR Logical_Operator_out189_out1;

  Logical_Operator_out314_out1 <= Logical_Operator_out182_out1 XOR Logical_Operator_out190_out1;

  Logical_Operator_out315_out1 <= Logical_Operator_out183_out1 XOR Logical_Operator_out191_out1;

  Logical_Operator_out316_out1 <= Logical_Operator_out184_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out317_out1 <= Logical_Operator_out119_out1 XOR Logical_Operator_out127_out1;

  Logical_Operator_out318_out1 <= Logical_Operator_out120_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out319_out1 <= Logical_Operator_out56_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out320_out1 <= in112 XOR in128;

  Logical_Operator_out321_out1 <= Logical_Operator_out257_out1 XOR Logical_Operator_out273_out1;

  Logical_Operator_out322_out1 <= Logical_Operator_out258_out1 XOR Logical_Operator_out274_out1;

  Logical_Operator_out323_out1 <= Logical_Operator_out259_out1 XOR Logical_Operator_out275_out1;

  Logical_Operator_out324_out1 <= Logical_Operator_out260_out1 XOR Logical_Operator_out276_out1;

  Logical_Operator_out325_out1 <= Logical_Operator_out261_out1 XOR Logical_Operator_out277_out1;

  Logical_Operator_out326_out1 <= Logical_Operator_out262_out1 XOR Logical_Operator_out278_out1;

  Logical_Operator_out327_out1 <= Logical_Operator_out263_out1 XOR Logical_Operator_out279_out1;

  Logical_Operator_out328_out1 <= Logical_Operator_out264_out1 XOR Logical_Operator_out280_out1;

  Logical_Operator_out329_out1 <= Logical_Operator_out265_out1 XOR Logical_Operator_out281_out1;

  Logical_Operator_out330_out1 <= Logical_Operator_out266_out1 XOR Logical_Operator_out282_out1;

  Logical_Operator_out331_out1 <= Logical_Operator_out267_out1 XOR Logical_Operator_out283_out1;

  Logical_Operator_out332_out1 <= Logical_Operator_out268_out1 XOR Logical_Operator_out284_out1;

  Logical_Operator_out333_out1 <= Logical_Operator_out269_out1 XOR Logical_Operator_out285_out1;

  Logical_Operator_out334_out1 <= Logical_Operator_out270_out1 XOR Logical_Operator_out286_out1;

  Logical_Operator_out335_out1 <= Logical_Operator_out271_out1 XOR Logical_Operator_out287_out1;

  Logical_Operator_out336_out1 <= Logical_Operator_out272_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out337_out1 <= Logical_Operator_out201_out1 XOR Logical_Operator_out217_out1;

  Logical_Operator_out338_out1 <= Logical_Operator_out202_out1 XOR Logical_Operator_out218_out1;

  Logical_Operator_out339_out1 <= Logical_Operator_out203_out1 XOR Logical_Operator_out219_out1;

  Logical_Operator_out340_out1 <= Logical_Operator_out204_out1 XOR Logical_Operator_out220_out1;

  Logical_Operator_out341_out1 <= Logical_Operator_out205_out1 XOR Logical_Operator_out221_out1;

  Logical_Operator_out342_out1 <= Logical_Operator_out206_out1 XOR Logical_Operator_out222_out1;

  Logical_Operator_out343_out1 <= Logical_Operator_out207_out1 XOR Logical_Operator_out223_out1;

  Logical_Operator_out344_out1 <= Logical_Operator_out208_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out345_out1 <= Logical_Operator_out141_out1 XOR Logical_Operator_out157_out1;

  Logical_Operator_out346_out1 <= Logical_Operator_out142_out1 XOR Logical_Operator_out158_out1;

  Logical_Operator_out347_out1 <= Logical_Operator_out143_out1 XOR Logical_Operator_out159_out1;

  Logical_Operator_out348_out1 <= Logical_Operator_out144_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out349_out1 <= Logical_Operator_out79_out1 XOR Logical_Operator_out95_out1;

  Logical_Operator_out350_out1 <= Logical_Operator_out80_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out351_out1 <= Logical_Operator_out16_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out352_out1 <= in32 XOR in64;

  Logical_Operator_out353_out1 <= Logical_Operator_out289_out1 XOR Logical_Operator_out305_out1;

  Logical_Operator_out354_out1 <= Logical_Operator_out290_out1 XOR Logical_Operator_out306_out1;

  Logical_Operator_out355_out1 <= Logical_Operator_out291_out1 XOR Logical_Operator_out307_out1;

  Logical_Operator_out356_out1 <= Logical_Operator_out292_out1 XOR Logical_Operator_out308_out1;

  Logical_Operator_out357_out1 <= Logical_Operator_out293_out1 XOR Logical_Operator_out309_out1;

  Logical_Operator_out358_out1 <= Logical_Operator_out294_out1 XOR Logical_Operator_out310_out1;

  Logical_Operator_out359_out1 <= Logical_Operator_out295_out1 XOR Logical_Operator_out311_out1;

  Logical_Operator_out360_out1 <= Logical_Operator_out296_out1 XOR Logical_Operator_out312_out1;

  Logical_Operator_out361_out1 <= Logical_Operator_out297_out1 XOR Logical_Operator_out313_out1;

  Logical_Operator_out362_out1 <= Logical_Operator_out298_out1 XOR Logical_Operator_out314_out1;

  Logical_Operator_out363_out1 <= Logical_Operator_out299_out1 XOR Logical_Operator_out315_out1;

  Logical_Operator_out364_out1 <= Logical_Operator_out300_out1 XOR Logical_Operator_out316_out1;

  Logical_Operator_out365_out1 <= Logical_Operator_out301_out1 XOR Logical_Operator_out317_out1;

  Logical_Operator_out366_out1 <= Logical_Operator_out302_out1 XOR Logical_Operator_out318_out1;

  Logical_Operator_out367_out1 <= Logical_Operator_out303_out1 XOR Logical_Operator_out319_out1;

  Logical_Operator_out368_out1 <= Logical_Operator_out304_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out369_out1 <= Logical_Operator_out233_out1 XOR Logical_Operator_out249_out1;

  Logical_Operator_out370_out1 <= Logical_Operator_out234_out1 XOR Logical_Operator_out250_out1;

  Logical_Operator_out371_out1 <= Logical_Operator_out235_out1 XOR Logical_Operator_out251_out1;

  Logical_Operator_out372_out1 <= Logical_Operator_out236_out1 XOR Logical_Operator_out252_out1;

  Logical_Operator_out373_out1 <= Logical_Operator_out237_out1 XOR Logical_Operator_out253_out1;

  Logical_Operator_out374_out1 <= Logical_Operator_out238_out1 XOR Logical_Operator_out254_out1;

  Logical_Operator_out375_out1 <= Logical_Operator_out239_out1 XOR Logical_Operator_out255_out1;

  Logical_Operator_out376_out1 <= Logical_Operator_out240_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out377_out1 <= Logical_Operator_out173_out1 XOR Logical_Operator_out189_out1;

  Logical_Operator_out378_out1 <= Logical_Operator_out174_out1 XOR Logical_Operator_out190_out1;

  Logical_Operator_out379_out1 <= Logical_Operator_out175_out1 XOR Logical_Operator_out191_out1;

  Logical_Operator_out380_out1 <= Logical_Operator_out176_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out381_out1 <= Logical_Operator_out111_out1 XOR Logical_Operator_out127_out1;

  Logical_Operator_out382_out1 <= Logical_Operator_out112_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out383_out1 <= Logical_Operator_out48_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out384_out1 <= in96 XOR in128;

  Logical_Operator_out385_out1 <= Logical_Operator_out321_out1 XOR Logical_Operator_out353_out1;

  Logical_Operator_out386_out1 <= Logical_Operator_out322_out1 XOR Logical_Operator_out354_out1;

  Logical_Operator_out387_out1 <= Logical_Operator_out323_out1 XOR Logical_Operator_out355_out1;

  Logical_Operator_out388_out1 <= Logical_Operator_out324_out1 XOR Logical_Operator_out356_out1;

  Logical_Operator_out389_out1 <= Logical_Operator_out325_out1 XOR Logical_Operator_out357_out1;

  Logical_Operator_out390_out1 <= Logical_Operator_out326_out1 XOR Logical_Operator_out358_out1;

  Logical_Operator_out391_out1 <= Logical_Operator_out327_out1 XOR Logical_Operator_out359_out1;

  Logical_Operator_out392_out1 <= Logical_Operator_out328_out1 XOR Logical_Operator_out360_out1;

  Logical_Operator_out393_out1 <= Logical_Operator_out329_out1 XOR Logical_Operator_out361_out1;

  Logical_Operator_out394_out1 <= Logical_Operator_out330_out1 XOR Logical_Operator_out362_out1;

  Logical_Operator_out395_out1 <= Logical_Operator_out331_out1 XOR Logical_Operator_out363_out1;

  Logical_Operator_out396_out1 <= Logical_Operator_out332_out1 XOR Logical_Operator_out364_out1;

  Logical_Operator_out397_out1 <= Logical_Operator_out333_out1 XOR Logical_Operator_out365_out1;

  Logical_Operator_out398_out1 <= Logical_Operator_out334_out1 XOR Logical_Operator_out366_out1;

  Logical_Operator_out399_out1 <= Logical_Operator_out335_out1 XOR Logical_Operator_out367_out1;

  Logical_Operator_out400_out1 <= Logical_Operator_out336_out1 XOR Logical_Operator_out368_out1;

  Logical_Operator_out401_out1 <= Logical_Operator_out337_out1 XOR Logical_Operator_out369_out1;

  Logical_Operator_out402_out1 <= Logical_Operator_out338_out1 XOR Logical_Operator_out370_out1;

  Logical_Operator_out403_out1 <= Logical_Operator_out339_out1 XOR Logical_Operator_out371_out1;

  Logical_Operator_out404_out1 <= Logical_Operator_out340_out1 XOR Logical_Operator_out372_out1;

  Logical_Operator_out405_out1 <= Logical_Operator_out341_out1 XOR Logical_Operator_out373_out1;

  Logical_Operator_out406_out1 <= Logical_Operator_out342_out1 XOR Logical_Operator_out374_out1;

  Logical_Operator_out407_out1 <= Logical_Operator_out343_out1 XOR Logical_Operator_out375_out1;

  Logical_Operator_out408_out1 <= Logical_Operator_out344_out1 XOR Logical_Operator_out376_out1;

  Logical_Operator_out409_out1 <= Logical_Operator_out345_out1 XOR Logical_Operator_out377_out1;

  Logical_Operator_out410_out1 <= Logical_Operator_out346_out1 XOR Logical_Operator_out378_out1;

  Logical_Operator_out411_out1 <= Logical_Operator_out347_out1 XOR Logical_Operator_out379_out1;

  Logical_Operator_out412_out1 <= Logical_Operator_out348_out1 XOR Logical_Operator_out380_out1;

  Logical_Operator_out413_out1 <= Logical_Operator_out349_out1 XOR Logical_Operator_out381_out1;

  Logical_Operator_out414_out1 <= Logical_Operator_out350_out1 XOR Logical_Operator_out382_out1;

  Logical_Operator_out415_out1 <= Logical_Operator_out351_out1 XOR Logical_Operator_out383_out1;

  Logical_Operator_out416_out1 <= Logical_Operator_out352_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out417_out1 <= Logical_Operator_out273_out1 XOR Logical_Operator_out305_out1;

  Logical_Operator_out418_out1 <= Logical_Operator_out274_out1 XOR Logical_Operator_out306_out1;

  Logical_Operator_out419_out1 <= Logical_Operator_out275_out1 XOR Logical_Operator_out307_out1;

  Logical_Operator_out420_out1 <= Logical_Operator_out276_out1 XOR Logical_Operator_out308_out1;

  Logical_Operator_out421_out1 <= Logical_Operator_out277_out1 XOR Logical_Operator_out309_out1;

  Logical_Operator_out422_out1 <= Logical_Operator_out278_out1 XOR Logical_Operator_out310_out1;

  Logical_Operator_out423_out1 <= Logical_Operator_out279_out1 XOR Logical_Operator_out311_out1;

  Logical_Operator_out424_out1 <= Logical_Operator_out280_out1 XOR Logical_Operator_out312_out1;

  Logical_Operator_out425_out1 <= Logical_Operator_out281_out1 XOR Logical_Operator_out313_out1;

  Logical_Operator_out426_out1 <= Logical_Operator_out282_out1 XOR Logical_Operator_out314_out1;

  Logical_Operator_out427_out1 <= Logical_Operator_out283_out1 XOR Logical_Operator_out315_out1;

  Logical_Operator_out428_out1 <= Logical_Operator_out284_out1 XOR Logical_Operator_out316_out1;

  Logical_Operator_out429_out1 <= Logical_Operator_out285_out1 XOR Logical_Operator_out317_out1;

  Logical_Operator_out430_out1 <= Logical_Operator_out286_out1 XOR Logical_Operator_out318_out1;

  Logical_Operator_out431_out1 <= Logical_Operator_out287_out1 XOR Logical_Operator_out319_out1;

  Logical_Operator_out432_out1 <= Logical_Operator_out288_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out433_out1 <= Logical_Operator_out217_out1 XOR Logical_Operator_out249_out1;

  Logical_Operator_out434_out1 <= Logical_Operator_out218_out1 XOR Logical_Operator_out250_out1;

  Logical_Operator_out435_out1 <= Logical_Operator_out219_out1 XOR Logical_Operator_out251_out1;

  Logical_Operator_out436_out1 <= Logical_Operator_out220_out1 XOR Logical_Operator_out252_out1;

  Logical_Operator_out437_out1 <= Logical_Operator_out221_out1 XOR Logical_Operator_out253_out1;

  Logical_Operator_out438_out1 <= Logical_Operator_out222_out1 XOR Logical_Operator_out254_out1;

  Logical_Operator_out439_out1 <= Logical_Operator_out223_out1 XOR Logical_Operator_out255_out1;

  Logical_Operator_out440_out1 <= Logical_Operator_out224_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out441_out1 <= Logical_Operator_out157_out1 XOR Logical_Operator_out189_out1;

  Logical_Operator_out442_out1 <= Logical_Operator_out158_out1 XOR Logical_Operator_out190_out1;

  Logical_Operator_out443_out1 <= Logical_Operator_out159_out1 XOR Logical_Operator_out191_out1;

  Logical_Operator_out444_out1 <= Logical_Operator_out160_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out445_out1 <= Logical_Operator_out95_out1 XOR Logical_Operator_out127_out1;

  Logical_Operator_out446_out1 <= Logical_Operator_out96_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out447_out1 <= Logical_Operator_out32_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out448_out1 <= in64 XOR in128;

  out1 <= Logical_Operator_out385_out1;

  out2 <= Logical_Operator_out386_out1;

  out3 <= Logical_Operator_out387_out1;

  out4 <= Logical_Operator_out388_out1;

  out5 <= Logical_Operator_out389_out1;

  out6 <= Logical_Operator_out390_out1;

  out7 <= Logical_Operator_out391_out1;

  out8 <= Logical_Operator_out392_out1;

  out9 <= Logical_Operator_out393_out1;

  out10 <= Logical_Operator_out394_out1;

  out11 <= Logical_Operator_out395_out1;

  out12 <= Logical_Operator_out396_out1;

  out13 <= Logical_Operator_out397_out1;

  out14 <= Logical_Operator_out398_out1;

  out15 <= Logical_Operator_out399_out1;

  out16 <= Logical_Operator_out400_out1;

  out17 <= Logical_Operator_out401_out1;

  out18 <= Logical_Operator_out402_out1;

  out19 <= Logical_Operator_out403_out1;

  out20 <= Logical_Operator_out404_out1;

  out21 <= Logical_Operator_out405_out1;

  out22 <= Logical_Operator_out406_out1;

  out23 <= Logical_Operator_out407_out1;

  out24 <= Logical_Operator_out408_out1;

  out25 <= Logical_Operator_out409_out1;

  out26 <= Logical_Operator_out410_out1;

  out27 <= Logical_Operator_out411_out1;

  out28 <= Logical_Operator_out412_out1;

  out29 <= Logical_Operator_out413_out1;

  out30 <= Logical_Operator_out414_out1;

  out31 <= Logical_Operator_out415_out1;

  out32 <= Logical_Operator_out416_out1;

  out33 <= Logical_Operator_out417_out1;

  out34 <= Logical_Operator_out418_out1;

  out35 <= Logical_Operator_out419_out1;

  out36 <= Logical_Operator_out420_out1;

  out37 <= Logical_Operator_out421_out1;

  out38 <= Logical_Operator_out422_out1;

  out39 <= Logical_Operator_out423_out1;

  out40 <= Logical_Operator_out424_out1;

  out41 <= Logical_Operator_out425_out1;

  out42 <= Logical_Operator_out426_out1;

  out43 <= Logical_Operator_out427_out1;

  out44 <= Logical_Operator_out428_out1;

  out45 <= Logical_Operator_out429_out1;

  out46 <= Logical_Operator_out430_out1;

  out47 <= Logical_Operator_out431_out1;

  out48 <= Logical_Operator_out432_out1;

  out49 <= Logical_Operator_out433_out1;

  out50 <= Logical_Operator_out434_out1;

  out51 <= Logical_Operator_out435_out1;

  out52 <= Logical_Operator_out436_out1;

  out53 <= Logical_Operator_out437_out1;

  out54 <= Logical_Operator_out438_out1;

  out55 <= Logical_Operator_out439_out1;

  out56 <= Logical_Operator_out440_out1;

  out57 <= Logical_Operator_out441_out1;

  out58 <= Logical_Operator_out442_out1;

  out59 <= Logical_Operator_out443_out1;

  out60 <= Logical_Operator_out444_out1;

  out61 <= Logical_Operator_out445_out1;

  out62 <= Logical_Operator_out446_out1;

  out63 <= Logical_Operator_out447_out1;

  out64 <= Logical_Operator_out448_out1;

  out65 <= Logical_Operator_out353_out1;

  out66 <= Logical_Operator_out354_out1;

  out67 <= Logical_Operator_out355_out1;

  out68 <= Logical_Operator_out356_out1;

  out69 <= Logical_Operator_out357_out1;

  out70 <= Logical_Operator_out358_out1;

  out71 <= Logical_Operator_out359_out1;

  out72 <= Logical_Operator_out360_out1;

  out73 <= Logical_Operator_out361_out1;

  out74 <= Logical_Operator_out362_out1;

  out75 <= Logical_Operator_out363_out1;

  out76 <= Logical_Operator_out364_out1;

  out77 <= Logical_Operator_out365_out1;

  out78 <= Logical_Operator_out366_out1;

  out79 <= Logical_Operator_out367_out1;

  out80 <= Logical_Operator_out368_out1;

  out81 <= Logical_Operator_out369_out1;

  out82 <= Logical_Operator_out370_out1;

  out83 <= Logical_Operator_out371_out1;

  out84 <= Logical_Operator_out372_out1;

  out85 <= Logical_Operator_out373_out1;

  out86 <= Logical_Operator_out374_out1;

  out87 <= Logical_Operator_out375_out1;

  out88 <= Logical_Operator_out376_out1;

  out89 <= Logical_Operator_out377_out1;

  out90 <= Logical_Operator_out378_out1;

  out91 <= Logical_Operator_out379_out1;

  out92 <= Logical_Operator_out380_out1;

  out93 <= Logical_Operator_out381_out1;

  out94 <= Logical_Operator_out382_out1;

  out95 <= Logical_Operator_out383_out1;

  out96 <= Logical_Operator_out384_out1;

  out97 <= Logical_Operator_out305_out1;

  out98 <= Logical_Operator_out306_out1;

  out99 <= Logical_Operator_out307_out1;

  out100 <= Logical_Operator_out308_out1;

  out101 <= Logical_Operator_out309_out1;

  out102 <= Logical_Operator_out310_out1;

  out103 <= Logical_Operator_out311_out1;

  out104 <= Logical_Operator_out312_out1;

  out105 <= Logical_Operator_out313_out1;

  out106 <= Logical_Operator_out314_out1;

  out107 <= Logical_Operator_out315_out1;

  out108 <= Logical_Operator_out316_out1;

  out109 <= Logical_Operator_out317_out1;

  out110 <= Logical_Operator_out318_out1;

  out111 <= Logical_Operator_out319_out1;

  out112 <= Logical_Operator_out320_out1;

  out113 <= Logical_Operator_out249_out1;

  out114 <= Logical_Operator_out250_out1;

  out115 <= Logical_Operator_out251_out1;

  out116 <= Logical_Operator_out252_out1;

  out117 <= Logical_Operator_out253_out1;

  out118 <= Logical_Operator_out254_out1;

  out119 <= Logical_Operator_out255_out1;

  out120 <= Logical_Operator_out256_out1;

  out121 <= Logical_Operator_out189_out1;

  out122 <= Logical_Operator_out190_out1;

  out123 <= Logical_Operator_out191_out1;

  out124 <= Logical_Operator_out192_out1;

  out125 <= Logical_Operator_out127_out1;

  out126 <= Logical_Operator_out128_out1;

  out127 <= Logical_Operator_out64_out1;

  out128 <= in128;

END rtl;
