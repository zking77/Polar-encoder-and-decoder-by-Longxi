LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY encoderN256 IS
PORT( 
	in1                               :   IN    std_logic;
	in2                               :   IN    std_logic;
	in3                               :   IN    std_logic;
	in4                               :   IN    std_logic;
	in5                               :   IN    std_logic;
	in6                               :   IN    std_logic;
	in7                               :   IN    std_logic;
	in8                               :   IN    std_logic;
	in9                               :   IN    std_logic;
	in10                               :   IN    std_logic;
	in11                               :   IN    std_logic;
	in12                               :   IN    std_logic;
	in13                               :   IN    std_logic;
	in14                               :   IN    std_logic;
	in15                               :   IN    std_logic;
	in16                               :   IN    std_logic;
	in17                               :   IN    std_logic;
	in18                               :   IN    std_logic;
	in19                               :   IN    std_logic;
	in20                               :   IN    std_logic;
	in21                               :   IN    std_logic;
	in22                               :   IN    std_logic;
	in23                               :   IN    std_logic;
	in24                               :   IN    std_logic;
	in25                               :   IN    std_logic;
	in26                               :   IN    std_logic;
	in27                               :   IN    std_logic;
	in28                               :   IN    std_logic;
	in29                               :   IN    std_logic;
	in30                               :   IN    std_logic;
	in31                               :   IN    std_logic;
	in32                               :   IN    std_logic;
	in33                               :   IN    std_logic;
	in34                               :   IN    std_logic;
	in35                               :   IN    std_logic;
	in36                               :   IN    std_logic;
	in37                               :   IN    std_logic;
	in38                               :   IN    std_logic;
	in39                               :   IN    std_logic;
	in40                               :   IN    std_logic;
	in41                               :   IN    std_logic;
	in42                               :   IN    std_logic;
	in43                               :   IN    std_logic;
	in44                               :   IN    std_logic;
	in45                               :   IN    std_logic;
	in46                               :   IN    std_logic;
	in47                               :   IN    std_logic;
	in48                               :   IN    std_logic;
	in49                               :   IN    std_logic;
	in50                               :   IN    std_logic;
	in51                               :   IN    std_logic;
	in52                               :   IN    std_logic;
	in53                               :   IN    std_logic;
	in54                               :   IN    std_logic;
	in55                               :   IN    std_logic;
	in56                               :   IN    std_logic;
	in57                               :   IN    std_logic;
	in58                               :   IN    std_logic;
	in59                               :   IN    std_logic;
	in60                               :   IN    std_logic;
	in61                               :   IN    std_logic;
	in62                               :   IN    std_logic;
	in63                               :   IN    std_logic;
	in64                               :   IN    std_logic;
	in65                               :   IN    std_logic;
	in66                               :   IN    std_logic;
	in67                               :   IN    std_logic;
	in68                               :   IN    std_logic;
	in69                               :   IN    std_logic;
	in70                               :   IN    std_logic;
	in71                               :   IN    std_logic;
	in72                               :   IN    std_logic;
	in73                               :   IN    std_logic;
	in74                               :   IN    std_logic;
	in75                               :   IN    std_logic;
	in76                               :   IN    std_logic;
	in77                               :   IN    std_logic;
	in78                               :   IN    std_logic;
	in79                               :   IN    std_logic;
	in80                               :   IN    std_logic;
	in81                               :   IN    std_logic;
	in82                               :   IN    std_logic;
	in83                               :   IN    std_logic;
	in84                               :   IN    std_logic;
	in85                               :   IN    std_logic;
	in86                               :   IN    std_logic;
	in87                               :   IN    std_logic;
	in88                               :   IN    std_logic;
	in89                               :   IN    std_logic;
	in90                               :   IN    std_logic;
	in91                               :   IN    std_logic;
	in92                               :   IN    std_logic;
	in93                               :   IN    std_logic;
	in94                               :   IN    std_logic;
	in95                               :   IN    std_logic;
	in96                               :   IN    std_logic;
	in97                               :   IN    std_logic;
	in98                               :   IN    std_logic;
	in99                               :   IN    std_logic;
	in100                               :   IN    std_logic;
	in101                               :   IN    std_logic;
	in102                               :   IN    std_logic;
	in103                               :   IN    std_logic;
	in104                               :   IN    std_logic;
	in105                               :   IN    std_logic;
	in106                               :   IN    std_logic;
	in107                               :   IN    std_logic;
	in108                               :   IN    std_logic;
	in109                               :   IN    std_logic;
	in110                               :   IN    std_logic;
	in111                               :   IN    std_logic;
	in112                               :   IN    std_logic;
	in113                               :   IN    std_logic;
	in114                               :   IN    std_logic;
	in115                               :   IN    std_logic;
	in116                               :   IN    std_logic;
	in117                               :   IN    std_logic;
	in118                               :   IN    std_logic;
	in119                               :   IN    std_logic;
	in120                               :   IN    std_logic;
	in121                               :   IN    std_logic;
	in122                               :   IN    std_logic;
	in123                               :   IN    std_logic;
	in124                               :   IN    std_logic;
	in125                               :   IN    std_logic;
	in126                               :   IN    std_logic;
	in127                               :   IN    std_logic;
	in128                               :   IN    std_logic;
	in129                               :   IN    std_logic;
	in130                               :   IN    std_logic;
	in131                               :   IN    std_logic;
	in132                               :   IN    std_logic;
	in133                               :   IN    std_logic;
	in134                               :   IN    std_logic;
	in135                               :   IN    std_logic;
	in136                               :   IN    std_logic;
	in137                               :   IN    std_logic;
	in138                               :   IN    std_logic;
	in139                               :   IN    std_logic;
	in140                               :   IN    std_logic;
	in141                               :   IN    std_logic;
	in142                               :   IN    std_logic;
	in143                               :   IN    std_logic;
	in144                               :   IN    std_logic;
	in145                               :   IN    std_logic;
	in146                               :   IN    std_logic;
	in147                               :   IN    std_logic;
	in148                               :   IN    std_logic;
	in149                               :   IN    std_logic;
	in150                               :   IN    std_logic;
	in151                               :   IN    std_logic;
	in152                               :   IN    std_logic;
	in153                               :   IN    std_logic;
	in154                               :   IN    std_logic;
	in155                               :   IN    std_logic;
	in156                               :   IN    std_logic;
	in157                               :   IN    std_logic;
	in158                               :   IN    std_logic;
	in159                               :   IN    std_logic;
	in160                               :   IN    std_logic;
	in161                               :   IN    std_logic;
	in162                               :   IN    std_logic;
	in163                               :   IN    std_logic;
	in164                               :   IN    std_logic;
	in165                               :   IN    std_logic;
	in166                               :   IN    std_logic;
	in167                               :   IN    std_logic;
	in168                               :   IN    std_logic;
	in169                               :   IN    std_logic;
	in170                               :   IN    std_logic;
	in171                               :   IN    std_logic;
	in172                               :   IN    std_logic;
	in173                               :   IN    std_logic;
	in174                               :   IN    std_logic;
	in175                               :   IN    std_logic;
	in176                               :   IN    std_logic;
	in177                               :   IN    std_logic;
	in178                               :   IN    std_logic;
	in179                               :   IN    std_logic;
	in180                               :   IN    std_logic;
	in181                               :   IN    std_logic;
	in182                               :   IN    std_logic;
	in183                               :   IN    std_logic;
	in184                               :   IN    std_logic;
	in185                               :   IN    std_logic;
	in186                               :   IN    std_logic;
	in187                               :   IN    std_logic;
	in188                               :   IN    std_logic;
	in189                               :   IN    std_logic;
	in190                               :   IN    std_logic;
	in191                               :   IN    std_logic;
	in192                               :   IN    std_logic;
	in193                               :   IN    std_logic;
	in194                               :   IN    std_logic;
	in195                               :   IN    std_logic;
	in196                               :   IN    std_logic;
	in197                               :   IN    std_logic;
	in198                               :   IN    std_logic;
	in199                               :   IN    std_logic;
	in200                               :   IN    std_logic;
	in201                               :   IN    std_logic;
	in202                               :   IN    std_logic;
	in203                               :   IN    std_logic;
	in204                               :   IN    std_logic;
	in205                               :   IN    std_logic;
	in206                               :   IN    std_logic;
	in207                               :   IN    std_logic;
	in208                               :   IN    std_logic;
	in209                               :   IN    std_logic;
	in210                               :   IN    std_logic;
	in211                               :   IN    std_logic;
	in212                               :   IN    std_logic;
	in213                               :   IN    std_logic;
	in214                               :   IN    std_logic;
	in215                               :   IN    std_logic;
	in216                               :   IN    std_logic;
	in217                               :   IN    std_logic;
	in218                               :   IN    std_logic;
	in219                               :   IN    std_logic;
	in220                               :   IN    std_logic;
	in221                               :   IN    std_logic;
	in222                               :   IN    std_logic;
	in223                               :   IN    std_logic;
	in224                               :   IN    std_logic;
	in225                               :   IN    std_logic;
	in226                               :   IN    std_logic;
	in227                               :   IN    std_logic;
	in228                               :   IN    std_logic;
	in229                               :   IN    std_logic;
	in230                               :   IN    std_logic;
	in231                               :   IN    std_logic;
	in232                               :   IN    std_logic;
	in233                               :   IN    std_logic;
	in234                               :   IN    std_logic;
	in235                               :   IN    std_logic;
	in236                               :   IN    std_logic;
	in237                               :   IN    std_logic;
	in238                               :   IN    std_logic;
	in239                               :   IN    std_logic;
	in240                               :   IN    std_logic;
	in241                               :   IN    std_logic;
	in242                               :   IN    std_logic;
	in243                               :   IN    std_logic;
	in244                               :   IN    std_logic;
	in245                               :   IN    std_logic;
	in246                               :   IN    std_logic;
	in247                               :   IN    std_logic;
	in248                               :   IN    std_logic;
	in249                               :   IN    std_logic;
	in250                               :   IN    std_logic;
	in251                               :   IN    std_logic;
	in252                               :   IN    std_logic;
	in253                               :   IN    std_logic;
	in254                               :   IN    std_logic;
	in255                               :   IN    std_logic;
	in256                               :   IN    std_logic;
	out1                               :   OUT    std_logic;
	out2                               :   OUT    std_logic;
	out3                               :   OUT    std_logic;
	out4                               :   OUT    std_logic;
	out5                               :   OUT    std_logic;
	out6                               :   OUT    std_logic;
	out7                               :   OUT    std_logic;
	out8                               :   OUT    std_logic;
	out9                               :   OUT    std_logic;
	out10                               :   OUT    std_logic;
	out11                               :   OUT    std_logic;
	out12                               :   OUT    std_logic;
	out13                               :   OUT    std_logic;
	out14                               :   OUT    std_logic;
	out15                               :   OUT    std_logic;
	out16                               :   OUT    std_logic;
	out17                               :   OUT    std_logic;
	out18                               :   OUT    std_logic;
	out19                               :   OUT    std_logic;
	out20                               :   OUT    std_logic;
	out21                               :   OUT    std_logic;
	out22                               :   OUT    std_logic;
	out23                               :   OUT    std_logic;
	out24                               :   OUT    std_logic;
	out25                               :   OUT    std_logic;
	out26                               :   OUT    std_logic;
	out27                               :   OUT    std_logic;
	out28                               :   OUT    std_logic;
	out29                               :   OUT    std_logic;
	out30                               :   OUT    std_logic;
	out31                               :   OUT    std_logic;
	out32                               :   OUT    std_logic;
	out33                               :   OUT    std_logic;
	out34                               :   OUT    std_logic;
	out35                               :   OUT    std_logic;
	out36                               :   OUT    std_logic;
	out37                               :   OUT    std_logic;
	out38                               :   OUT    std_logic;
	out39                               :   OUT    std_logic;
	out40                               :   OUT    std_logic;
	out41                               :   OUT    std_logic;
	out42                               :   OUT    std_logic;
	out43                               :   OUT    std_logic;
	out44                               :   OUT    std_logic;
	out45                               :   OUT    std_logic;
	out46                               :   OUT    std_logic;
	out47                               :   OUT    std_logic;
	out48                               :   OUT    std_logic;
	out49                               :   OUT    std_logic;
	out50                               :   OUT    std_logic;
	out51                               :   OUT    std_logic;
	out52                               :   OUT    std_logic;
	out53                               :   OUT    std_logic;
	out54                               :   OUT    std_logic;
	out55                               :   OUT    std_logic;
	out56                               :   OUT    std_logic;
	out57                               :   OUT    std_logic;
	out58                               :   OUT    std_logic;
	out59                               :   OUT    std_logic;
	out60                               :   OUT    std_logic;
	out61                               :   OUT    std_logic;
	out62                               :   OUT    std_logic;
	out63                               :   OUT    std_logic;
	out64                               :   OUT    std_logic;
	out65                               :   OUT    std_logic;
	out66                               :   OUT    std_logic;
	out67                               :   OUT    std_logic;
	out68                               :   OUT    std_logic;
	out69                               :   OUT    std_logic;
	out70                               :   OUT    std_logic;
	out71                               :   OUT    std_logic;
	out72                               :   OUT    std_logic;
	out73                               :   OUT    std_logic;
	out74                               :   OUT    std_logic;
	out75                               :   OUT    std_logic;
	out76                               :   OUT    std_logic;
	out77                               :   OUT    std_logic;
	out78                               :   OUT    std_logic;
	out79                               :   OUT    std_logic;
	out80                               :   OUT    std_logic;
	out81                               :   OUT    std_logic;
	out82                               :   OUT    std_logic;
	out83                               :   OUT    std_logic;
	out84                               :   OUT    std_logic;
	out85                               :   OUT    std_logic;
	out86                               :   OUT    std_logic;
	out87                               :   OUT    std_logic;
	out88                               :   OUT    std_logic;
	out89                               :   OUT    std_logic;
	out90                               :   OUT    std_logic;
	out91                               :   OUT    std_logic;
	out92                               :   OUT    std_logic;
	out93                               :   OUT    std_logic;
	out94                               :   OUT    std_logic;
	out95                               :   OUT    std_logic;
	out96                               :   OUT    std_logic;
	out97                               :   OUT    std_logic;
	out98                               :   OUT    std_logic;
	out99                               :   OUT    std_logic;
	out100                               :   OUT    std_logic;
	out101                               :   OUT    std_logic;
	out102                               :   OUT    std_logic;
	out103                               :   OUT    std_logic;
	out104                               :   OUT    std_logic;
	out105                               :   OUT    std_logic;
	out106                               :   OUT    std_logic;
	out107                               :   OUT    std_logic;
	out108                               :   OUT    std_logic;
	out109                               :   OUT    std_logic;
	out110                               :   OUT    std_logic;
	out111                               :   OUT    std_logic;
	out112                               :   OUT    std_logic;
	out113                               :   OUT    std_logic;
	out114                               :   OUT    std_logic;
	out115                               :   OUT    std_logic;
	out116                               :   OUT    std_logic;
	out117                               :   OUT    std_logic;
	out118                               :   OUT    std_logic;
	out119                               :   OUT    std_logic;
	out120                               :   OUT    std_logic;
	out121                               :   OUT    std_logic;
	out122                               :   OUT    std_logic;
	out123                               :   OUT    std_logic;
	out124                               :   OUT    std_logic;
	out125                               :   OUT    std_logic;
	out126                               :   OUT    std_logic;
	out127                               :   OUT    std_logic;
	out128                               :   OUT    std_logic;
	out129                               :   OUT    std_logic;
	out130                               :   OUT    std_logic;
	out131                               :   OUT    std_logic;
	out132                               :   OUT    std_logic;
	out133                               :   OUT    std_logic;
	out134                               :   OUT    std_logic;
	out135                               :   OUT    std_logic;
	out136                               :   OUT    std_logic;
	out137                               :   OUT    std_logic;
	out138                               :   OUT    std_logic;
	out139                               :   OUT    std_logic;
	out140                               :   OUT    std_logic;
	out141                               :   OUT    std_logic;
	out142                               :   OUT    std_logic;
	out143                               :   OUT    std_logic;
	out144                               :   OUT    std_logic;
	out145                               :   OUT    std_logic;
	out146                               :   OUT    std_logic;
	out147                               :   OUT    std_logic;
	out148                               :   OUT    std_logic;
	out149                               :   OUT    std_logic;
	out150                               :   OUT    std_logic;
	out151                               :   OUT    std_logic;
	out152                               :   OUT    std_logic;
	out153                               :   OUT    std_logic;
	out154                               :   OUT    std_logic;
	out155                               :   OUT    std_logic;
	out156                               :   OUT    std_logic;
	out157                               :   OUT    std_logic;
	out158                               :   OUT    std_logic;
	out159                               :   OUT    std_logic;
	out160                               :   OUT    std_logic;
	out161                               :   OUT    std_logic;
	out162                               :   OUT    std_logic;
	out163                               :   OUT    std_logic;
	out164                               :   OUT    std_logic;
	out165                               :   OUT    std_logic;
	out166                               :   OUT    std_logic;
	out167                               :   OUT    std_logic;
	out168                               :   OUT    std_logic;
	out169                               :   OUT    std_logic;
	out170                               :   OUT    std_logic;
	out171                               :   OUT    std_logic;
	out172                               :   OUT    std_logic;
	out173                               :   OUT    std_logic;
	out174                               :   OUT    std_logic;
	out175                               :   OUT    std_logic;
	out176                               :   OUT    std_logic;
	out177                               :   OUT    std_logic;
	out178                               :   OUT    std_logic;
	out179                               :   OUT    std_logic;
	out180                               :   OUT    std_logic;
	out181                               :   OUT    std_logic;
	out182                               :   OUT    std_logic;
	out183                               :   OUT    std_logic;
	out184                               :   OUT    std_logic;
	out185                               :   OUT    std_logic;
	out186                               :   OUT    std_logic;
	out187                               :   OUT    std_logic;
	out188                               :   OUT    std_logic;
	out189                               :   OUT    std_logic;
	out190                               :   OUT    std_logic;
	out191                               :   OUT    std_logic;
	out192                               :   OUT    std_logic;
	out193                               :   OUT    std_logic;
	out194                               :   OUT    std_logic;
	out195                               :   OUT    std_logic;
	out196                               :   OUT    std_logic;
	out197                               :   OUT    std_logic;
	out198                               :   OUT    std_logic;
	out199                               :   OUT    std_logic;
	out200                               :   OUT    std_logic;
	out201                               :   OUT    std_logic;
	out202                               :   OUT    std_logic;
	out203                               :   OUT    std_logic;
	out204                               :   OUT    std_logic;
	out205                               :   OUT    std_logic;
	out206                               :   OUT    std_logic;
	out207                               :   OUT    std_logic;
	out208                               :   OUT    std_logic;
	out209                               :   OUT    std_logic;
	out210                               :   OUT    std_logic;
	out211                               :   OUT    std_logic;
	out212                               :   OUT    std_logic;
	out213                               :   OUT    std_logic;
	out214                               :   OUT    std_logic;
	out215                               :   OUT    std_logic;
	out216                               :   OUT    std_logic;
	out217                               :   OUT    std_logic;
	out218                               :   OUT    std_logic;
	out219                               :   OUT    std_logic;
	out220                               :   OUT    std_logic;
	out221                               :   OUT    std_logic;
	out222                               :   OUT    std_logic;
	out223                               :   OUT    std_logic;
	out224                               :   OUT    std_logic;
	out225                               :   OUT    std_logic;
	out226                               :   OUT    std_logic;
	out227                               :   OUT    std_logic;
	out228                               :   OUT    std_logic;
	out229                               :   OUT    std_logic;
	out230                               :   OUT    std_logic;
	out231                               :   OUT    std_logic;
	out232                               :   OUT    std_logic;
	out233                               :   OUT    std_logic;
	out234                               :   OUT    std_logic;
	out235                               :   OUT    std_logic;
	out236                               :   OUT    std_logic;
	out237                               :   OUT    std_logic;
	out238                               :   OUT    std_logic;
	out239                               :   OUT    std_logic;
	out240                               :   OUT    std_logic;
	out241                               :   OUT    std_logic;
	out242                               :   OUT    std_logic;
	out243                               :   OUT    std_logic;
	out244                               :   OUT    std_logic;
	out245                               :   OUT    std_logic;
	out246                               :   OUT    std_logic;
	out247                               :   OUT    std_logic;
	out248                               :   OUT    std_logic;
	out249                               :   OUT    std_logic;
	out250                               :   OUT    std_logic;
	out251                               :   OUT    std_logic;
	out252                               :   OUT    std_logic;
	out253                               :   OUT    std_logic;
	out254                               :   OUT    std_logic;
	out255                               :   OUT    std_logic;
	out256                               :   OUT    std_logic
	);
END encoderN256;

ARCHITECTURE rtl OF encoderN256 IS

  SIGNAL Logical_Operator_out1_out1            : std_logic;
  SIGNAL Logical_Operator_out2_out1            : std_logic;
  SIGNAL Logical_Operator_out3_out1            : std_logic;
  SIGNAL Logical_Operator_out4_out1            : std_logic;
  SIGNAL Logical_Operator_out5_out1            : std_logic;
  SIGNAL Logical_Operator_out6_out1            : std_logic;
  SIGNAL Logical_Operator_out7_out1            : std_logic;
  SIGNAL Logical_Operator_out8_out1            : std_logic;
  SIGNAL Logical_Operator_out9_out1            : std_logic;
  SIGNAL Logical_Operator_out10_out1            : std_logic;
  SIGNAL Logical_Operator_out11_out1            : std_logic;
  SIGNAL Logical_Operator_out12_out1            : std_logic;
  SIGNAL Logical_Operator_out13_out1            : std_logic;
  SIGNAL Logical_Operator_out14_out1            : std_logic;
  SIGNAL Logical_Operator_out15_out1            : std_logic;
  SIGNAL Logical_Operator_out16_out1            : std_logic;
  SIGNAL Logical_Operator_out17_out1            : std_logic;
  SIGNAL Logical_Operator_out18_out1            : std_logic;
  SIGNAL Logical_Operator_out19_out1            : std_logic;
  SIGNAL Logical_Operator_out20_out1            : std_logic;
  SIGNAL Logical_Operator_out21_out1            : std_logic;
  SIGNAL Logical_Operator_out22_out1            : std_logic;
  SIGNAL Logical_Operator_out23_out1            : std_logic;
  SIGNAL Logical_Operator_out24_out1            : std_logic;
  SIGNAL Logical_Operator_out25_out1            : std_logic;
  SIGNAL Logical_Operator_out26_out1            : std_logic;
  SIGNAL Logical_Operator_out27_out1            : std_logic;
  SIGNAL Logical_Operator_out28_out1            : std_logic;
  SIGNAL Logical_Operator_out29_out1            : std_logic;
  SIGNAL Logical_Operator_out30_out1            : std_logic;
  SIGNAL Logical_Operator_out31_out1            : std_logic;
  SIGNAL Logical_Operator_out32_out1            : std_logic;
  SIGNAL Logical_Operator_out33_out1            : std_logic;
  SIGNAL Logical_Operator_out34_out1            : std_logic;
  SIGNAL Logical_Operator_out35_out1            : std_logic;
  SIGNAL Logical_Operator_out36_out1            : std_logic;
  SIGNAL Logical_Operator_out37_out1            : std_logic;
  SIGNAL Logical_Operator_out38_out1            : std_logic;
  SIGNAL Logical_Operator_out39_out1            : std_logic;
  SIGNAL Logical_Operator_out40_out1            : std_logic;
  SIGNAL Logical_Operator_out41_out1            : std_logic;
  SIGNAL Logical_Operator_out42_out1            : std_logic;
  SIGNAL Logical_Operator_out43_out1            : std_logic;
  SIGNAL Logical_Operator_out44_out1            : std_logic;
  SIGNAL Logical_Operator_out45_out1            : std_logic;
  SIGNAL Logical_Operator_out46_out1            : std_logic;
  SIGNAL Logical_Operator_out47_out1            : std_logic;
  SIGNAL Logical_Operator_out48_out1            : std_logic;
  SIGNAL Logical_Operator_out49_out1            : std_logic;
  SIGNAL Logical_Operator_out50_out1            : std_logic;
  SIGNAL Logical_Operator_out51_out1            : std_logic;
  SIGNAL Logical_Operator_out52_out1            : std_logic;
  SIGNAL Logical_Operator_out53_out1            : std_logic;
  SIGNAL Logical_Operator_out54_out1            : std_logic;
  SIGNAL Logical_Operator_out55_out1            : std_logic;
  SIGNAL Logical_Operator_out56_out1            : std_logic;
  SIGNAL Logical_Operator_out57_out1            : std_logic;
  SIGNAL Logical_Operator_out58_out1            : std_logic;
  SIGNAL Logical_Operator_out59_out1            : std_logic;
  SIGNAL Logical_Operator_out60_out1            : std_logic;
  SIGNAL Logical_Operator_out61_out1            : std_logic;
  SIGNAL Logical_Operator_out62_out1            : std_logic;
  SIGNAL Logical_Operator_out63_out1            : std_logic;
  SIGNAL Logical_Operator_out64_out1            : std_logic;
  SIGNAL Logical_Operator_out65_out1            : std_logic;
  SIGNAL Logical_Operator_out66_out1            : std_logic;
  SIGNAL Logical_Operator_out67_out1            : std_logic;
  SIGNAL Logical_Operator_out68_out1            : std_logic;
  SIGNAL Logical_Operator_out69_out1            : std_logic;
  SIGNAL Logical_Operator_out70_out1            : std_logic;
  SIGNAL Logical_Operator_out71_out1            : std_logic;
  SIGNAL Logical_Operator_out72_out1            : std_logic;
  SIGNAL Logical_Operator_out73_out1            : std_logic;
  SIGNAL Logical_Operator_out74_out1            : std_logic;
  SIGNAL Logical_Operator_out75_out1            : std_logic;
  SIGNAL Logical_Operator_out76_out1            : std_logic;
  SIGNAL Logical_Operator_out77_out1            : std_logic;
  SIGNAL Logical_Operator_out78_out1            : std_logic;
  SIGNAL Logical_Operator_out79_out1            : std_logic;
  SIGNAL Logical_Operator_out80_out1            : std_logic;
  SIGNAL Logical_Operator_out81_out1            : std_logic;
  SIGNAL Logical_Operator_out82_out1            : std_logic;
  SIGNAL Logical_Operator_out83_out1            : std_logic;
  SIGNAL Logical_Operator_out84_out1            : std_logic;
  SIGNAL Logical_Operator_out85_out1            : std_logic;
  SIGNAL Logical_Operator_out86_out1            : std_logic;
  SIGNAL Logical_Operator_out87_out1            : std_logic;
  SIGNAL Logical_Operator_out88_out1            : std_logic;
  SIGNAL Logical_Operator_out89_out1            : std_logic;
  SIGNAL Logical_Operator_out90_out1            : std_logic;
  SIGNAL Logical_Operator_out91_out1            : std_logic;
  SIGNAL Logical_Operator_out92_out1            : std_logic;
  SIGNAL Logical_Operator_out93_out1            : std_logic;
  SIGNAL Logical_Operator_out94_out1            : std_logic;
  SIGNAL Logical_Operator_out95_out1            : std_logic;
  SIGNAL Logical_Operator_out96_out1            : std_logic;
  SIGNAL Logical_Operator_out97_out1            : std_logic;
  SIGNAL Logical_Operator_out98_out1            : std_logic;
  SIGNAL Logical_Operator_out99_out1            : std_logic;
  SIGNAL Logical_Operator_out100_out1            : std_logic;
  SIGNAL Logical_Operator_out101_out1            : std_logic;
  SIGNAL Logical_Operator_out102_out1            : std_logic;
  SIGNAL Logical_Operator_out103_out1            : std_logic;
  SIGNAL Logical_Operator_out104_out1            : std_logic;
  SIGNAL Logical_Operator_out105_out1            : std_logic;
  SIGNAL Logical_Operator_out106_out1            : std_logic;
  SIGNAL Logical_Operator_out107_out1            : std_logic;
  SIGNAL Logical_Operator_out108_out1            : std_logic;
  SIGNAL Logical_Operator_out109_out1            : std_logic;
  SIGNAL Logical_Operator_out110_out1            : std_logic;
  SIGNAL Logical_Operator_out111_out1            : std_logic;
  SIGNAL Logical_Operator_out112_out1            : std_logic;
  SIGNAL Logical_Operator_out113_out1            : std_logic;
  SIGNAL Logical_Operator_out114_out1            : std_logic;
  SIGNAL Logical_Operator_out115_out1            : std_logic;
  SIGNAL Logical_Operator_out116_out1            : std_logic;
  SIGNAL Logical_Operator_out117_out1            : std_logic;
  SIGNAL Logical_Operator_out118_out1            : std_logic;
  SIGNAL Logical_Operator_out119_out1            : std_logic;
  SIGNAL Logical_Operator_out120_out1            : std_logic;
  SIGNAL Logical_Operator_out121_out1            : std_logic;
  SIGNAL Logical_Operator_out122_out1            : std_logic;
  SIGNAL Logical_Operator_out123_out1            : std_logic;
  SIGNAL Logical_Operator_out124_out1            : std_logic;
  SIGNAL Logical_Operator_out125_out1            : std_logic;
  SIGNAL Logical_Operator_out126_out1            : std_logic;
  SIGNAL Logical_Operator_out127_out1            : std_logic;
  SIGNAL Logical_Operator_out128_out1            : std_logic;
  SIGNAL Logical_Operator_out129_out1            : std_logic;
  SIGNAL Logical_Operator_out130_out1            : std_logic;
  SIGNAL Logical_Operator_out131_out1            : std_logic;
  SIGNAL Logical_Operator_out132_out1            : std_logic;
  SIGNAL Logical_Operator_out133_out1            : std_logic;
  SIGNAL Logical_Operator_out134_out1            : std_logic;
  SIGNAL Logical_Operator_out135_out1            : std_logic;
  SIGNAL Logical_Operator_out136_out1            : std_logic;
  SIGNAL Logical_Operator_out137_out1            : std_logic;
  SIGNAL Logical_Operator_out138_out1            : std_logic;
  SIGNAL Logical_Operator_out139_out1            : std_logic;
  SIGNAL Logical_Operator_out140_out1            : std_logic;
  SIGNAL Logical_Operator_out141_out1            : std_logic;
  SIGNAL Logical_Operator_out142_out1            : std_logic;
  SIGNAL Logical_Operator_out143_out1            : std_logic;
  SIGNAL Logical_Operator_out144_out1            : std_logic;
  SIGNAL Logical_Operator_out145_out1            : std_logic;
  SIGNAL Logical_Operator_out146_out1            : std_logic;
  SIGNAL Logical_Operator_out147_out1            : std_logic;
  SIGNAL Logical_Operator_out148_out1            : std_logic;
  SIGNAL Logical_Operator_out149_out1            : std_logic;
  SIGNAL Logical_Operator_out150_out1            : std_logic;
  SIGNAL Logical_Operator_out151_out1            : std_logic;
  SIGNAL Logical_Operator_out152_out1            : std_logic;
  SIGNAL Logical_Operator_out153_out1            : std_logic;
  SIGNAL Logical_Operator_out154_out1            : std_logic;
  SIGNAL Logical_Operator_out155_out1            : std_logic;
  SIGNAL Logical_Operator_out156_out1            : std_logic;
  SIGNAL Logical_Operator_out157_out1            : std_logic;
  SIGNAL Logical_Operator_out158_out1            : std_logic;
  SIGNAL Logical_Operator_out159_out1            : std_logic;
  SIGNAL Logical_Operator_out160_out1            : std_logic;
  SIGNAL Logical_Operator_out161_out1            : std_logic;
  SIGNAL Logical_Operator_out162_out1            : std_logic;
  SIGNAL Logical_Operator_out163_out1            : std_logic;
  SIGNAL Logical_Operator_out164_out1            : std_logic;
  SIGNAL Logical_Operator_out165_out1            : std_logic;
  SIGNAL Logical_Operator_out166_out1            : std_logic;
  SIGNAL Logical_Operator_out167_out1            : std_logic;
  SIGNAL Logical_Operator_out168_out1            : std_logic;
  SIGNAL Logical_Operator_out169_out1            : std_logic;
  SIGNAL Logical_Operator_out170_out1            : std_logic;
  SIGNAL Logical_Operator_out171_out1            : std_logic;
  SIGNAL Logical_Operator_out172_out1            : std_logic;
  SIGNAL Logical_Operator_out173_out1            : std_logic;
  SIGNAL Logical_Operator_out174_out1            : std_logic;
  SIGNAL Logical_Operator_out175_out1            : std_logic;
  SIGNAL Logical_Operator_out176_out1            : std_logic;
  SIGNAL Logical_Operator_out177_out1            : std_logic;
  SIGNAL Logical_Operator_out178_out1            : std_logic;
  SIGNAL Logical_Operator_out179_out1            : std_logic;
  SIGNAL Logical_Operator_out180_out1            : std_logic;
  SIGNAL Logical_Operator_out181_out1            : std_logic;
  SIGNAL Logical_Operator_out182_out1            : std_logic;
  SIGNAL Logical_Operator_out183_out1            : std_logic;
  SIGNAL Logical_Operator_out184_out1            : std_logic;
  SIGNAL Logical_Operator_out185_out1            : std_logic;
  SIGNAL Logical_Operator_out186_out1            : std_logic;
  SIGNAL Logical_Operator_out187_out1            : std_logic;
  SIGNAL Logical_Operator_out188_out1            : std_logic;
  SIGNAL Logical_Operator_out189_out1            : std_logic;
  SIGNAL Logical_Operator_out190_out1            : std_logic;
  SIGNAL Logical_Operator_out191_out1            : std_logic;
  SIGNAL Logical_Operator_out192_out1            : std_logic;
  SIGNAL Logical_Operator_out193_out1            : std_logic;
  SIGNAL Logical_Operator_out194_out1            : std_logic;
  SIGNAL Logical_Operator_out195_out1            : std_logic;
  SIGNAL Logical_Operator_out196_out1            : std_logic;
  SIGNAL Logical_Operator_out197_out1            : std_logic;
  SIGNAL Logical_Operator_out198_out1            : std_logic;
  SIGNAL Logical_Operator_out199_out1            : std_logic;
  SIGNAL Logical_Operator_out200_out1            : std_logic;
  SIGNAL Logical_Operator_out201_out1            : std_logic;
  SIGNAL Logical_Operator_out202_out1            : std_logic;
  SIGNAL Logical_Operator_out203_out1            : std_logic;
  SIGNAL Logical_Operator_out204_out1            : std_logic;
  SIGNAL Logical_Operator_out205_out1            : std_logic;
  SIGNAL Logical_Operator_out206_out1            : std_logic;
  SIGNAL Logical_Operator_out207_out1            : std_logic;
  SIGNAL Logical_Operator_out208_out1            : std_logic;
  SIGNAL Logical_Operator_out209_out1            : std_logic;
  SIGNAL Logical_Operator_out210_out1            : std_logic;
  SIGNAL Logical_Operator_out211_out1            : std_logic;
  SIGNAL Logical_Operator_out212_out1            : std_logic;
  SIGNAL Logical_Operator_out213_out1            : std_logic;
  SIGNAL Logical_Operator_out214_out1            : std_logic;
  SIGNAL Logical_Operator_out215_out1            : std_logic;
  SIGNAL Logical_Operator_out216_out1            : std_logic;
  SIGNAL Logical_Operator_out217_out1            : std_logic;
  SIGNAL Logical_Operator_out218_out1            : std_logic;
  SIGNAL Logical_Operator_out219_out1            : std_logic;
  SIGNAL Logical_Operator_out220_out1            : std_logic;
  SIGNAL Logical_Operator_out221_out1            : std_logic;
  SIGNAL Logical_Operator_out222_out1            : std_logic;
  SIGNAL Logical_Operator_out223_out1            : std_logic;
  SIGNAL Logical_Operator_out224_out1            : std_logic;
  SIGNAL Logical_Operator_out225_out1            : std_logic;
  SIGNAL Logical_Operator_out226_out1            : std_logic;
  SIGNAL Logical_Operator_out227_out1            : std_logic;
  SIGNAL Logical_Operator_out228_out1            : std_logic;
  SIGNAL Logical_Operator_out229_out1            : std_logic;
  SIGNAL Logical_Operator_out230_out1            : std_logic;
  SIGNAL Logical_Operator_out231_out1            : std_logic;
  SIGNAL Logical_Operator_out232_out1            : std_logic;
  SIGNAL Logical_Operator_out233_out1            : std_logic;
  SIGNAL Logical_Operator_out234_out1            : std_logic;
  SIGNAL Logical_Operator_out235_out1            : std_logic;
  SIGNAL Logical_Operator_out236_out1            : std_logic;
  SIGNAL Logical_Operator_out237_out1            : std_logic;
  SIGNAL Logical_Operator_out238_out1            : std_logic;
  SIGNAL Logical_Operator_out239_out1            : std_logic;
  SIGNAL Logical_Operator_out240_out1            : std_logic;
  SIGNAL Logical_Operator_out241_out1            : std_logic;
  SIGNAL Logical_Operator_out242_out1            : std_logic;
  SIGNAL Logical_Operator_out243_out1            : std_logic;
  SIGNAL Logical_Operator_out244_out1            : std_logic;
  SIGNAL Logical_Operator_out245_out1            : std_logic;
  SIGNAL Logical_Operator_out246_out1            : std_logic;
  SIGNAL Logical_Operator_out247_out1            : std_logic;
  SIGNAL Logical_Operator_out248_out1            : std_logic;
  SIGNAL Logical_Operator_out249_out1            : std_logic;
  SIGNAL Logical_Operator_out250_out1            : std_logic;
  SIGNAL Logical_Operator_out251_out1            : std_logic;
  SIGNAL Logical_Operator_out252_out1            : std_logic;
  SIGNAL Logical_Operator_out253_out1            : std_logic;
  SIGNAL Logical_Operator_out254_out1            : std_logic;
  SIGNAL Logical_Operator_out255_out1            : std_logic;
  SIGNAL Logical_Operator_out256_out1            : std_logic;
  SIGNAL Logical_Operator_out257_out1            : std_logic;
  SIGNAL Logical_Operator_out258_out1            : std_logic;
  SIGNAL Logical_Operator_out259_out1            : std_logic;
  SIGNAL Logical_Operator_out260_out1            : std_logic;
  SIGNAL Logical_Operator_out261_out1            : std_logic;
  SIGNAL Logical_Operator_out262_out1            : std_logic;
  SIGNAL Logical_Operator_out263_out1            : std_logic;
  SIGNAL Logical_Operator_out264_out1            : std_logic;
  SIGNAL Logical_Operator_out265_out1            : std_logic;
  SIGNAL Logical_Operator_out266_out1            : std_logic;
  SIGNAL Logical_Operator_out267_out1            : std_logic;
  SIGNAL Logical_Operator_out268_out1            : std_logic;
  SIGNAL Logical_Operator_out269_out1            : std_logic;
  SIGNAL Logical_Operator_out270_out1            : std_logic;
  SIGNAL Logical_Operator_out271_out1            : std_logic;
  SIGNAL Logical_Operator_out272_out1            : std_logic;
  SIGNAL Logical_Operator_out273_out1            : std_logic;
  SIGNAL Logical_Operator_out274_out1            : std_logic;
  SIGNAL Logical_Operator_out275_out1            : std_logic;
  SIGNAL Logical_Operator_out276_out1            : std_logic;
  SIGNAL Logical_Operator_out277_out1            : std_logic;
  SIGNAL Logical_Operator_out278_out1            : std_logic;
  SIGNAL Logical_Operator_out279_out1            : std_logic;
  SIGNAL Logical_Operator_out280_out1            : std_logic;
  SIGNAL Logical_Operator_out281_out1            : std_logic;
  SIGNAL Logical_Operator_out282_out1            : std_logic;
  SIGNAL Logical_Operator_out283_out1            : std_logic;
  SIGNAL Logical_Operator_out284_out1            : std_logic;
  SIGNAL Logical_Operator_out285_out1            : std_logic;
  SIGNAL Logical_Operator_out286_out1            : std_logic;
  SIGNAL Logical_Operator_out287_out1            : std_logic;
  SIGNAL Logical_Operator_out288_out1            : std_logic;
  SIGNAL Logical_Operator_out289_out1            : std_logic;
  SIGNAL Logical_Operator_out290_out1            : std_logic;
  SIGNAL Logical_Operator_out291_out1            : std_logic;
  SIGNAL Logical_Operator_out292_out1            : std_logic;
  SIGNAL Logical_Operator_out293_out1            : std_logic;
  SIGNAL Logical_Operator_out294_out1            : std_logic;
  SIGNAL Logical_Operator_out295_out1            : std_logic;
  SIGNAL Logical_Operator_out296_out1            : std_logic;
  SIGNAL Logical_Operator_out297_out1            : std_logic;
  SIGNAL Logical_Operator_out298_out1            : std_logic;
  SIGNAL Logical_Operator_out299_out1            : std_logic;
  SIGNAL Logical_Operator_out300_out1            : std_logic;
  SIGNAL Logical_Operator_out301_out1            : std_logic;
  SIGNAL Logical_Operator_out302_out1            : std_logic;
  SIGNAL Logical_Operator_out303_out1            : std_logic;
  SIGNAL Logical_Operator_out304_out1            : std_logic;
  SIGNAL Logical_Operator_out305_out1            : std_logic;
  SIGNAL Logical_Operator_out306_out1            : std_logic;
  SIGNAL Logical_Operator_out307_out1            : std_logic;
  SIGNAL Logical_Operator_out308_out1            : std_logic;
  SIGNAL Logical_Operator_out309_out1            : std_logic;
  SIGNAL Logical_Operator_out310_out1            : std_logic;
  SIGNAL Logical_Operator_out311_out1            : std_logic;
  SIGNAL Logical_Operator_out312_out1            : std_logic;
  SIGNAL Logical_Operator_out313_out1            : std_logic;
  SIGNAL Logical_Operator_out314_out1            : std_logic;
  SIGNAL Logical_Operator_out315_out1            : std_logic;
  SIGNAL Logical_Operator_out316_out1            : std_logic;
  SIGNAL Logical_Operator_out317_out1            : std_logic;
  SIGNAL Logical_Operator_out318_out1            : std_logic;
  SIGNAL Logical_Operator_out319_out1            : std_logic;
  SIGNAL Logical_Operator_out320_out1            : std_logic;
  SIGNAL Logical_Operator_out321_out1            : std_logic;
  SIGNAL Logical_Operator_out322_out1            : std_logic;
  SIGNAL Logical_Operator_out323_out1            : std_logic;
  SIGNAL Logical_Operator_out324_out1            : std_logic;
  SIGNAL Logical_Operator_out325_out1            : std_logic;
  SIGNAL Logical_Operator_out326_out1            : std_logic;
  SIGNAL Logical_Operator_out327_out1            : std_logic;
  SIGNAL Logical_Operator_out328_out1            : std_logic;
  SIGNAL Logical_Operator_out329_out1            : std_logic;
  SIGNAL Logical_Operator_out330_out1            : std_logic;
  SIGNAL Logical_Operator_out331_out1            : std_logic;
  SIGNAL Logical_Operator_out332_out1            : std_logic;
  SIGNAL Logical_Operator_out333_out1            : std_logic;
  SIGNAL Logical_Operator_out334_out1            : std_logic;
  SIGNAL Logical_Operator_out335_out1            : std_logic;
  SIGNAL Logical_Operator_out336_out1            : std_logic;
  SIGNAL Logical_Operator_out337_out1            : std_logic;
  SIGNAL Logical_Operator_out338_out1            : std_logic;
  SIGNAL Logical_Operator_out339_out1            : std_logic;
  SIGNAL Logical_Operator_out340_out1            : std_logic;
  SIGNAL Logical_Operator_out341_out1            : std_logic;
  SIGNAL Logical_Operator_out342_out1            : std_logic;
  SIGNAL Logical_Operator_out343_out1            : std_logic;
  SIGNAL Logical_Operator_out344_out1            : std_logic;
  SIGNAL Logical_Operator_out345_out1            : std_logic;
  SIGNAL Logical_Operator_out346_out1            : std_logic;
  SIGNAL Logical_Operator_out347_out1            : std_logic;
  SIGNAL Logical_Operator_out348_out1            : std_logic;
  SIGNAL Logical_Operator_out349_out1            : std_logic;
  SIGNAL Logical_Operator_out350_out1            : std_logic;
  SIGNAL Logical_Operator_out351_out1            : std_logic;
  SIGNAL Logical_Operator_out352_out1            : std_logic;
  SIGNAL Logical_Operator_out353_out1            : std_logic;
  SIGNAL Logical_Operator_out354_out1            : std_logic;
  SIGNAL Logical_Operator_out355_out1            : std_logic;
  SIGNAL Logical_Operator_out356_out1            : std_logic;
  SIGNAL Logical_Operator_out357_out1            : std_logic;
  SIGNAL Logical_Operator_out358_out1            : std_logic;
  SIGNAL Logical_Operator_out359_out1            : std_logic;
  SIGNAL Logical_Operator_out360_out1            : std_logic;
  SIGNAL Logical_Operator_out361_out1            : std_logic;
  SIGNAL Logical_Operator_out362_out1            : std_logic;
  SIGNAL Logical_Operator_out363_out1            : std_logic;
  SIGNAL Logical_Operator_out364_out1            : std_logic;
  SIGNAL Logical_Operator_out365_out1            : std_logic;
  SIGNAL Logical_Operator_out366_out1            : std_logic;
  SIGNAL Logical_Operator_out367_out1            : std_logic;
  SIGNAL Logical_Operator_out368_out1            : std_logic;
  SIGNAL Logical_Operator_out369_out1            : std_logic;
  SIGNAL Logical_Operator_out370_out1            : std_logic;
  SIGNAL Logical_Operator_out371_out1            : std_logic;
  SIGNAL Logical_Operator_out372_out1            : std_logic;
  SIGNAL Logical_Operator_out373_out1            : std_logic;
  SIGNAL Logical_Operator_out374_out1            : std_logic;
  SIGNAL Logical_Operator_out375_out1            : std_logic;
  SIGNAL Logical_Operator_out376_out1            : std_logic;
  SIGNAL Logical_Operator_out377_out1            : std_logic;
  SIGNAL Logical_Operator_out378_out1            : std_logic;
  SIGNAL Logical_Operator_out379_out1            : std_logic;
  SIGNAL Logical_Operator_out380_out1            : std_logic;
  SIGNAL Logical_Operator_out381_out1            : std_logic;
  SIGNAL Logical_Operator_out382_out1            : std_logic;
  SIGNAL Logical_Operator_out383_out1            : std_logic;
  SIGNAL Logical_Operator_out384_out1            : std_logic;
  SIGNAL Logical_Operator_out385_out1            : std_logic;
  SIGNAL Logical_Operator_out386_out1            : std_logic;
  SIGNAL Logical_Operator_out387_out1            : std_logic;
  SIGNAL Logical_Operator_out388_out1            : std_logic;
  SIGNAL Logical_Operator_out389_out1            : std_logic;
  SIGNAL Logical_Operator_out390_out1            : std_logic;
  SIGNAL Logical_Operator_out391_out1            : std_logic;
  SIGNAL Logical_Operator_out392_out1            : std_logic;
  SIGNAL Logical_Operator_out393_out1            : std_logic;
  SIGNAL Logical_Operator_out394_out1            : std_logic;
  SIGNAL Logical_Operator_out395_out1            : std_logic;
  SIGNAL Logical_Operator_out396_out1            : std_logic;
  SIGNAL Logical_Operator_out397_out1            : std_logic;
  SIGNAL Logical_Operator_out398_out1            : std_logic;
  SIGNAL Logical_Operator_out399_out1            : std_logic;
  SIGNAL Logical_Operator_out400_out1            : std_logic;
  SIGNAL Logical_Operator_out401_out1            : std_logic;
  SIGNAL Logical_Operator_out402_out1            : std_logic;
  SIGNAL Logical_Operator_out403_out1            : std_logic;
  SIGNAL Logical_Operator_out404_out1            : std_logic;
  SIGNAL Logical_Operator_out405_out1            : std_logic;
  SIGNAL Logical_Operator_out406_out1            : std_logic;
  SIGNAL Logical_Operator_out407_out1            : std_logic;
  SIGNAL Logical_Operator_out408_out1            : std_logic;
  SIGNAL Logical_Operator_out409_out1            : std_logic;
  SIGNAL Logical_Operator_out410_out1            : std_logic;
  SIGNAL Logical_Operator_out411_out1            : std_logic;
  SIGNAL Logical_Operator_out412_out1            : std_logic;
  SIGNAL Logical_Operator_out413_out1            : std_logic;
  SIGNAL Logical_Operator_out414_out1            : std_logic;
  SIGNAL Logical_Operator_out415_out1            : std_logic;
  SIGNAL Logical_Operator_out416_out1            : std_logic;
  SIGNAL Logical_Operator_out417_out1            : std_logic;
  SIGNAL Logical_Operator_out418_out1            : std_logic;
  SIGNAL Logical_Operator_out419_out1            : std_logic;
  SIGNAL Logical_Operator_out420_out1            : std_logic;
  SIGNAL Logical_Operator_out421_out1            : std_logic;
  SIGNAL Logical_Operator_out422_out1            : std_logic;
  SIGNAL Logical_Operator_out423_out1            : std_logic;
  SIGNAL Logical_Operator_out424_out1            : std_logic;
  SIGNAL Logical_Operator_out425_out1            : std_logic;
  SIGNAL Logical_Operator_out426_out1            : std_logic;
  SIGNAL Logical_Operator_out427_out1            : std_logic;
  SIGNAL Logical_Operator_out428_out1            : std_logic;
  SIGNAL Logical_Operator_out429_out1            : std_logic;
  SIGNAL Logical_Operator_out430_out1            : std_logic;
  SIGNAL Logical_Operator_out431_out1            : std_logic;
  SIGNAL Logical_Operator_out432_out1            : std_logic;
  SIGNAL Logical_Operator_out433_out1            : std_logic;
  SIGNAL Logical_Operator_out434_out1            : std_logic;
  SIGNAL Logical_Operator_out435_out1            : std_logic;
  SIGNAL Logical_Operator_out436_out1            : std_logic;
  SIGNAL Logical_Operator_out437_out1            : std_logic;
  SIGNAL Logical_Operator_out438_out1            : std_logic;
  SIGNAL Logical_Operator_out439_out1            : std_logic;
  SIGNAL Logical_Operator_out440_out1            : std_logic;
  SIGNAL Logical_Operator_out441_out1            : std_logic;
  SIGNAL Logical_Operator_out442_out1            : std_logic;
  SIGNAL Logical_Operator_out443_out1            : std_logic;
  SIGNAL Logical_Operator_out444_out1            : std_logic;
  SIGNAL Logical_Operator_out445_out1            : std_logic;
  SIGNAL Logical_Operator_out446_out1            : std_logic;
  SIGNAL Logical_Operator_out447_out1            : std_logic;
  SIGNAL Logical_Operator_out448_out1            : std_logic;
  SIGNAL Logical_Operator_out449_out1            : std_logic;
  SIGNAL Logical_Operator_out450_out1            : std_logic;
  SIGNAL Logical_Operator_out451_out1            : std_logic;
  SIGNAL Logical_Operator_out452_out1            : std_logic;
  SIGNAL Logical_Operator_out453_out1            : std_logic;
  SIGNAL Logical_Operator_out454_out1            : std_logic;
  SIGNAL Logical_Operator_out455_out1            : std_logic;
  SIGNAL Logical_Operator_out456_out1            : std_logic;
  SIGNAL Logical_Operator_out457_out1            : std_logic;
  SIGNAL Logical_Operator_out458_out1            : std_logic;
  SIGNAL Logical_Operator_out459_out1            : std_logic;
  SIGNAL Logical_Operator_out460_out1            : std_logic;
  SIGNAL Logical_Operator_out461_out1            : std_logic;
  SIGNAL Logical_Operator_out462_out1            : std_logic;
  SIGNAL Logical_Operator_out463_out1            : std_logic;
  SIGNAL Logical_Operator_out464_out1            : std_logic;
  SIGNAL Logical_Operator_out465_out1            : std_logic;
  SIGNAL Logical_Operator_out466_out1            : std_logic;
  SIGNAL Logical_Operator_out467_out1            : std_logic;
  SIGNAL Logical_Operator_out468_out1            : std_logic;
  SIGNAL Logical_Operator_out469_out1            : std_logic;
  SIGNAL Logical_Operator_out470_out1            : std_logic;
  SIGNAL Logical_Operator_out471_out1            : std_logic;
  SIGNAL Logical_Operator_out472_out1            : std_logic;
  SIGNAL Logical_Operator_out473_out1            : std_logic;
  SIGNAL Logical_Operator_out474_out1            : std_logic;
  SIGNAL Logical_Operator_out475_out1            : std_logic;
  SIGNAL Logical_Operator_out476_out1            : std_logic;
  SIGNAL Logical_Operator_out477_out1            : std_logic;
  SIGNAL Logical_Operator_out478_out1            : std_logic;
  SIGNAL Logical_Operator_out479_out1            : std_logic;
  SIGNAL Logical_Operator_out480_out1            : std_logic;
  SIGNAL Logical_Operator_out481_out1            : std_logic;
  SIGNAL Logical_Operator_out482_out1            : std_logic;
  SIGNAL Logical_Operator_out483_out1            : std_logic;
  SIGNAL Logical_Operator_out484_out1            : std_logic;
  SIGNAL Logical_Operator_out485_out1            : std_logic;
  SIGNAL Logical_Operator_out486_out1            : std_logic;
  SIGNAL Logical_Operator_out487_out1            : std_logic;
  SIGNAL Logical_Operator_out488_out1            : std_logic;
  SIGNAL Logical_Operator_out489_out1            : std_logic;
  SIGNAL Logical_Operator_out490_out1            : std_logic;
  SIGNAL Logical_Operator_out491_out1            : std_logic;
  SIGNAL Logical_Operator_out492_out1            : std_logic;
  SIGNAL Logical_Operator_out493_out1            : std_logic;
  SIGNAL Logical_Operator_out494_out1            : std_logic;
  SIGNAL Logical_Operator_out495_out1            : std_logic;
  SIGNAL Logical_Operator_out496_out1            : std_logic;
  SIGNAL Logical_Operator_out497_out1            : std_logic;
  SIGNAL Logical_Operator_out498_out1            : std_logic;
  SIGNAL Logical_Operator_out499_out1            : std_logic;
  SIGNAL Logical_Operator_out500_out1            : std_logic;
  SIGNAL Logical_Operator_out501_out1            : std_logic;
  SIGNAL Logical_Operator_out502_out1            : std_logic;
  SIGNAL Logical_Operator_out503_out1            : std_logic;
  SIGNAL Logical_Operator_out504_out1            : std_logic;
  SIGNAL Logical_Operator_out505_out1            : std_logic;
  SIGNAL Logical_Operator_out506_out1            : std_logic;
  SIGNAL Logical_Operator_out507_out1            : std_logic;
  SIGNAL Logical_Operator_out508_out1            : std_logic;
  SIGNAL Logical_Operator_out509_out1            : std_logic;
  SIGNAL Logical_Operator_out510_out1            : std_logic;
  SIGNAL Logical_Operator_out511_out1            : std_logic;
  SIGNAL Logical_Operator_out512_out1            : std_logic;
  SIGNAL Logical_Operator_out513_out1            : std_logic;
  SIGNAL Logical_Operator_out514_out1            : std_logic;
  SIGNAL Logical_Operator_out515_out1            : std_logic;
  SIGNAL Logical_Operator_out516_out1            : std_logic;
  SIGNAL Logical_Operator_out517_out1            : std_logic;
  SIGNAL Logical_Operator_out518_out1            : std_logic;
  SIGNAL Logical_Operator_out519_out1            : std_logic;
  SIGNAL Logical_Operator_out520_out1            : std_logic;
  SIGNAL Logical_Operator_out521_out1            : std_logic;
  SIGNAL Logical_Operator_out522_out1            : std_logic;
  SIGNAL Logical_Operator_out523_out1            : std_logic;
  SIGNAL Logical_Operator_out524_out1            : std_logic;
  SIGNAL Logical_Operator_out525_out1            : std_logic;
  SIGNAL Logical_Operator_out526_out1            : std_logic;
  SIGNAL Logical_Operator_out527_out1            : std_logic;
  SIGNAL Logical_Operator_out528_out1            : std_logic;
  SIGNAL Logical_Operator_out529_out1            : std_logic;
  SIGNAL Logical_Operator_out530_out1            : std_logic;
  SIGNAL Logical_Operator_out531_out1            : std_logic;
  SIGNAL Logical_Operator_out532_out1            : std_logic;
  SIGNAL Logical_Operator_out533_out1            : std_logic;
  SIGNAL Logical_Operator_out534_out1            : std_logic;
  SIGNAL Logical_Operator_out535_out1            : std_logic;
  SIGNAL Logical_Operator_out536_out1            : std_logic;
  SIGNAL Logical_Operator_out537_out1            : std_logic;
  SIGNAL Logical_Operator_out538_out1            : std_logic;
  SIGNAL Logical_Operator_out539_out1            : std_logic;
  SIGNAL Logical_Operator_out540_out1            : std_logic;
  SIGNAL Logical_Operator_out541_out1            : std_logic;
  SIGNAL Logical_Operator_out542_out1            : std_logic;
  SIGNAL Logical_Operator_out543_out1            : std_logic;
  SIGNAL Logical_Operator_out544_out1            : std_logic;
  SIGNAL Logical_Operator_out545_out1            : std_logic;
  SIGNAL Logical_Operator_out546_out1            : std_logic;
  SIGNAL Logical_Operator_out547_out1            : std_logic;
  SIGNAL Logical_Operator_out548_out1            : std_logic;
  SIGNAL Logical_Operator_out549_out1            : std_logic;
  SIGNAL Logical_Operator_out550_out1            : std_logic;
  SIGNAL Logical_Operator_out551_out1            : std_logic;
  SIGNAL Logical_Operator_out552_out1            : std_logic;
  SIGNAL Logical_Operator_out553_out1            : std_logic;
  SIGNAL Logical_Operator_out554_out1            : std_logic;
  SIGNAL Logical_Operator_out555_out1            : std_logic;
  SIGNAL Logical_Operator_out556_out1            : std_logic;
  SIGNAL Logical_Operator_out557_out1            : std_logic;
  SIGNAL Logical_Operator_out558_out1            : std_logic;
  SIGNAL Logical_Operator_out559_out1            : std_logic;
  SIGNAL Logical_Operator_out560_out1            : std_logic;
  SIGNAL Logical_Operator_out561_out1            : std_logic;
  SIGNAL Logical_Operator_out562_out1            : std_logic;
  SIGNAL Logical_Operator_out563_out1            : std_logic;
  SIGNAL Logical_Operator_out564_out1            : std_logic;
  SIGNAL Logical_Operator_out565_out1            : std_logic;
  SIGNAL Logical_Operator_out566_out1            : std_logic;
  SIGNAL Logical_Operator_out567_out1            : std_logic;
  SIGNAL Logical_Operator_out568_out1            : std_logic;
  SIGNAL Logical_Operator_out569_out1            : std_logic;
  SIGNAL Logical_Operator_out570_out1            : std_logic;
  SIGNAL Logical_Operator_out571_out1            : std_logic;
  SIGNAL Logical_Operator_out572_out1            : std_logic;
  SIGNAL Logical_Operator_out573_out1            : std_logic;
  SIGNAL Logical_Operator_out574_out1            : std_logic;
  SIGNAL Logical_Operator_out575_out1            : std_logic;
  SIGNAL Logical_Operator_out576_out1            : std_logic;
  SIGNAL Logical_Operator_out577_out1            : std_logic;
  SIGNAL Logical_Operator_out578_out1            : std_logic;
  SIGNAL Logical_Operator_out579_out1            : std_logic;
  SIGNAL Logical_Operator_out580_out1            : std_logic;
  SIGNAL Logical_Operator_out581_out1            : std_logic;
  SIGNAL Logical_Operator_out582_out1            : std_logic;
  SIGNAL Logical_Operator_out583_out1            : std_logic;
  SIGNAL Logical_Operator_out584_out1            : std_logic;
  SIGNAL Logical_Operator_out585_out1            : std_logic;
  SIGNAL Logical_Operator_out586_out1            : std_logic;
  SIGNAL Logical_Operator_out587_out1            : std_logic;
  SIGNAL Logical_Operator_out588_out1            : std_logic;
  SIGNAL Logical_Operator_out589_out1            : std_logic;
  SIGNAL Logical_Operator_out590_out1            : std_logic;
  SIGNAL Logical_Operator_out591_out1            : std_logic;
  SIGNAL Logical_Operator_out592_out1            : std_logic;
  SIGNAL Logical_Operator_out593_out1            : std_logic;
  SIGNAL Logical_Operator_out594_out1            : std_logic;
  SIGNAL Logical_Operator_out595_out1            : std_logic;
  SIGNAL Logical_Operator_out596_out1            : std_logic;
  SIGNAL Logical_Operator_out597_out1            : std_logic;
  SIGNAL Logical_Operator_out598_out1            : std_logic;
  SIGNAL Logical_Operator_out599_out1            : std_logic;
  SIGNAL Logical_Operator_out600_out1            : std_logic;
  SIGNAL Logical_Operator_out601_out1            : std_logic;
  SIGNAL Logical_Operator_out602_out1            : std_logic;
  SIGNAL Logical_Operator_out603_out1            : std_logic;
  SIGNAL Logical_Operator_out604_out1            : std_logic;
  SIGNAL Logical_Operator_out605_out1            : std_logic;
  SIGNAL Logical_Operator_out606_out1            : std_logic;
  SIGNAL Logical_Operator_out607_out1            : std_logic;
  SIGNAL Logical_Operator_out608_out1            : std_logic;
  SIGNAL Logical_Operator_out609_out1            : std_logic;
  SIGNAL Logical_Operator_out610_out1            : std_logic;
  SIGNAL Logical_Operator_out611_out1            : std_logic;
  SIGNAL Logical_Operator_out612_out1            : std_logic;
  SIGNAL Logical_Operator_out613_out1            : std_logic;
  SIGNAL Logical_Operator_out614_out1            : std_logic;
  SIGNAL Logical_Operator_out615_out1            : std_logic;
  SIGNAL Logical_Operator_out616_out1            : std_logic;
  SIGNAL Logical_Operator_out617_out1            : std_logic;
  SIGNAL Logical_Operator_out618_out1            : std_logic;
  SIGNAL Logical_Operator_out619_out1            : std_logic;
  SIGNAL Logical_Operator_out620_out1            : std_logic;
  SIGNAL Logical_Operator_out621_out1            : std_logic;
  SIGNAL Logical_Operator_out622_out1            : std_logic;
  SIGNAL Logical_Operator_out623_out1            : std_logic;
  SIGNAL Logical_Operator_out624_out1            : std_logic;
  SIGNAL Logical_Operator_out625_out1            : std_logic;
  SIGNAL Logical_Operator_out626_out1            : std_logic;
  SIGNAL Logical_Operator_out627_out1            : std_logic;
  SIGNAL Logical_Operator_out628_out1            : std_logic;
  SIGNAL Logical_Operator_out629_out1            : std_logic;
  SIGNAL Logical_Operator_out630_out1            : std_logic;
  SIGNAL Logical_Operator_out631_out1            : std_logic;
  SIGNAL Logical_Operator_out632_out1            : std_logic;
  SIGNAL Logical_Operator_out633_out1            : std_logic;
  SIGNAL Logical_Operator_out634_out1            : std_logic;
  SIGNAL Logical_Operator_out635_out1            : std_logic;
  SIGNAL Logical_Operator_out636_out1            : std_logic;
  SIGNAL Logical_Operator_out637_out1            : std_logic;
  SIGNAL Logical_Operator_out638_out1            : std_logic;
  SIGNAL Logical_Operator_out639_out1            : std_logic;
  SIGNAL Logical_Operator_out640_out1            : std_logic;
  SIGNAL Logical_Operator_out641_out1            : std_logic;
  SIGNAL Logical_Operator_out642_out1            : std_logic;
  SIGNAL Logical_Operator_out643_out1            : std_logic;
  SIGNAL Logical_Operator_out644_out1            : std_logic;
  SIGNAL Logical_Operator_out645_out1            : std_logic;
  SIGNAL Logical_Operator_out646_out1            : std_logic;
  SIGNAL Logical_Operator_out647_out1            : std_logic;
  SIGNAL Logical_Operator_out648_out1            : std_logic;
  SIGNAL Logical_Operator_out649_out1            : std_logic;
  SIGNAL Logical_Operator_out650_out1            : std_logic;
  SIGNAL Logical_Operator_out651_out1            : std_logic;
  SIGNAL Logical_Operator_out652_out1            : std_logic;
  SIGNAL Logical_Operator_out653_out1            : std_logic;
  SIGNAL Logical_Operator_out654_out1            : std_logic;
  SIGNAL Logical_Operator_out655_out1            : std_logic;
  SIGNAL Logical_Operator_out656_out1            : std_logic;
  SIGNAL Logical_Operator_out657_out1            : std_logic;
  SIGNAL Logical_Operator_out658_out1            : std_logic;
  SIGNAL Logical_Operator_out659_out1            : std_logic;
  SIGNAL Logical_Operator_out660_out1            : std_logic;
  SIGNAL Logical_Operator_out661_out1            : std_logic;
  SIGNAL Logical_Operator_out662_out1            : std_logic;
  SIGNAL Logical_Operator_out663_out1            : std_logic;
  SIGNAL Logical_Operator_out664_out1            : std_logic;
  SIGNAL Logical_Operator_out665_out1            : std_logic;
  SIGNAL Logical_Operator_out666_out1            : std_logic;
  SIGNAL Logical_Operator_out667_out1            : std_logic;
  SIGNAL Logical_Operator_out668_out1            : std_logic;
  SIGNAL Logical_Operator_out669_out1            : std_logic;
  SIGNAL Logical_Operator_out670_out1            : std_logic;
  SIGNAL Logical_Operator_out671_out1            : std_logic;
  SIGNAL Logical_Operator_out672_out1            : std_logic;
  SIGNAL Logical_Operator_out673_out1            : std_logic;
  SIGNAL Logical_Operator_out674_out1            : std_logic;
  SIGNAL Logical_Operator_out675_out1            : std_logic;
  SIGNAL Logical_Operator_out676_out1            : std_logic;
  SIGNAL Logical_Operator_out677_out1            : std_logic;
  SIGNAL Logical_Operator_out678_out1            : std_logic;
  SIGNAL Logical_Operator_out679_out1            : std_logic;
  SIGNAL Logical_Operator_out680_out1            : std_logic;
  SIGNAL Logical_Operator_out681_out1            : std_logic;
  SIGNAL Logical_Operator_out682_out1            : std_logic;
  SIGNAL Logical_Operator_out683_out1            : std_logic;
  SIGNAL Logical_Operator_out684_out1            : std_logic;
  SIGNAL Logical_Operator_out685_out1            : std_logic;
  SIGNAL Logical_Operator_out686_out1            : std_logic;
  SIGNAL Logical_Operator_out687_out1            : std_logic;
  SIGNAL Logical_Operator_out688_out1            : std_logic;
  SIGNAL Logical_Operator_out689_out1            : std_logic;
  SIGNAL Logical_Operator_out690_out1            : std_logic;
  SIGNAL Logical_Operator_out691_out1            : std_logic;
  SIGNAL Logical_Operator_out692_out1            : std_logic;
  SIGNAL Logical_Operator_out693_out1            : std_logic;
  SIGNAL Logical_Operator_out694_out1            : std_logic;
  SIGNAL Logical_Operator_out695_out1            : std_logic;
  SIGNAL Logical_Operator_out696_out1            : std_logic;
  SIGNAL Logical_Operator_out697_out1            : std_logic;
  SIGNAL Logical_Operator_out698_out1            : std_logic;
  SIGNAL Logical_Operator_out699_out1            : std_logic;
  SIGNAL Logical_Operator_out700_out1            : std_logic;
  SIGNAL Logical_Operator_out701_out1            : std_logic;
  SIGNAL Logical_Operator_out702_out1            : std_logic;
  SIGNAL Logical_Operator_out703_out1            : std_logic;
  SIGNAL Logical_Operator_out704_out1            : std_logic;
  SIGNAL Logical_Operator_out705_out1            : std_logic;
  SIGNAL Logical_Operator_out706_out1            : std_logic;
  SIGNAL Logical_Operator_out707_out1            : std_logic;
  SIGNAL Logical_Operator_out708_out1            : std_logic;
  SIGNAL Logical_Operator_out709_out1            : std_logic;
  SIGNAL Logical_Operator_out710_out1            : std_logic;
  SIGNAL Logical_Operator_out711_out1            : std_logic;
  SIGNAL Logical_Operator_out712_out1            : std_logic;
  SIGNAL Logical_Operator_out713_out1            : std_logic;
  SIGNAL Logical_Operator_out714_out1            : std_logic;
  SIGNAL Logical_Operator_out715_out1            : std_logic;
  SIGNAL Logical_Operator_out716_out1            : std_logic;
  SIGNAL Logical_Operator_out717_out1            : std_logic;
  SIGNAL Logical_Operator_out718_out1            : std_logic;
  SIGNAL Logical_Operator_out719_out1            : std_logic;
  SIGNAL Logical_Operator_out720_out1            : std_logic;
  SIGNAL Logical_Operator_out721_out1            : std_logic;
  SIGNAL Logical_Operator_out722_out1            : std_logic;
  SIGNAL Logical_Operator_out723_out1            : std_logic;
  SIGNAL Logical_Operator_out724_out1            : std_logic;
  SIGNAL Logical_Operator_out725_out1            : std_logic;
  SIGNAL Logical_Operator_out726_out1            : std_logic;
  SIGNAL Logical_Operator_out727_out1            : std_logic;
  SIGNAL Logical_Operator_out728_out1            : std_logic;
  SIGNAL Logical_Operator_out729_out1            : std_logic;
  SIGNAL Logical_Operator_out730_out1            : std_logic;
  SIGNAL Logical_Operator_out731_out1            : std_logic;
  SIGNAL Logical_Operator_out732_out1            : std_logic;
  SIGNAL Logical_Operator_out733_out1            : std_logic;
  SIGNAL Logical_Operator_out734_out1            : std_logic;
  SIGNAL Logical_Operator_out735_out1            : std_logic;
  SIGNAL Logical_Operator_out736_out1            : std_logic;
  SIGNAL Logical_Operator_out737_out1            : std_logic;
  SIGNAL Logical_Operator_out738_out1            : std_logic;
  SIGNAL Logical_Operator_out739_out1            : std_logic;
  SIGNAL Logical_Operator_out740_out1            : std_logic;
  SIGNAL Logical_Operator_out741_out1            : std_logic;
  SIGNAL Logical_Operator_out742_out1            : std_logic;
  SIGNAL Logical_Operator_out743_out1            : std_logic;
  SIGNAL Logical_Operator_out744_out1            : std_logic;
  SIGNAL Logical_Operator_out745_out1            : std_logic;
  SIGNAL Logical_Operator_out746_out1            : std_logic;
  SIGNAL Logical_Operator_out747_out1            : std_logic;
  SIGNAL Logical_Operator_out748_out1            : std_logic;
  SIGNAL Logical_Operator_out749_out1            : std_logic;
  SIGNAL Logical_Operator_out750_out1            : std_logic;
  SIGNAL Logical_Operator_out751_out1            : std_logic;
  SIGNAL Logical_Operator_out752_out1            : std_logic;
  SIGNAL Logical_Operator_out753_out1            : std_logic;
  SIGNAL Logical_Operator_out754_out1            : std_logic;
  SIGNAL Logical_Operator_out755_out1            : std_logic;
  SIGNAL Logical_Operator_out756_out1            : std_logic;
  SIGNAL Logical_Operator_out757_out1            : std_logic;
  SIGNAL Logical_Operator_out758_out1            : std_logic;
  SIGNAL Logical_Operator_out759_out1            : std_logic;
  SIGNAL Logical_Operator_out760_out1            : std_logic;
  SIGNAL Logical_Operator_out761_out1            : std_logic;
  SIGNAL Logical_Operator_out762_out1            : std_logic;
  SIGNAL Logical_Operator_out763_out1            : std_logic;
  SIGNAL Logical_Operator_out764_out1            : std_logic;
  SIGNAL Logical_Operator_out765_out1            : std_logic;
  SIGNAL Logical_Operator_out766_out1            : std_logic;
  SIGNAL Logical_Operator_out767_out1            : std_logic;
  SIGNAL Logical_Operator_out768_out1            : std_logic;
  SIGNAL Logical_Operator_out769_out1            : std_logic;
  SIGNAL Logical_Operator_out770_out1            : std_logic;
  SIGNAL Logical_Operator_out771_out1            : std_logic;
  SIGNAL Logical_Operator_out772_out1            : std_logic;
  SIGNAL Logical_Operator_out773_out1            : std_logic;
  SIGNAL Logical_Operator_out774_out1            : std_logic;
  SIGNAL Logical_Operator_out775_out1            : std_logic;
  SIGNAL Logical_Operator_out776_out1            : std_logic;
  SIGNAL Logical_Operator_out777_out1            : std_logic;
  SIGNAL Logical_Operator_out778_out1            : std_logic;
  SIGNAL Logical_Operator_out779_out1            : std_logic;
  SIGNAL Logical_Operator_out780_out1            : std_logic;
  SIGNAL Logical_Operator_out781_out1            : std_logic;
  SIGNAL Logical_Operator_out782_out1            : std_logic;
  SIGNAL Logical_Operator_out783_out1            : std_logic;
  SIGNAL Logical_Operator_out784_out1            : std_logic;
  SIGNAL Logical_Operator_out785_out1            : std_logic;
  SIGNAL Logical_Operator_out786_out1            : std_logic;
  SIGNAL Logical_Operator_out787_out1            : std_logic;
  SIGNAL Logical_Operator_out788_out1            : std_logic;
  SIGNAL Logical_Operator_out789_out1            : std_logic;
  SIGNAL Logical_Operator_out790_out1            : std_logic;
  SIGNAL Logical_Operator_out791_out1            : std_logic;
  SIGNAL Logical_Operator_out792_out1            : std_logic;
  SIGNAL Logical_Operator_out793_out1            : std_logic;
  SIGNAL Logical_Operator_out794_out1            : std_logic;
  SIGNAL Logical_Operator_out795_out1            : std_logic;
  SIGNAL Logical_Operator_out796_out1            : std_logic;
  SIGNAL Logical_Operator_out797_out1            : std_logic;
  SIGNAL Logical_Operator_out798_out1            : std_logic;
  SIGNAL Logical_Operator_out799_out1            : std_logic;
  SIGNAL Logical_Operator_out800_out1            : std_logic;
  SIGNAL Logical_Operator_out801_out1            : std_logic;
  SIGNAL Logical_Operator_out802_out1            : std_logic;
  SIGNAL Logical_Operator_out803_out1            : std_logic;
  SIGNAL Logical_Operator_out804_out1            : std_logic;
  SIGNAL Logical_Operator_out805_out1            : std_logic;
  SIGNAL Logical_Operator_out806_out1            : std_logic;
  SIGNAL Logical_Operator_out807_out1            : std_logic;
  SIGNAL Logical_Operator_out808_out1            : std_logic;
  SIGNAL Logical_Operator_out809_out1            : std_logic;
  SIGNAL Logical_Operator_out810_out1            : std_logic;
  SIGNAL Logical_Operator_out811_out1            : std_logic;
  SIGNAL Logical_Operator_out812_out1            : std_logic;
  SIGNAL Logical_Operator_out813_out1            : std_logic;
  SIGNAL Logical_Operator_out814_out1            : std_logic;
  SIGNAL Logical_Operator_out815_out1            : std_logic;
  SIGNAL Logical_Operator_out816_out1            : std_logic;
  SIGNAL Logical_Operator_out817_out1            : std_logic;
  SIGNAL Logical_Operator_out818_out1            : std_logic;
  SIGNAL Logical_Operator_out819_out1            : std_logic;
  SIGNAL Logical_Operator_out820_out1            : std_logic;
  SIGNAL Logical_Operator_out821_out1            : std_logic;
  SIGNAL Logical_Operator_out822_out1            : std_logic;
  SIGNAL Logical_Operator_out823_out1            : std_logic;
  SIGNAL Logical_Operator_out824_out1            : std_logic;
  SIGNAL Logical_Operator_out825_out1            : std_logic;
  SIGNAL Logical_Operator_out826_out1            : std_logic;
  SIGNAL Logical_Operator_out827_out1            : std_logic;
  SIGNAL Logical_Operator_out828_out1            : std_logic;
  SIGNAL Logical_Operator_out829_out1            : std_logic;
  SIGNAL Logical_Operator_out830_out1            : std_logic;
  SIGNAL Logical_Operator_out831_out1            : std_logic;
  SIGNAL Logical_Operator_out832_out1            : std_logic;
  SIGNAL Logical_Operator_out833_out1            : std_logic;
  SIGNAL Logical_Operator_out834_out1            : std_logic;
  SIGNAL Logical_Operator_out835_out1            : std_logic;
  SIGNAL Logical_Operator_out836_out1            : std_logic;
  SIGNAL Logical_Operator_out837_out1            : std_logic;
  SIGNAL Logical_Operator_out838_out1            : std_logic;
  SIGNAL Logical_Operator_out839_out1            : std_logic;
  SIGNAL Logical_Operator_out840_out1            : std_logic;
  SIGNAL Logical_Operator_out841_out1            : std_logic;
  SIGNAL Logical_Operator_out842_out1            : std_logic;
  SIGNAL Logical_Operator_out843_out1            : std_logic;
  SIGNAL Logical_Operator_out844_out1            : std_logic;
  SIGNAL Logical_Operator_out845_out1            : std_logic;
  SIGNAL Logical_Operator_out846_out1            : std_logic;
  SIGNAL Logical_Operator_out847_out1            : std_logic;
  SIGNAL Logical_Operator_out848_out1            : std_logic;
  SIGNAL Logical_Operator_out849_out1            : std_logic;
  SIGNAL Logical_Operator_out850_out1            : std_logic;
  SIGNAL Logical_Operator_out851_out1            : std_logic;
  SIGNAL Logical_Operator_out852_out1            : std_logic;
  SIGNAL Logical_Operator_out853_out1            : std_logic;
  SIGNAL Logical_Operator_out854_out1            : std_logic;
  SIGNAL Logical_Operator_out855_out1            : std_logic;
  SIGNAL Logical_Operator_out856_out1            : std_logic;
  SIGNAL Logical_Operator_out857_out1            : std_logic;
  SIGNAL Logical_Operator_out858_out1            : std_logic;
  SIGNAL Logical_Operator_out859_out1            : std_logic;
  SIGNAL Logical_Operator_out860_out1            : std_logic;
  SIGNAL Logical_Operator_out861_out1            : std_logic;
  SIGNAL Logical_Operator_out862_out1            : std_logic;
  SIGNAL Logical_Operator_out863_out1            : std_logic;
  SIGNAL Logical_Operator_out864_out1            : std_logic;
  SIGNAL Logical_Operator_out865_out1            : std_logic;
  SIGNAL Logical_Operator_out866_out1            : std_logic;
  SIGNAL Logical_Operator_out867_out1            : std_logic;
  SIGNAL Logical_Operator_out868_out1            : std_logic;
  SIGNAL Logical_Operator_out869_out1            : std_logic;
  SIGNAL Logical_Operator_out870_out1            : std_logic;
  SIGNAL Logical_Operator_out871_out1            : std_logic;
  SIGNAL Logical_Operator_out872_out1            : std_logic;
  SIGNAL Logical_Operator_out873_out1            : std_logic;
  SIGNAL Logical_Operator_out874_out1            : std_logic;
  SIGNAL Logical_Operator_out875_out1            : std_logic;
  SIGNAL Logical_Operator_out876_out1            : std_logic;
  SIGNAL Logical_Operator_out877_out1            : std_logic;
  SIGNAL Logical_Operator_out878_out1            : std_logic;
  SIGNAL Logical_Operator_out879_out1            : std_logic;
  SIGNAL Logical_Operator_out880_out1            : std_logic;
  SIGNAL Logical_Operator_out881_out1            : std_logic;
  SIGNAL Logical_Operator_out882_out1            : std_logic;
  SIGNAL Logical_Operator_out883_out1            : std_logic;
  SIGNAL Logical_Operator_out884_out1            : std_logic;
  SIGNAL Logical_Operator_out885_out1            : std_logic;
  SIGNAL Logical_Operator_out886_out1            : std_logic;
  SIGNAL Logical_Operator_out887_out1            : std_logic;
  SIGNAL Logical_Operator_out888_out1            : std_logic;
  SIGNAL Logical_Operator_out889_out1            : std_logic;
  SIGNAL Logical_Operator_out890_out1            : std_logic;
  SIGNAL Logical_Operator_out891_out1            : std_logic;
  SIGNAL Logical_Operator_out892_out1            : std_logic;
  SIGNAL Logical_Operator_out893_out1            : std_logic;
  SIGNAL Logical_Operator_out894_out1            : std_logic;
  SIGNAL Logical_Operator_out895_out1            : std_logic;
  SIGNAL Logical_Operator_out896_out1            : std_logic;
  SIGNAL Logical_Operator_out897_out1            : std_logic;
  SIGNAL Logical_Operator_out898_out1            : std_logic;
  SIGNAL Logical_Operator_out899_out1            : std_logic;
  SIGNAL Logical_Operator_out900_out1            : std_logic;
  SIGNAL Logical_Operator_out901_out1            : std_logic;
  SIGNAL Logical_Operator_out902_out1            : std_logic;
  SIGNAL Logical_Operator_out903_out1            : std_logic;
  SIGNAL Logical_Operator_out904_out1            : std_logic;
  SIGNAL Logical_Operator_out905_out1            : std_logic;
  SIGNAL Logical_Operator_out906_out1            : std_logic;
  SIGNAL Logical_Operator_out907_out1            : std_logic;
  SIGNAL Logical_Operator_out908_out1            : std_logic;
  SIGNAL Logical_Operator_out909_out1            : std_logic;
  SIGNAL Logical_Operator_out910_out1            : std_logic;
  SIGNAL Logical_Operator_out911_out1            : std_logic;
  SIGNAL Logical_Operator_out912_out1            : std_logic;
  SIGNAL Logical_Operator_out913_out1            : std_logic;
  SIGNAL Logical_Operator_out914_out1            : std_logic;
  SIGNAL Logical_Operator_out915_out1            : std_logic;
  SIGNAL Logical_Operator_out916_out1            : std_logic;
  SIGNAL Logical_Operator_out917_out1            : std_logic;
  SIGNAL Logical_Operator_out918_out1            : std_logic;
  SIGNAL Logical_Operator_out919_out1            : std_logic;
  SIGNAL Logical_Operator_out920_out1            : std_logic;
  SIGNAL Logical_Operator_out921_out1            : std_logic;
  SIGNAL Logical_Operator_out922_out1            : std_logic;
  SIGNAL Logical_Operator_out923_out1            : std_logic;
  SIGNAL Logical_Operator_out924_out1            : std_logic;
  SIGNAL Logical_Operator_out925_out1            : std_logic;
  SIGNAL Logical_Operator_out926_out1            : std_logic;
  SIGNAL Logical_Operator_out927_out1            : std_logic;
  SIGNAL Logical_Operator_out928_out1            : std_logic;
  SIGNAL Logical_Operator_out929_out1            : std_logic;
  SIGNAL Logical_Operator_out930_out1            : std_logic;
  SIGNAL Logical_Operator_out931_out1            : std_logic;
  SIGNAL Logical_Operator_out932_out1            : std_logic;
  SIGNAL Logical_Operator_out933_out1            : std_logic;
  SIGNAL Logical_Operator_out934_out1            : std_logic;
  SIGNAL Logical_Operator_out935_out1            : std_logic;
  SIGNAL Logical_Operator_out936_out1            : std_logic;
  SIGNAL Logical_Operator_out937_out1            : std_logic;
  SIGNAL Logical_Operator_out938_out1            : std_logic;
  SIGNAL Logical_Operator_out939_out1            : std_logic;
  SIGNAL Logical_Operator_out940_out1            : std_logic;
  SIGNAL Logical_Operator_out941_out1            : std_logic;
  SIGNAL Logical_Operator_out942_out1            : std_logic;
  SIGNAL Logical_Operator_out943_out1            : std_logic;
  SIGNAL Logical_Operator_out944_out1            : std_logic;
  SIGNAL Logical_Operator_out945_out1            : std_logic;
  SIGNAL Logical_Operator_out946_out1            : std_logic;
  SIGNAL Logical_Operator_out947_out1            : std_logic;
  SIGNAL Logical_Operator_out948_out1            : std_logic;
  SIGNAL Logical_Operator_out949_out1            : std_logic;
  SIGNAL Logical_Operator_out950_out1            : std_logic;
  SIGNAL Logical_Operator_out951_out1            : std_logic;
  SIGNAL Logical_Operator_out952_out1            : std_logic;
  SIGNAL Logical_Operator_out953_out1            : std_logic;
  SIGNAL Logical_Operator_out954_out1            : std_logic;
  SIGNAL Logical_Operator_out955_out1            : std_logic;
  SIGNAL Logical_Operator_out956_out1            : std_logic;
  SIGNAL Logical_Operator_out957_out1            : std_logic;
  SIGNAL Logical_Operator_out958_out1            : std_logic;
  SIGNAL Logical_Operator_out959_out1            : std_logic;
  SIGNAL Logical_Operator_out960_out1            : std_logic;
  SIGNAL Logical_Operator_out961_out1            : std_logic;
  SIGNAL Logical_Operator_out962_out1            : std_logic;
  SIGNAL Logical_Operator_out963_out1            : std_logic;
  SIGNAL Logical_Operator_out964_out1            : std_logic;
  SIGNAL Logical_Operator_out965_out1            : std_logic;
  SIGNAL Logical_Operator_out966_out1            : std_logic;
  SIGNAL Logical_Operator_out967_out1            : std_logic;
  SIGNAL Logical_Operator_out968_out1            : std_logic;
  SIGNAL Logical_Operator_out969_out1            : std_logic;
  SIGNAL Logical_Operator_out970_out1            : std_logic;
  SIGNAL Logical_Operator_out971_out1            : std_logic;
  SIGNAL Logical_Operator_out972_out1            : std_logic;
  SIGNAL Logical_Operator_out973_out1            : std_logic;
  SIGNAL Logical_Operator_out974_out1            : std_logic;
  SIGNAL Logical_Operator_out975_out1            : std_logic;
  SIGNAL Logical_Operator_out976_out1            : std_logic;
  SIGNAL Logical_Operator_out977_out1            : std_logic;
  SIGNAL Logical_Operator_out978_out1            : std_logic;
  SIGNAL Logical_Operator_out979_out1            : std_logic;
  SIGNAL Logical_Operator_out980_out1            : std_logic;
  SIGNAL Logical_Operator_out981_out1            : std_logic;
  SIGNAL Logical_Operator_out982_out1            : std_logic;
  SIGNAL Logical_Operator_out983_out1            : std_logic;
  SIGNAL Logical_Operator_out984_out1            : std_logic;
  SIGNAL Logical_Operator_out985_out1            : std_logic;
  SIGNAL Logical_Operator_out986_out1            : std_logic;
  SIGNAL Logical_Operator_out987_out1            : std_logic;
  SIGNAL Logical_Operator_out988_out1            : std_logic;
  SIGNAL Logical_Operator_out989_out1            : std_logic;
  SIGNAL Logical_Operator_out990_out1            : std_logic;
  SIGNAL Logical_Operator_out991_out1            : std_logic;
  SIGNAL Logical_Operator_out992_out1            : std_logic;
  SIGNAL Logical_Operator_out993_out1            : std_logic;
  SIGNAL Logical_Operator_out994_out1            : std_logic;
  SIGNAL Logical_Operator_out995_out1            : std_logic;
  SIGNAL Logical_Operator_out996_out1            : std_logic;
  SIGNAL Logical_Operator_out997_out1            : std_logic;
  SIGNAL Logical_Operator_out998_out1            : std_logic;
  SIGNAL Logical_Operator_out999_out1            : std_logic;
  SIGNAL Logical_Operator_out1000_out1            : std_logic;
  SIGNAL Logical_Operator_out1001_out1            : std_logic;
  SIGNAL Logical_Operator_out1002_out1            : std_logic;
  SIGNAL Logical_Operator_out1003_out1            : std_logic;
  SIGNAL Logical_Operator_out1004_out1            : std_logic;
  SIGNAL Logical_Operator_out1005_out1            : std_logic;
  SIGNAL Logical_Operator_out1006_out1            : std_logic;
  SIGNAL Logical_Operator_out1007_out1            : std_logic;
  SIGNAL Logical_Operator_out1008_out1            : std_logic;
  SIGNAL Logical_Operator_out1009_out1            : std_logic;
  SIGNAL Logical_Operator_out1010_out1            : std_logic;
  SIGNAL Logical_Operator_out1011_out1            : std_logic;
  SIGNAL Logical_Operator_out1012_out1            : std_logic;
  SIGNAL Logical_Operator_out1013_out1            : std_logic;
  SIGNAL Logical_Operator_out1014_out1            : std_logic;
  SIGNAL Logical_Operator_out1015_out1            : std_logic;
  SIGNAL Logical_Operator_out1016_out1            : std_logic;
  SIGNAL Logical_Operator_out1017_out1            : std_logic;
  SIGNAL Logical_Operator_out1018_out1            : std_logic;
  SIGNAL Logical_Operator_out1019_out1            : std_logic;
  SIGNAL Logical_Operator_out1020_out1            : std_logic;
  SIGNAL Logical_Operator_out1021_out1            : std_logic;
  SIGNAL Logical_Operator_out1022_out1            : std_logic;
  SIGNAL Logical_Operator_out1023_out1            : std_logic;
  SIGNAL Logical_Operator_out1024_out1            : std_logic;

BEGIN

  Logical_Operator_out1_out1 <= in1 XOR in2;

  Logical_Operator_out2_out1 <= in3 XOR in4;

  Logical_Operator_out3_out1 <= in5 XOR in6;

  Logical_Operator_out4_out1 <= in7 XOR in8;

  Logical_Operator_out5_out1 <= in9 XOR in10;

  Logical_Operator_out6_out1 <= in11 XOR in12;

  Logical_Operator_out7_out1 <= in13 XOR in14;

  Logical_Operator_out8_out1 <= in15 XOR in16;

  Logical_Operator_out9_out1 <= in17 XOR in18;

  Logical_Operator_out10_out1 <= in19 XOR in20;

  Logical_Operator_out11_out1 <= in21 XOR in22;

  Logical_Operator_out12_out1 <= in23 XOR in24;

  Logical_Operator_out13_out1 <= in25 XOR in26;

  Logical_Operator_out14_out1 <= in27 XOR in28;

  Logical_Operator_out15_out1 <= in29 XOR in30;

  Logical_Operator_out16_out1 <= in31 XOR in32;

  Logical_Operator_out17_out1 <= in33 XOR in34;

  Logical_Operator_out18_out1 <= in35 XOR in36;

  Logical_Operator_out19_out1 <= in37 XOR in38;

  Logical_Operator_out20_out1 <= in39 XOR in40;

  Logical_Operator_out21_out1 <= in41 XOR in42;

  Logical_Operator_out22_out1 <= in43 XOR in44;

  Logical_Operator_out23_out1 <= in45 XOR in46;

  Logical_Operator_out24_out1 <= in47 XOR in48;

  Logical_Operator_out25_out1 <= in49 XOR in50;

  Logical_Operator_out26_out1 <= in51 XOR in52;

  Logical_Operator_out27_out1 <= in53 XOR in54;

  Logical_Operator_out28_out1 <= in55 XOR in56;

  Logical_Operator_out29_out1 <= in57 XOR in58;

  Logical_Operator_out30_out1 <= in59 XOR in60;

  Logical_Operator_out31_out1 <= in61 XOR in62;

  Logical_Operator_out32_out1 <= in63 XOR in64;

  Logical_Operator_out33_out1 <= in65 XOR in66;

  Logical_Operator_out34_out1 <= in67 XOR in68;

  Logical_Operator_out35_out1 <= in69 XOR in70;

  Logical_Operator_out36_out1 <= in71 XOR in72;

  Logical_Operator_out37_out1 <= in73 XOR in74;

  Logical_Operator_out38_out1 <= in75 XOR in76;

  Logical_Operator_out39_out1 <= in77 XOR in78;

  Logical_Operator_out40_out1 <= in79 XOR in80;

  Logical_Operator_out41_out1 <= in81 XOR in82;

  Logical_Operator_out42_out1 <= in83 XOR in84;

  Logical_Operator_out43_out1 <= in85 XOR in86;

  Logical_Operator_out44_out1 <= in87 XOR in88;

  Logical_Operator_out45_out1 <= in89 XOR in90;

  Logical_Operator_out46_out1 <= in91 XOR in92;

  Logical_Operator_out47_out1 <= in93 XOR in94;

  Logical_Operator_out48_out1 <= in95 XOR in96;

  Logical_Operator_out49_out1 <= in97 XOR in98;

  Logical_Operator_out50_out1 <= in99 XOR in100;

  Logical_Operator_out51_out1 <= in101 XOR in102;

  Logical_Operator_out52_out1 <= in103 XOR in104;

  Logical_Operator_out53_out1 <= in105 XOR in106;

  Logical_Operator_out54_out1 <= in107 XOR in108;

  Logical_Operator_out55_out1 <= in109 XOR in110;

  Logical_Operator_out56_out1 <= in111 XOR in112;

  Logical_Operator_out57_out1 <= in113 XOR in114;

  Logical_Operator_out58_out1 <= in115 XOR in116;

  Logical_Operator_out59_out1 <= in117 XOR in118;

  Logical_Operator_out60_out1 <= in119 XOR in120;

  Logical_Operator_out61_out1 <= in121 XOR in122;

  Logical_Operator_out62_out1 <= in123 XOR in124;

  Logical_Operator_out63_out1 <= in125 XOR in126;

  Logical_Operator_out64_out1 <= in127 XOR in128;

  Logical_Operator_out65_out1 <= in129 XOR in130;

  Logical_Operator_out66_out1 <= in131 XOR in132;

  Logical_Operator_out67_out1 <= in133 XOR in134;

  Logical_Operator_out68_out1 <= in135 XOR in136;

  Logical_Operator_out69_out1 <= in137 XOR in138;

  Logical_Operator_out70_out1 <= in139 XOR in140;

  Logical_Operator_out71_out1 <= in141 XOR in142;

  Logical_Operator_out72_out1 <= in143 XOR in144;

  Logical_Operator_out73_out1 <= in145 XOR in146;

  Logical_Operator_out74_out1 <= in147 XOR in148;

  Logical_Operator_out75_out1 <= in149 XOR in150;

  Logical_Operator_out76_out1 <= in151 XOR in152;

  Logical_Operator_out77_out1 <= in153 XOR in154;

  Logical_Operator_out78_out1 <= in155 XOR in156;

  Logical_Operator_out79_out1 <= in157 XOR in158;

  Logical_Operator_out80_out1 <= in159 XOR in160;

  Logical_Operator_out81_out1 <= in161 XOR in162;

  Logical_Operator_out82_out1 <= in163 XOR in164;

  Logical_Operator_out83_out1 <= in165 XOR in166;

  Logical_Operator_out84_out1 <= in167 XOR in168;

  Logical_Operator_out85_out1 <= in169 XOR in170;

  Logical_Operator_out86_out1 <= in171 XOR in172;

  Logical_Operator_out87_out1 <= in173 XOR in174;

  Logical_Operator_out88_out1 <= in175 XOR in176;

  Logical_Operator_out89_out1 <= in177 XOR in178;

  Logical_Operator_out90_out1 <= in179 XOR in180;

  Logical_Operator_out91_out1 <= in181 XOR in182;

  Logical_Operator_out92_out1 <= in183 XOR in184;

  Logical_Operator_out93_out1 <= in185 XOR in186;

  Logical_Operator_out94_out1 <= in187 XOR in188;

  Logical_Operator_out95_out1 <= in189 XOR in190;

  Logical_Operator_out96_out1 <= in191 XOR in192;

  Logical_Operator_out97_out1 <= in193 XOR in194;

  Logical_Operator_out98_out1 <= in195 XOR in196;

  Logical_Operator_out99_out1 <= in197 XOR in198;

  Logical_Operator_out100_out1 <= in199 XOR in200;

  Logical_Operator_out101_out1 <= in201 XOR in202;

  Logical_Operator_out102_out1 <= in203 XOR in204;

  Logical_Operator_out103_out1 <= in205 XOR in206;

  Logical_Operator_out104_out1 <= in207 XOR in208;

  Logical_Operator_out105_out1 <= in209 XOR in210;

  Logical_Operator_out106_out1 <= in211 XOR in212;

  Logical_Operator_out107_out1 <= in213 XOR in214;

  Logical_Operator_out108_out1 <= in215 XOR in216;

  Logical_Operator_out109_out1 <= in217 XOR in218;

  Logical_Operator_out110_out1 <= in219 XOR in220;

  Logical_Operator_out111_out1 <= in221 XOR in222;

  Logical_Operator_out112_out1 <= in223 XOR in224;

  Logical_Operator_out113_out1 <= in225 XOR in226;

  Logical_Operator_out114_out1 <= in227 XOR in228;

  Logical_Operator_out115_out1 <= in229 XOR in230;

  Logical_Operator_out116_out1 <= in231 XOR in232;

  Logical_Operator_out117_out1 <= in233 XOR in234;

  Logical_Operator_out118_out1 <= in235 XOR in236;

  Logical_Operator_out119_out1 <= in237 XOR in238;

  Logical_Operator_out120_out1 <= in239 XOR in240;

  Logical_Operator_out121_out1 <= in241 XOR in242;

  Logical_Operator_out122_out1 <= in243 XOR in244;

  Logical_Operator_out123_out1 <= in245 XOR in246;

  Logical_Operator_out124_out1 <= in247 XOR in248;

  Logical_Operator_out125_out1 <= in249 XOR in250;

  Logical_Operator_out126_out1 <= in251 XOR in252;

  Logical_Operator_out127_out1 <= in253 XOR in254;

  Logical_Operator_out128_out1 <= in255 XOR in256;

  Logical_Operator_out129_out1 <= Logical_Operator_out1_out1 XOR Logical_Operator_out2_out1;

  Logical_Operator_out130_out1 <= in2 XOR in4;

  Logical_Operator_out131_out1 <= Logical_Operator_out3_out1 XOR Logical_Operator_out4_out1;

  Logical_Operator_out132_out1 <= in6 XOR in8;

  Logical_Operator_out133_out1 <= Logical_Operator_out5_out1 XOR Logical_Operator_out6_out1;

  Logical_Operator_out134_out1 <= in10 XOR in12;

  Logical_Operator_out135_out1 <= Logical_Operator_out7_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out136_out1 <= in14 XOR in16;

  Logical_Operator_out137_out1 <= Logical_Operator_out9_out1 XOR Logical_Operator_out10_out1;

  Logical_Operator_out138_out1 <= in18 XOR in20;

  Logical_Operator_out139_out1 <= Logical_Operator_out11_out1 XOR Logical_Operator_out12_out1;

  Logical_Operator_out140_out1 <= in22 XOR in24;

  Logical_Operator_out141_out1 <= Logical_Operator_out13_out1 XOR Logical_Operator_out14_out1;

  Logical_Operator_out142_out1 <= in26 XOR in28;

  Logical_Operator_out143_out1 <= Logical_Operator_out15_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out144_out1 <= in30 XOR in32;

  Logical_Operator_out145_out1 <= Logical_Operator_out17_out1 XOR Logical_Operator_out18_out1;

  Logical_Operator_out146_out1 <= in34 XOR in36;

  Logical_Operator_out147_out1 <= Logical_Operator_out19_out1 XOR Logical_Operator_out20_out1;

  Logical_Operator_out148_out1 <= in38 XOR in40;

  Logical_Operator_out149_out1 <= Logical_Operator_out21_out1 XOR Logical_Operator_out22_out1;

  Logical_Operator_out150_out1 <= in42 XOR in44;

  Logical_Operator_out151_out1 <= Logical_Operator_out23_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out152_out1 <= in46 XOR in48;

  Logical_Operator_out153_out1 <= Logical_Operator_out25_out1 XOR Logical_Operator_out26_out1;

  Logical_Operator_out154_out1 <= in50 XOR in52;

  Logical_Operator_out155_out1 <= Logical_Operator_out27_out1 XOR Logical_Operator_out28_out1;

  Logical_Operator_out156_out1 <= in54 XOR in56;

  Logical_Operator_out157_out1 <= Logical_Operator_out29_out1 XOR Logical_Operator_out30_out1;

  Logical_Operator_out158_out1 <= in58 XOR in60;

  Logical_Operator_out159_out1 <= Logical_Operator_out31_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out160_out1 <= in62 XOR in64;

  Logical_Operator_out161_out1 <= Logical_Operator_out33_out1 XOR Logical_Operator_out34_out1;

  Logical_Operator_out162_out1 <= in66 XOR in68;

  Logical_Operator_out163_out1 <= Logical_Operator_out35_out1 XOR Logical_Operator_out36_out1;

  Logical_Operator_out164_out1 <= in70 XOR in72;

  Logical_Operator_out165_out1 <= Logical_Operator_out37_out1 XOR Logical_Operator_out38_out1;

  Logical_Operator_out166_out1 <= in74 XOR in76;

  Logical_Operator_out167_out1 <= Logical_Operator_out39_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out168_out1 <= in78 XOR in80;

  Logical_Operator_out169_out1 <= Logical_Operator_out41_out1 XOR Logical_Operator_out42_out1;

  Logical_Operator_out170_out1 <= in82 XOR in84;

  Logical_Operator_out171_out1 <= Logical_Operator_out43_out1 XOR Logical_Operator_out44_out1;

  Logical_Operator_out172_out1 <= in86 XOR in88;

  Logical_Operator_out173_out1 <= Logical_Operator_out45_out1 XOR Logical_Operator_out46_out1;

  Logical_Operator_out174_out1 <= in90 XOR in92;

  Logical_Operator_out175_out1 <= Logical_Operator_out47_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out176_out1 <= in94 XOR in96;

  Logical_Operator_out177_out1 <= Logical_Operator_out49_out1 XOR Logical_Operator_out50_out1;

  Logical_Operator_out178_out1 <= in98 XOR in100;

  Logical_Operator_out179_out1 <= Logical_Operator_out51_out1 XOR Logical_Operator_out52_out1;

  Logical_Operator_out180_out1 <= in102 XOR in104;

  Logical_Operator_out181_out1 <= Logical_Operator_out53_out1 XOR Logical_Operator_out54_out1;

  Logical_Operator_out182_out1 <= in106 XOR in108;

  Logical_Operator_out183_out1 <= Logical_Operator_out55_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out184_out1 <= in110 XOR in112;

  Logical_Operator_out185_out1 <= Logical_Operator_out57_out1 XOR Logical_Operator_out58_out1;

  Logical_Operator_out186_out1 <= in114 XOR in116;

  Logical_Operator_out187_out1 <= Logical_Operator_out59_out1 XOR Logical_Operator_out60_out1;

  Logical_Operator_out188_out1 <= in118 XOR in120;

  Logical_Operator_out189_out1 <= Logical_Operator_out61_out1 XOR Logical_Operator_out62_out1;

  Logical_Operator_out190_out1 <= in122 XOR in124;

  Logical_Operator_out191_out1 <= Logical_Operator_out63_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out192_out1 <= in126 XOR in128;

  Logical_Operator_out193_out1 <= Logical_Operator_out65_out1 XOR Logical_Operator_out66_out1;

  Logical_Operator_out194_out1 <= in130 XOR in132;

  Logical_Operator_out195_out1 <= Logical_Operator_out67_out1 XOR Logical_Operator_out68_out1;

  Logical_Operator_out196_out1 <= in134 XOR in136;

  Logical_Operator_out197_out1 <= Logical_Operator_out69_out1 XOR Logical_Operator_out70_out1;

  Logical_Operator_out198_out1 <= in138 XOR in140;

  Logical_Operator_out199_out1 <= Logical_Operator_out71_out1 XOR Logical_Operator_out72_out1;

  Logical_Operator_out200_out1 <= in142 XOR in144;

  Logical_Operator_out201_out1 <= Logical_Operator_out73_out1 XOR Logical_Operator_out74_out1;

  Logical_Operator_out202_out1 <= in146 XOR in148;

  Logical_Operator_out203_out1 <= Logical_Operator_out75_out1 XOR Logical_Operator_out76_out1;

  Logical_Operator_out204_out1 <= in150 XOR in152;

  Logical_Operator_out205_out1 <= Logical_Operator_out77_out1 XOR Logical_Operator_out78_out1;

  Logical_Operator_out206_out1 <= in154 XOR in156;

  Logical_Operator_out207_out1 <= Logical_Operator_out79_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out208_out1 <= in158 XOR in160;

  Logical_Operator_out209_out1 <= Logical_Operator_out81_out1 XOR Logical_Operator_out82_out1;

  Logical_Operator_out210_out1 <= in162 XOR in164;

  Logical_Operator_out211_out1 <= Logical_Operator_out83_out1 XOR Logical_Operator_out84_out1;

  Logical_Operator_out212_out1 <= in166 XOR in168;

  Logical_Operator_out213_out1 <= Logical_Operator_out85_out1 XOR Logical_Operator_out86_out1;

  Logical_Operator_out214_out1 <= in170 XOR in172;

  Logical_Operator_out215_out1 <= Logical_Operator_out87_out1 XOR Logical_Operator_out88_out1;

  Logical_Operator_out216_out1 <= in174 XOR in176;

  Logical_Operator_out217_out1 <= Logical_Operator_out89_out1 XOR Logical_Operator_out90_out1;

  Logical_Operator_out218_out1 <= in178 XOR in180;

  Logical_Operator_out219_out1 <= Logical_Operator_out91_out1 XOR Logical_Operator_out92_out1;

  Logical_Operator_out220_out1 <= in182 XOR in184;

  Logical_Operator_out221_out1 <= Logical_Operator_out93_out1 XOR Logical_Operator_out94_out1;

  Logical_Operator_out222_out1 <= in186 XOR in188;

  Logical_Operator_out223_out1 <= Logical_Operator_out95_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out224_out1 <= in190 XOR in192;

  Logical_Operator_out225_out1 <= Logical_Operator_out97_out1 XOR Logical_Operator_out98_out1;

  Logical_Operator_out226_out1 <= in194 XOR in196;

  Logical_Operator_out227_out1 <= Logical_Operator_out99_out1 XOR Logical_Operator_out100_out1;

  Logical_Operator_out228_out1 <= in198 XOR in200;

  Logical_Operator_out229_out1 <= Logical_Operator_out101_out1 XOR Logical_Operator_out102_out1;

  Logical_Operator_out230_out1 <= in202 XOR in204;

  Logical_Operator_out231_out1 <= Logical_Operator_out103_out1 XOR Logical_Operator_out104_out1;

  Logical_Operator_out232_out1 <= in206 XOR in208;

  Logical_Operator_out233_out1 <= Logical_Operator_out105_out1 XOR Logical_Operator_out106_out1;

  Logical_Operator_out234_out1 <= in210 XOR in212;

  Logical_Operator_out235_out1 <= Logical_Operator_out107_out1 XOR Logical_Operator_out108_out1;

  Logical_Operator_out236_out1 <= in214 XOR in216;

  Logical_Operator_out237_out1 <= Logical_Operator_out109_out1 XOR Logical_Operator_out110_out1;

  Logical_Operator_out238_out1 <= in218 XOR in220;

  Logical_Operator_out239_out1 <= Logical_Operator_out111_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out240_out1 <= in222 XOR in224;

  Logical_Operator_out241_out1 <= Logical_Operator_out113_out1 XOR Logical_Operator_out114_out1;

  Logical_Operator_out242_out1 <= in226 XOR in228;

  Logical_Operator_out243_out1 <= Logical_Operator_out115_out1 XOR Logical_Operator_out116_out1;

  Logical_Operator_out244_out1 <= in230 XOR in232;

  Logical_Operator_out245_out1 <= Logical_Operator_out117_out1 XOR Logical_Operator_out118_out1;

  Logical_Operator_out246_out1 <= in234 XOR in236;

  Logical_Operator_out247_out1 <= Logical_Operator_out119_out1 XOR Logical_Operator_out120_out1;

  Logical_Operator_out248_out1 <= in238 XOR in240;

  Logical_Operator_out249_out1 <= Logical_Operator_out121_out1 XOR Logical_Operator_out122_out1;

  Logical_Operator_out250_out1 <= in242 XOR in244;

  Logical_Operator_out251_out1 <= Logical_Operator_out123_out1 XOR Logical_Operator_out124_out1;

  Logical_Operator_out252_out1 <= in246 XOR in248;

  Logical_Operator_out253_out1 <= Logical_Operator_out125_out1 XOR Logical_Operator_out126_out1;

  Logical_Operator_out254_out1 <= in250 XOR in252;

  Logical_Operator_out255_out1 <= Logical_Operator_out127_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out256_out1 <= in254 XOR in256;

  Logical_Operator_out257_out1 <= Logical_Operator_out129_out1 XOR Logical_Operator_out131_out1;

  Logical_Operator_out258_out1 <= Logical_Operator_out130_out1 XOR Logical_Operator_out132_out1;

  Logical_Operator_out259_out1 <= Logical_Operator_out2_out1 XOR Logical_Operator_out4_out1;

  Logical_Operator_out260_out1 <= in4 XOR in8;

  Logical_Operator_out261_out1 <= Logical_Operator_out133_out1 XOR Logical_Operator_out135_out1;

  Logical_Operator_out262_out1 <= Logical_Operator_out134_out1 XOR Logical_Operator_out136_out1;

  Logical_Operator_out263_out1 <= Logical_Operator_out6_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out264_out1 <= in12 XOR in16;

  Logical_Operator_out265_out1 <= Logical_Operator_out137_out1 XOR Logical_Operator_out139_out1;

  Logical_Operator_out266_out1 <= Logical_Operator_out138_out1 XOR Logical_Operator_out140_out1;

  Logical_Operator_out267_out1 <= Logical_Operator_out10_out1 XOR Logical_Operator_out12_out1;

  Logical_Operator_out268_out1 <= in20 XOR in24;

  Logical_Operator_out269_out1 <= Logical_Operator_out141_out1 XOR Logical_Operator_out143_out1;

  Logical_Operator_out270_out1 <= Logical_Operator_out142_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out271_out1 <= Logical_Operator_out14_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out272_out1 <= in28 XOR in32;

  Logical_Operator_out273_out1 <= Logical_Operator_out145_out1 XOR Logical_Operator_out147_out1;

  Logical_Operator_out274_out1 <= Logical_Operator_out146_out1 XOR Logical_Operator_out148_out1;

  Logical_Operator_out275_out1 <= Logical_Operator_out18_out1 XOR Logical_Operator_out20_out1;

  Logical_Operator_out276_out1 <= in36 XOR in40;

  Logical_Operator_out277_out1 <= Logical_Operator_out149_out1 XOR Logical_Operator_out151_out1;

  Logical_Operator_out278_out1 <= Logical_Operator_out150_out1 XOR Logical_Operator_out152_out1;

  Logical_Operator_out279_out1 <= Logical_Operator_out22_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out280_out1 <= in44 XOR in48;

  Logical_Operator_out281_out1 <= Logical_Operator_out153_out1 XOR Logical_Operator_out155_out1;

  Logical_Operator_out282_out1 <= Logical_Operator_out154_out1 XOR Logical_Operator_out156_out1;

  Logical_Operator_out283_out1 <= Logical_Operator_out26_out1 XOR Logical_Operator_out28_out1;

  Logical_Operator_out284_out1 <= in52 XOR in56;

  Logical_Operator_out285_out1 <= Logical_Operator_out157_out1 XOR Logical_Operator_out159_out1;

  Logical_Operator_out286_out1 <= Logical_Operator_out158_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out287_out1 <= Logical_Operator_out30_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out288_out1 <= in60 XOR in64;

  Logical_Operator_out289_out1 <= Logical_Operator_out161_out1 XOR Logical_Operator_out163_out1;

  Logical_Operator_out290_out1 <= Logical_Operator_out162_out1 XOR Logical_Operator_out164_out1;

  Logical_Operator_out291_out1 <= Logical_Operator_out34_out1 XOR Logical_Operator_out36_out1;

  Logical_Operator_out292_out1 <= in68 XOR in72;

  Logical_Operator_out293_out1 <= Logical_Operator_out165_out1 XOR Logical_Operator_out167_out1;

  Logical_Operator_out294_out1 <= Logical_Operator_out166_out1 XOR Logical_Operator_out168_out1;

  Logical_Operator_out295_out1 <= Logical_Operator_out38_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out296_out1 <= in76 XOR in80;

  Logical_Operator_out297_out1 <= Logical_Operator_out169_out1 XOR Logical_Operator_out171_out1;

  Logical_Operator_out298_out1 <= Logical_Operator_out170_out1 XOR Logical_Operator_out172_out1;

  Logical_Operator_out299_out1 <= Logical_Operator_out42_out1 XOR Logical_Operator_out44_out1;

  Logical_Operator_out300_out1 <= in84 XOR in88;

  Logical_Operator_out301_out1 <= Logical_Operator_out173_out1 XOR Logical_Operator_out175_out1;

  Logical_Operator_out302_out1 <= Logical_Operator_out174_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out303_out1 <= Logical_Operator_out46_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out304_out1 <= in92 XOR in96;

  Logical_Operator_out305_out1 <= Logical_Operator_out177_out1 XOR Logical_Operator_out179_out1;

  Logical_Operator_out306_out1 <= Logical_Operator_out178_out1 XOR Logical_Operator_out180_out1;

  Logical_Operator_out307_out1 <= Logical_Operator_out50_out1 XOR Logical_Operator_out52_out1;

  Logical_Operator_out308_out1 <= in100 XOR in104;

  Logical_Operator_out309_out1 <= Logical_Operator_out181_out1 XOR Logical_Operator_out183_out1;

  Logical_Operator_out310_out1 <= Logical_Operator_out182_out1 XOR Logical_Operator_out184_out1;

  Logical_Operator_out311_out1 <= Logical_Operator_out54_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out312_out1 <= in108 XOR in112;

  Logical_Operator_out313_out1 <= Logical_Operator_out185_out1 XOR Logical_Operator_out187_out1;

  Logical_Operator_out314_out1 <= Logical_Operator_out186_out1 XOR Logical_Operator_out188_out1;

  Logical_Operator_out315_out1 <= Logical_Operator_out58_out1 XOR Logical_Operator_out60_out1;

  Logical_Operator_out316_out1 <= in116 XOR in120;

  Logical_Operator_out317_out1 <= Logical_Operator_out189_out1 XOR Logical_Operator_out191_out1;

  Logical_Operator_out318_out1 <= Logical_Operator_out190_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out319_out1 <= Logical_Operator_out62_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out320_out1 <= in124 XOR in128;

  Logical_Operator_out321_out1 <= Logical_Operator_out193_out1 XOR Logical_Operator_out195_out1;

  Logical_Operator_out322_out1 <= Logical_Operator_out194_out1 XOR Logical_Operator_out196_out1;

  Logical_Operator_out323_out1 <= Logical_Operator_out66_out1 XOR Logical_Operator_out68_out1;

  Logical_Operator_out324_out1 <= in132 XOR in136;

  Logical_Operator_out325_out1 <= Logical_Operator_out197_out1 XOR Logical_Operator_out199_out1;

  Logical_Operator_out326_out1 <= Logical_Operator_out198_out1 XOR Logical_Operator_out200_out1;

  Logical_Operator_out327_out1 <= Logical_Operator_out70_out1 XOR Logical_Operator_out72_out1;

  Logical_Operator_out328_out1 <= in140 XOR in144;

  Logical_Operator_out329_out1 <= Logical_Operator_out201_out1 XOR Logical_Operator_out203_out1;

  Logical_Operator_out330_out1 <= Logical_Operator_out202_out1 XOR Logical_Operator_out204_out1;

  Logical_Operator_out331_out1 <= Logical_Operator_out74_out1 XOR Logical_Operator_out76_out1;

  Logical_Operator_out332_out1 <= in148 XOR in152;

  Logical_Operator_out333_out1 <= Logical_Operator_out205_out1 XOR Logical_Operator_out207_out1;

  Logical_Operator_out334_out1 <= Logical_Operator_out206_out1 XOR Logical_Operator_out208_out1;

  Logical_Operator_out335_out1 <= Logical_Operator_out78_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out336_out1 <= in156 XOR in160;

  Logical_Operator_out337_out1 <= Logical_Operator_out209_out1 XOR Logical_Operator_out211_out1;

  Logical_Operator_out338_out1 <= Logical_Operator_out210_out1 XOR Logical_Operator_out212_out1;

  Logical_Operator_out339_out1 <= Logical_Operator_out82_out1 XOR Logical_Operator_out84_out1;

  Logical_Operator_out340_out1 <= in164 XOR in168;

  Logical_Operator_out341_out1 <= Logical_Operator_out213_out1 XOR Logical_Operator_out215_out1;

  Logical_Operator_out342_out1 <= Logical_Operator_out214_out1 XOR Logical_Operator_out216_out1;

  Logical_Operator_out343_out1 <= Logical_Operator_out86_out1 XOR Logical_Operator_out88_out1;

  Logical_Operator_out344_out1 <= in172 XOR in176;

  Logical_Operator_out345_out1 <= Logical_Operator_out217_out1 XOR Logical_Operator_out219_out1;

  Logical_Operator_out346_out1 <= Logical_Operator_out218_out1 XOR Logical_Operator_out220_out1;

  Logical_Operator_out347_out1 <= Logical_Operator_out90_out1 XOR Logical_Operator_out92_out1;

  Logical_Operator_out348_out1 <= in180 XOR in184;

  Logical_Operator_out349_out1 <= Logical_Operator_out221_out1 XOR Logical_Operator_out223_out1;

  Logical_Operator_out350_out1 <= Logical_Operator_out222_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out351_out1 <= Logical_Operator_out94_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out352_out1 <= in188 XOR in192;

  Logical_Operator_out353_out1 <= Logical_Operator_out225_out1 XOR Logical_Operator_out227_out1;

  Logical_Operator_out354_out1 <= Logical_Operator_out226_out1 XOR Logical_Operator_out228_out1;

  Logical_Operator_out355_out1 <= Logical_Operator_out98_out1 XOR Logical_Operator_out100_out1;

  Logical_Operator_out356_out1 <= in196 XOR in200;

  Logical_Operator_out357_out1 <= Logical_Operator_out229_out1 XOR Logical_Operator_out231_out1;

  Logical_Operator_out358_out1 <= Logical_Operator_out230_out1 XOR Logical_Operator_out232_out1;

  Logical_Operator_out359_out1 <= Logical_Operator_out102_out1 XOR Logical_Operator_out104_out1;

  Logical_Operator_out360_out1 <= in204 XOR in208;

  Logical_Operator_out361_out1 <= Logical_Operator_out233_out1 XOR Logical_Operator_out235_out1;

  Logical_Operator_out362_out1 <= Logical_Operator_out234_out1 XOR Logical_Operator_out236_out1;

  Logical_Operator_out363_out1 <= Logical_Operator_out106_out1 XOR Logical_Operator_out108_out1;

  Logical_Operator_out364_out1 <= in212 XOR in216;

  Logical_Operator_out365_out1 <= Logical_Operator_out237_out1 XOR Logical_Operator_out239_out1;

  Logical_Operator_out366_out1 <= Logical_Operator_out238_out1 XOR Logical_Operator_out240_out1;

  Logical_Operator_out367_out1 <= Logical_Operator_out110_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out368_out1 <= in220 XOR in224;

  Logical_Operator_out369_out1 <= Logical_Operator_out241_out1 XOR Logical_Operator_out243_out1;

  Logical_Operator_out370_out1 <= Logical_Operator_out242_out1 XOR Logical_Operator_out244_out1;

  Logical_Operator_out371_out1 <= Logical_Operator_out114_out1 XOR Logical_Operator_out116_out1;

  Logical_Operator_out372_out1 <= in228 XOR in232;

  Logical_Operator_out373_out1 <= Logical_Operator_out245_out1 XOR Logical_Operator_out247_out1;

  Logical_Operator_out374_out1 <= Logical_Operator_out246_out1 XOR Logical_Operator_out248_out1;

  Logical_Operator_out375_out1 <= Logical_Operator_out118_out1 XOR Logical_Operator_out120_out1;

  Logical_Operator_out376_out1 <= in236 XOR in240;

  Logical_Operator_out377_out1 <= Logical_Operator_out249_out1 XOR Logical_Operator_out251_out1;

  Logical_Operator_out378_out1 <= Logical_Operator_out250_out1 XOR Logical_Operator_out252_out1;

  Logical_Operator_out379_out1 <= Logical_Operator_out122_out1 XOR Logical_Operator_out124_out1;

  Logical_Operator_out380_out1 <= in244 XOR in248;

  Logical_Operator_out381_out1 <= Logical_Operator_out253_out1 XOR Logical_Operator_out255_out1;

  Logical_Operator_out382_out1 <= Logical_Operator_out254_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out383_out1 <= Logical_Operator_out126_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out384_out1 <= in252 XOR in256;

  Logical_Operator_out385_out1 <= Logical_Operator_out257_out1 XOR Logical_Operator_out261_out1;

  Logical_Operator_out386_out1 <= Logical_Operator_out258_out1 XOR Logical_Operator_out262_out1;

  Logical_Operator_out387_out1 <= Logical_Operator_out259_out1 XOR Logical_Operator_out263_out1;

  Logical_Operator_out388_out1 <= Logical_Operator_out260_out1 XOR Logical_Operator_out264_out1;

  Logical_Operator_out389_out1 <= Logical_Operator_out131_out1 XOR Logical_Operator_out135_out1;

  Logical_Operator_out390_out1 <= Logical_Operator_out132_out1 XOR Logical_Operator_out136_out1;

  Logical_Operator_out391_out1 <= Logical_Operator_out4_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out392_out1 <= in8 XOR in16;

  Logical_Operator_out393_out1 <= Logical_Operator_out265_out1 XOR Logical_Operator_out269_out1;

  Logical_Operator_out394_out1 <= Logical_Operator_out266_out1 XOR Logical_Operator_out270_out1;

  Logical_Operator_out395_out1 <= Logical_Operator_out267_out1 XOR Logical_Operator_out271_out1;

  Logical_Operator_out396_out1 <= Logical_Operator_out268_out1 XOR Logical_Operator_out272_out1;

  Logical_Operator_out397_out1 <= Logical_Operator_out139_out1 XOR Logical_Operator_out143_out1;

  Logical_Operator_out398_out1 <= Logical_Operator_out140_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out399_out1 <= Logical_Operator_out12_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out400_out1 <= in24 XOR in32;

  Logical_Operator_out401_out1 <= Logical_Operator_out273_out1 XOR Logical_Operator_out277_out1;

  Logical_Operator_out402_out1 <= Logical_Operator_out274_out1 XOR Logical_Operator_out278_out1;

  Logical_Operator_out403_out1 <= Logical_Operator_out275_out1 XOR Logical_Operator_out279_out1;

  Logical_Operator_out404_out1 <= Logical_Operator_out276_out1 XOR Logical_Operator_out280_out1;

  Logical_Operator_out405_out1 <= Logical_Operator_out147_out1 XOR Logical_Operator_out151_out1;

  Logical_Operator_out406_out1 <= Logical_Operator_out148_out1 XOR Logical_Operator_out152_out1;

  Logical_Operator_out407_out1 <= Logical_Operator_out20_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out408_out1 <= in40 XOR in48;

  Logical_Operator_out409_out1 <= Logical_Operator_out281_out1 XOR Logical_Operator_out285_out1;

  Logical_Operator_out410_out1 <= Logical_Operator_out282_out1 XOR Logical_Operator_out286_out1;

  Logical_Operator_out411_out1 <= Logical_Operator_out283_out1 XOR Logical_Operator_out287_out1;

  Logical_Operator_out412_out1 <= Logical_Operator_out284_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out413_out1 <= Logical_Operator_out155_out1 XOR Logical_Operator_out159_out1;

  Logical_Operator_out414_out1 <= Logical_Operator_out156_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out415_out1 <= Logical_Operator_out28_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out416_out1 <= in56 XOR in64;

  Logical_Operator_out417_out1 <= Logical_Operator_out289_out1 XOR Logical_Operator_out293_out1;

  Logical_Operator_out418_out1 <= Logical_Operator_out290_out1 XOR Logical_Operator_out294_out1;

  Logical_Operator_out419_out1 <= Logical_Operator_out291_out1 XOR Logical_Operator_out295_out1;

  Logical_Operator_out420_out1 <= Logical_Operator_out292_out1 XOR Logical_Operator_out296_out1;

  Logical_Operator_out421_out1 <= Logical_Operator_out163_out1 XOR Logical_Operator_out167_out1;

  Logical_Operator_out422_out1 <= Logical_Operator_out164_out1 XOR Logical_Operator_out168_out1;

  Logical_Operator_out423_out1 <= Logical_Operator_out36_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out424_out1 <= in72 XOR in80;

  Logical_Operator_out425_out1 <= Logical_Operator_out297_out1 XOR Logical_Operator_out301_out1;

  Logical_Operator_out426_out1 <= Logical_Operator_out298_out1 XOR Logical_Operator_out302_out1;

  Logical_Operator_out427_out1 <= Logical_Operator_out299_out1 XOR Logical_Operator_out303_out1;

  Logical_Operator_out428_out1 <= Logical_Operator_out300_out1 XOR Logical_Operator_out304_out1;

  Logical_Operator_out429_out1 <= Logical_Operator_out171_out1 XOR Logical_Operator_out175_out1;

  Logical_Operator_out430_out1 <= Logical_Operator_out172_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out431_out1 <= Logical_Operator_out44_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out432_out1 <= in88 XOR in96;

  Logical_Operator_out433_out1 <= Logical_Operator_out305_out1 XOR Logical_Operator_out309_out1;

  Logical_Operator_out434_out1 <= Logical_Operator_out306_out1 XOR Logical_Operator_out310_out1;

  Logical_Operator_out435_out1 <= Logical_Operator_out307_out1 XOR Logical_Operator_out311_out1;

  Logical_Operator_out436_out1 <= Logical_Operator_out308_out1 XOR Logical_Operator_out312_out1;

  Logical_Operator_out437_out1 <= Logical_Operator_out179_out1 XOR Logical_Operator_out183_out1;

  Logical_Operator_out438_out1 <= Logical_Operator_out180_out1 XOR Logical_Operator_out184_out1;

  Logical_Operator_out439_out1 <= Logical_Operator_out52_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out440_out1 <= in104 XOR in112;

  Logical_Operator_out441_out1 <= Logical_Operator_out313_out1 XOR Logical_Operator_out317_out1;

  Logical_Operator_out442_out1 <= Logical_Operator_out314_out1 XOR Logical_Operator_out318_out1;

  Logical_Operator_out443_out1 <= Logical_Operator_out315_out1 XOR Logical_Operator_out319_out1;

  Logical_Operator_out444_out1 <= Logical_Operator_out316_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out445_out1 <= Logical_Operator_out187_out1 XOR Logical_Operator_out191_out1;

  Logical_Operator_out446_out1 <= Logical_Operator_out188_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out447_out1 <= Logical_Operator_out60_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out448_out1 <= in120 XOR in128;

  Logical_Operator_out449_out1 <= Logical_Operator_out321_out1 XOR Logical_Operator_out325_out1;

  Logical_Operator_out450_out1 <= Logical_Operator_out322_out1 XOR Logical_Operator_out326_out1;

  Logical_Operator_out451_out1 <= Logical_Operator_out323_out1 XOR Logical_Operator_out327_out1;

  Logical_Operator_out452_out1 <= Logical_Operator_out324_out1 XOR Logical_Operator_out328_out1;

  Logical_Operator_out453_out1 <= Logical_Operator_out195_out1 XOR Logical_Operator_out199_out1;

  Logical_Operator_out454_out1 <= Logical_Operator_out196_out1 XOR Logical_Operator_out200_out1;

  Logical_Operator_out455_out1 <= Logical_Operator_out68_out1 XOR Logical_Operator_out72_out1;

  Logical_Operator_out456_out1 <= in136 XOR in144;

  Logical_Operator_out457_out1 <= Logical_Operator_out329_out1 XOR Logical_Operator_out333_out1;

  Logical_Operator_out458_out1 <= Logical_Operator_out330_out1 XOR Logical_Operator_out334_out1;

  Logical_Operator_out459_out1 <= Logical_Operator_out331_out1 XOR Logical_Operator_out335_out1;

  Logical_Operator_out460_out1 <= Logical_Operator_out332_out1 XOR Logical_Operator_out336_out1;

  Logical_Operator_out461_out1 <= Logical_Operator_out203_out1 XOR Logical_Operator_out207_out1;

  Logical_Operator_out462_out1 <= Logical_Operator_out204_out1 XOR Logical_Operator_out208_out1;

  Logical_Operator_out463_out1 <= Logical_Operator_out76_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out464_out1 <= in152 XOR in160;

  Logical_Operator_out465_out1 <= Logical_Operator_out337_out1 XOR Logical_Operator_out341_out1;

  Logical_Operator_out466_out1 <= Logical_Operator_out338_out1 XOR Logical_Operator_out342_out1;

  Logical_Operator_out467_out1 <= Logical_Operator_out339_out1 XOR Logical_Operator_out343_out1;

  Logical_Operator_out468_out1 <= Logical_Operator_out340_out1 XOR Logical_Operator_out344_out1;

  Logical_Operator_out469_out1 <= Logical_Operator_out211_out1 XOR Logical_Operator_out215_out1;

  Logical_Operator_out470_out1 <= Logical_Operator_out212_out1 XOR Logical_Operator_out216_out1;

  Logical_Operator_out471_out1 <= Logical_Operator_out84_out1 XOR Logical_Operator_out88_out1;

  Logical_Operator_out472_out1 <= in168 XOR in176;

  Logical_Operator_out473_out1 <= Logical_Operator_out345_out1 XOR Logical_Operator_out349_out1;

  Logical_Operator_out474_out1 <= Logical_Operator_out346_out1 XOR Logical_Operator_out350_out1;

  Logical_Operator_out475_out1 <= Logical_Operator_out347_out1 XOR Logical_Operator_out351_out1;

  Logical_Operator_out476_out1 <= Logical_Operator_out348_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out477_out1 <= Logical_Operator_out219_out1 XOR Logical_Operator_out223_out1;

  Logical_Operator_out478_out1 <= Logical_Operator_out220_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out479_out1 <= Logical_Operator_out92_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out480_out1 <= in184 XOR in192;

  Logical_Operator_out481_out1 <= Logical_Operator_out353_out1 XOR Logical_Operator_out357_out1;

  Logical_Operator_out482_out1 <= Logical_Operator_out354_out1 XOR Logical_Operator_out358_out1;

  Logical_Operator_out483_out1 <= Logical_Operator_out355_out1 XOR Logical_Operator_out359_out1;

  Logical_Operator_out484_out1 <= Logical_Operator_out356_out1 XOR Logical_Operator_out360_out1;

  Logical_Operator_out485_out1 <= Logical_Operator_out227_out1 XOR Logical_Operator_out231_out1;

  Logical_Operator_out486_out1 <= Logical_Operator_out228_out1 XOR Logical_Operator_out232_out1;

  Logical_Operator_out487_out1 <= Logical_Operator_out100_out1 XOR Logical_Operator_out104_out1;

  Logical_Operator_out488_out1 <= in200 XOR in208;

  Logical_Operator_out489_out1 <= Logical_Operator_out361_out1 XOR Logical_Operator_out365_out1;

  Logical_Operator_out490_out1 <= Logical_Operator_out362_out1 XOR Logical_Operator_out366_out1;

  Logical_Operator_out491_out1 <= Logical_Operator_out363_out1 XOR Logical_Operator_out367_out1;

  Logical_Operator_out492_out1 <= Logical_Operator_out364_out1 XOR Logical_Operator_out368_out1;

  Logical_Operator_out493_out1 <= Logical_Operator_out235_out1 XOR Logical_Operator_out239_out1;

  Logical_Operator_out494_out1 <= Logical_Operator_out236_out1 XOR Logical_Operator_out240_out1;

  Logical_Operator_out495_out1 <= Logical_Operator_out108_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out496_out1 <= in216 XOR in224;

  Logical_Operator_out497_out1 <= Logical_Operator_out369_out1 XOR Logical_Operator_out373_out1;

  Logical_Operator_out498_out1 <= Logical_Operator_out370_out1 XOR Logical_Operator_out374_out1;

  Logical_Operator_out499_out1 <= Logical_Operator_out371_out1 XOR Logical_Operator_out375_out1;

  Logical_Operator_out500_out1 <= Logical_Operator_out372_out1 XOR Logical_Operator_out376_out1;

  Logical_Operator_out501_out1 <= Logical_Operator_out243_out1 XOR Logical_Operator_out247_out1;

  Logical_Operator_out502_out1 <= Logical_Operator_out244_out1 XOR Logical_Operator_out248_out1;

  Logical_Operator_out503_out1 <= Logical_Operator_out116_out1 XOR Logical_Operator_out120_out1;

  Logical_Operator_out504_out1 <= in232 XOR in240;

  Logical_Operator_out505_out1 <= Logical_Operator_out377_out1 XOR Logical_Operator_out381_out1;

  Logical_Operator_out506_out1 <= Logical_Operator_out378_out1 XOR Logical_Operator_out382_out1;

  Logical_Operator_out507_out1 <= Logical_Operator_out379_out1 XOR Logical_Operator_out383_out1;

  Logical_Operator_out508_out1 <= Logical_Operator_out380_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out509_out1 <= Logical_Operator_out251_out1 XOR Logical_Operator_out255_out1;

  Logical_Operator_out510_out1 <= Logical_Operator_out252_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out511_out1 <= Logical_Operator_out124_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out512_out1 <= in248 XOR in256;

  Logical_Operator_out513_out1 <= Logical_Operator_out385_out1 XOR Logical_Operator_out393_out1;

  Logical_Operator_out514_out1 <= Logical_Operator_out386_out1 XOR Logical_Operator_out394_out1;

  Logical_Operator_out515_out1 <= Logical_Operator_out387_out1 XOR Logical_Operator_out395_out1;

  Logical_Operator_out516_out1 <= Logical_Operator_out388_out1 XOR Logical_Operator_out396_out1;

  Logical_Operator_out517_out1 <= Logical_Operator_out389_out1 XOR Logical_Operator_out397_out1;

  Logical_Operator_out518_out1 <= Logical_Operator_out390_out1 XOR Logical_Operator_out398_out1;

  Logical_Operator_out519_out1 <= Logical_Operator_out391_out1 XOR Logical_Operator_out399_out1;

  Logical_Operator_out520_out1 <= Logical_Operator_out392_out1 XOR Logical_Operator_out400_out1;

  Logical_Operator_out521_out1 <= Logical_Operator_out261_out1 XOR Logical_Operator_out269_out1;

  Logical_Operator_out522_out1 <= Logical_Operator_out262_out1 XOR Logical_Operator_out270_out1;

  Logical_Operator_out523_out1 <= Logical_Operator_out263_out1 XOR Logical_Operator_out271_out1;

  Logical_Operator_out524_out1 <= Logical_Operator_out264_out1 XOR Logical_Operator_out272_out1;

  Logical_Operator_out525_out1 <= Logical_Operator_out135_out1 XOR Logical_Operator_out143_out1;

  Logical_Operator_out526_out1 <= Logical_Operator_out136_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out527_out1 <= Logical_Operator_out8_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out528_out1 <= in16 XOR in32;

  Logical_Operator_out529_out1 <= Logical_Operator_out401_out1 XOR Logical_Operator_out409_out1;

  Logical_Operator_out530_out1 <= Logical_Operator_out402_out1 XOR Logical_Operator_out410_out1;

  Logical_Operator_out531_out1 <= Logical_Operator_out403_out1 XOR Logical_Operator_out411_out1;

  Logical_Operator_out532_out1 <= Logical_Operator_out404_out1 XOR Logical_Operator_out412_out1;

  Logical_Operator_out533_out1 <= Logical_Operator_out405_out1 XOR Logical_Operator_out413_out1;

  Logical_Operator_out534_out1 <= Logical_Operator_out406_out1 XOR Logical_Operator_out414_out1;

  Logical_Operator_out535_out1 <= Logical_Operator_out407_out1 XOR Logical_Operator_out415_out1;

  Logical_Operator_out536_out1 <= Logical_Operator_out408_out1 XOR Logical_Operator_out416_out1;

  Logical_Operator_out537_out1 <= Logical_Operator_out277_out1 XOR Logical_Operator_out285_out1;

  Logical_Operator_out538_out1 <= Logical_Operator_out278_out1 XOR Logical_Operator_out286_out1;

  Logical_Operator_out539_out1 <= Logical_Operator_out279_out1 XOR Logical_Operator_out287_out1;

  Logical_Operator_out540_out1 <= Logical_Operator_out280_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out541_out1 <= Logical_Operator_out151_out1 XOR Logical_Operator_out159_out1;

  Logical_Operator_out542_out1 <= Logical_Operator_out152_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out543_out1 <= Logical_Operator_out24_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out544_out1 <= in48 XOR in64;

  Logical_Operator_out545_out1 <= Logical_Operator_out417_out1 XOR Logical_Operator_out425_out1;

  Logical_Operator_out546_out1 <= Logical_Operator_out418_out1 XOR Logical_Operator_out426_out1;

  Logical_Operator_out547_out1 <= Logical_Operator_out419_out1 XOR Logical_Operator_out427_out1;

  Logical_Operator_out548_out1 <= Logical_Operator_out420_out1 XOR Logical_Operator_out428_out1;

  Logical_Operator_out549_out1 <= Logical_Operator_out421_out1 XOR Logical_Operator_out429_out1;

  Logical_Operator_out550_out1 <= Logical_Operator_out422_out1 XOR Logical_Operator_out430_out1;

  Logical_Operator_out551_out1 <= Logical_Operator_out423_out1 XOR Logical_Operator_out431_out1;

  Logical_Operator_out552_out1 <= Logical_Operator_out424_out1 XOR Logical_Operator_out432_out1;

  Logical_Operator_out553_out1 <= Logical_Operator_out293_out1 XOR Logical_Operator_out301_out1;

  Logical_Operator_out554_out1 <= Logical_Operator_out294_out1 XOR Logical_Operator_out302_out1;

  Logical_Operator_out555_out1 <= Logical_Operator_out295_out1 XOR Logical_Operator_out303_out1;

  Logical_Operator_out556_out1 <= Logical_Operator_out296_out1 XOR Logical_Operator_out304_out1;

  Logical_Operator_out557_out1 <= Logical_Operator_out167_out1 XOR Logical_Operator_out175_out1;

  Logical_Operator_out558_out1 <= Logical_Operator_out168_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out559_out1 <= Logical_Operator_out40_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out560_out1 <= in80 XOR in96;

  Logical_Operator_out561_out1 <= Logical_Operator_out433_out1 XOR Logical_Operator_out441_out1;

  Logical_Operator_out562_out1 <= Logical_Operator_out434_out1 XOR Logical_Operator_out442_out1;

  Logical_Operator_out563_out1 <= Logical_Operator_out435_out1 XOR Logical_Operator_out443_out1;

  Logical_Operator_out564_out1 <= Logical_Operator_out436_out1 XOR Logical_Operator_out444_out1;

  Logical_Operator_out565_out1 <= Logical_Operator_out437_out1 XOR Logical_Operator_out445_out1;

  Logical_Operator_out566_out1 <= Logical_Operator_out438_out1 XOR Logical_Operator_out446_out1;

  Logical_Operator_out567_out1 <= Logical_Operator_out439_out1 XOR Logical_Operator_out447_out1;

  Logical_Operator_out568_out1 <= Logical_Operator_out440_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out569_out1 <= Logical_Operator_out309_out1 XOR Logical_Operator_out317_out1;

  Logical_Operator_out570_out1 <= Logical_Operator_out310_out1 XOR Logical_Operator_out318_out1;

  Logical_Operator_out571_out1 <= Logical_Operator_out311_out1 XOR Logical_Operator_out319_out1;

  Logical_Operator_out572_out1 <= Logical_Operator_out312_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out573_out1 <= Logical_Operator_out183_out1 XOR Logical_Operator_out191_out1;

  Logical_Operator_out574_out1 <= Logical_Operator_out184_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out575_out1 <= Logical_Operator_out56_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out576_out1 <= in112 XOR in128;

  Logical_Operator_out577_out1 <= Logical_Operator_out449_out1 XOR Logical_Operator_out457_out1;

  Logical_Operator_out578_out1 <= Logical_Operator_out450_out1 XOR Logical_Operator_out458_out1;

  Logical_Operator_out579_out1 <= Logical_Operator_out451_out1 XOR Logical_Operator_out459_out1;

  Logical_Operator_out580_out1 <= Logical_Operator_out452_out1 XOR Logical_Operator_out460_out1;

  Logical_Operator_out581_out1 <= Logical_Operator_out453_out1 XOR Logical_Operator_out461_out1;

  Logical_Operator_out582_out1 <= Logical_Operator_out454_out1 XOR Logical_Operator_out462_out1;

  Logical_Operator_out583_out1 <= Logical_Operator_out455_out1 XOR Logical_Operator_out463_out1;

  Logical_Operator_out584_out1 <= Logical_Operator_out456_out1 XOR Logical_Operator_out464_out1;

  Logical_Operator_out585_out1 <= Logical_Operator_out325_out1 XOR Logical_Operator_out333_out1;

  Logical_Operator_out586_out1 <= Logical_Operator_out326_out1 XOR Logical_Operator_out334_out1;

  Logical_Operator_out587_out1 <= Logical_Operator_out327_out1 XOR Logical_Operator_out335_out1;

  Logical_Operator_out588_out1 <= Logical_Operator_out328_out1 XOR Logical_Operator_out336_out1;

  Logical_Operator_out589_out1 <= Logical_Operator_out199_out1 XOR Logical_Operator_out207_out1;

  Logical_Operator_out590_out1 <= Logical_Operator_out200_out1 XOR Logical_Operator_out208_out1;

  Logical_Operator_out591_out1 <= Logical_Operator_out72_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out592_out1 <= in144 XOR in160;

  Logical_Operator_out593_out1 <= Logical_Operator_out465_out1 XOR Logical_Operator_out473_out1;

  Logical_Operator_out594_out1 <= Logical_Operator_out466_out1 XOR Logical_Operator_out474_out1;

  Logical_Operator_out595_out1 <= Logical_Operator_out467_out1 XOR Logical_Operator_out475_out1;

  Logical_Operator_out596_out1 <= Logical_Operator_out468_out1 XOR Logical_Operator_out476_out1;

  Logical_Operator_out597_out1 <= Logical_Operator_out469_out1 XOR Logical_Operator_out477_out1;

  Logical_Operator_out598_out1 <= Logical_Operator_out470_out1 XOR Logical_Operator_out478_out1;

  Logical_Operator_out599_out1 <= Logical_Operator_out471_out1 XOR Logical_Operator_out479_out1;

  Logical_Operator_out600_out1 <= Logical_Operator_out472_out1 XOR Logical_Operator_out480_out1;

  Logical_Operator_out601_out1 <= Logical_Operator_out341_out1 XOR Logical_Operator_out349_out1;

  Logical_Operator_out602_out1 <= Logical_Operator_out342_out1 XOR Logical_Operator_out350_out1;

  Logical_Operator_out603_out1 <= Logical_Operator_out343_out1 XOR Logical_Operator_out351_out1;

  Logical_Operator_out604_out1 <= Logical_Operator_out344_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out605_out1 <= Logical_Operator_out215_out1 XOR Logical_Operator_out223_out1;

  Logical_Operator_out606_out1 <= Logical_Operator_out216_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out607_out1 <= Logical_Operator_out88_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out608_out1 <= in176 XOR in192;

  Logical_Operator_out609_out1 <= Logical_Operator_out481_out1 XOR Logical_Operator_out489_out1;

  Logical_Operator_out610_out1 <= Logical_Operator_out482_out1 XOR Logical_Operator_out490_out1;

  Logical_Operator_out611_out1 <= Logical_Operator_out483_out1 XOR Logical_Operator_out491_out1;

  Logical_Operator_out612_out1 <= Logical_Operator_out484_out1 XOR Logical_Operator_out492_out1;

  Logical_Operator_out613_out1 <= Logical_Operator_out485_out1 XOR Logical_Operator_out493_out1;

  Logical_Operator_out614_out1 <= Logical_Operator_out486_out1 XOR Logical_Operator_out494_out1;

  Logical_Operator_out615_out1 <= Logical_Operator_out487_out1 XOR Logical_Operator_out495_out1;

  Logical_Operator_out616_out1 <= Logical_Operator_out488_out1 XOR Logical_Operator_out496_out1;

  Logical_Operator_out617_out1 <= Logical_Operator_out357_out1 XOR Logical_Operator_out365_out1;

  Logical_Operator_out618_out1 <= Logical_Operator_out358_out1 XOR Logical_Operator_out366_out1;

  Logical_Operator_out619_out1 <= Logical_Operator_out359_out1 XOR Logical_Operator_out367_out1;

  Logical_Operator_out620_out1 <= Logical_Operator_out360_out1 XOR Logical_Operator_out368_out1;

  Logical_Operator_out621_out1 <= Logical_Operator_out231_out1 XOR Logical_Operator_out239_out1;

  Logical_Operator_out622_out1 <= Logical_Operator_out232_out1 XOR Logical_Operator_out240_out1;

  Logical_Operator_out623_out1 <= Logical_Operator_out104_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out624_out1 <= in208 XOR in224;

  Logical_Operator_out625_out1 <= Logical_Operator_out497_out1 XOR Logical_Operator_out505_out1;

  Logical_Operator_out626_out1 <= Logical_Operator_out498_out1 XOR Logical_Operator_out506_out1;

  Logical_Operator_out627_out1 <= Logical_Operator_out499_out1 XOR Logical_Operator_out507_out1;

  Logical_Operator_out628_out1 <= Logical_Operator_out500_out1 XOR Logical_Operator_out508_out1;

  Logical_Operator_out629_out1 <= Logical_Operator_out501_out1 XOR Logical_Operator_out509_out1;

  Logical_Operator_out630_out1 <= Logical_Operator_out502_out1 XOR Logical_Operator_out510_out1;

  Logical_Operator_out631_out1 <= Logical_Operator_out503_out1 XOR Logical_Operator_out511_out1;

  Logical_Operator_out632_out1 <= Logical_Operator_out504_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out633_out1 <= Logical_Operator_out373_out1 XOR Logical_Operator_out381_out1;

  Logical_Operator_out634_out1 <= Logical_Operator_out374_out1 XOR Logical_Operator_out382_out1;

  Logical_Operator_out635_out1 <= Logical_Operator_out375_out1 XOR Logical_Operator_out383_out1;

  Logical_Operator_out636_out1 <= Logical_Operator_out376_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out637_out1 <= Logical_Operator_out247_out1 XOR Logical_Operator_out255_out1;

  Logical_Operator_out638_out1 <= Logical_Operator_out248_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out639_out1 <= Logical_Operator_out120_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out640_out1 <= in240 XOR in256;

  Logical_Operator_out641_out1 <= Logical_Operator_out513_out1 XOR Logical_Operator_out529_out1;

  Logical_Operator_out642_out1 <= Logical_Operator_out514_out1 XOR Logical_Operator_out530_out1;

  Logical_Operator_out643_out1 <= Logical_Operator_out515_out1 XOR Logical_Operator_out531_out1;

  Logical_Operator_out644_out1 <= Logical_Operator_out516_out1 XOR Logical_Operator_out532_out1;

  Logical_Operator_out645_out1 <= Logical_Operator_out517_out1 XOR Logical_Operator_out533_out1;

  Logical_Operator_out646_out1 <= Logical_Operator_out518_out1 XOR Logical_Operator_out534_out1;

  Logical_Operator_out647_out1 <= Logical_Operator_out519_out1 XOR Logical_Operator_out535_out1;

  Logical_Operator_out648_out1 <= Logical_Operator_out520_out1 XOR Logical_Operator_out536_out1;

  Logical_Operator_out649_out1 <= Logical_Operator_out521_out1 XOR Logical_Operator_out537_out1;

  Logical_Operator_out650_out1 <= Logical_Operator_out522_out1 XOR Logical_Operator_out538_out1;

  Logical_Operator_out651_out1 <= Logical_Operator_out523_out1 XOR Logical_Operator_out539_out1;

  Logical_Operator_out652_out1 <= Logical_Operator_out524_out1 XOR Logical_Operator_out540_out1;

  Logical_Operator_out653_out1 <= Logical_Operator_out525_out1 XOR Logical_Operator_out541_out1;

  Logical_Operator_out654_out1 <= Logical_Operator_out526_out1 XOR Logical_Operator_out542_out1;

  Logical_Operator_out655_out1 <= Logical_Operator_out527_out1 XOR Logical_Operator_out543_out1;

  Logical_Operator_out656_out1 <= Logical_Operator_out528_out1 XOR Logical_Operator_out544_out1;

  Logical_Operator_out657_out1 <= Logical_Operator_out393_out1 XOR Logical_Operator_out409_out1;

  Logical_Operator_out658_out1 <= Logical_Operator_out394_out1 XOR Logical_Operator_out410_out1;

  Logical_Operator_out659_out1 <= Logical_Operator_out395_out1 XOR Logical_Operator_out411_out1;

  Logical_Operator_out660_out1 <= Logical_Operator_out396_out1 XOR Logical_Operator_out412_out1;

  Logical_Operator_out661_out1 <= Logical_Operator_out397_out1 XOR Logical_Operator_out413_out1;

  Logical_Operator_out662_out1 <= Logical_Operator_out398_out1 XOR Logical_Operator_out414_out1;

  Logical_Operator_out663_out1 <= Logical_Operator_out399_out1 XOR Logical_Operator_out415_out1;

  Logical_Operator_out664_out1 <= Logical_Operator_out400_out1 XOR Logical_Operator_out416_out1;

  Logical_Operator_out665_out1 <= Logical_Operator_out269_out1 XOR Logical_Operator_out285_out1;

  Logical_Operator_out666_out1 <= Logical_Operator_out270_out1 XOR Logical_Operator_out286_out1;

  Logical_Operator_out667_out1 <= Logical_Operator_out271_out1 XOR Logical_Operator_out287_out1;

  Logical_Operator_out668_out1 <= Logical_Operator_out272_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out669_out1 <= Logical_Operator_out143_out1 XOR Logical_Operator_out159_out1;

  Logical_Operator_out670_out1 <= Logical_Operator_out144_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out671_out1 <= Logical_Operator_out16_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out672_out1 <= in32 XOR in64;

  Logical_Operator_out673_out1 <= Logical_Operator_out545_out1 XOR Logical_Operator_out561_out1;

  Logical_Operator_out674_out1 <= Logical_Operator_out546_out1 XOR Logical_Operator_out562_out1;

  Logical_Operator_out675_out1 <= Logical_Operator_out547_out1 XOR Logical_Operator_out563_out1;

  Logical_Operator_out676_out1 <= Logical_Operator_out548_out1 XOR Logical_Operator_out564_out1;

  Logical_Operator_out677_out1 <= Logical_Operator_out549_out1 XOR Logical_Operator_out565_out1;

  Logical_Operator_out678_out1 <= Logical_Operator_out550_out1 XOR Logical_Operator_out566_out1;

  Logical_Operator_out679_out1 <= Logical_Operator_out551_out1 XOR Logical_Operator_out567_out1;

  Logical_Operator_out680_out1 <= Logical_Operator_out552_out1 XOR Logical_Operator_out568_out1;

  Logical_Operator_out681_out1 <= Logical_Operator_out553_out1 XOR Logical_Operator_out569_out1;

  Logical_Operator_out682_out1 <= Logical_Operator_out554_out1 XOR Logical_Operator_out570_out1;

  Logical_Operator_out683_out1 <= Logical_Operator_out555_out1 XOR Logical_Operator_out571_out1;

  Logical_Operator_out684_out1 <= Logical_Operator_out556_out1 XOR Logical_Operator_out572_out1;

  Logical_Operator_out685_out1 <= Logical_Operator_out557_out1 XOR Logical_Operator_out573_out1;

  Logical_Operator_out686_out1 <= Logical_Operator_out558_out1 XOR Logical_Operator_out574_out1;

  Logical_Operator_out687_out1 <= Logical_Operator_out559_out1 XOR Logical_Operator_out575_out1;

  Logical_Operator_out688_out1 <= Logical_Operator_out560_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out689_out1 <= Logical_Operator_out425_out1 XOR Logical_Operator_out441_out1;

  Logical_Operator_out690_out1 <= Logical_Operator_out426_out1 XOR Logical_Operator_out442_out1;

  Logical_Operator_out691_out1 <= Logical_Operator_out427_out1 XOR Logical_Operator_out443_out1;

  Logical_Operator_out692_out1 <= Logical_Operator_out428_out1 XOR Logical_Operator_out444_out1;

  Logical_Operator_out693_out1 <= Logical_Operator_out429_out1 XOR Logical_Operator_out445_out1;

  Logical_Operator_out694_out1 <= Logical_Operator_out430_out1 XOR Logical_Operator_out446_out1;

  Logical_Operator_out695_out1 <= Logical_Operator_out431_out1 XOR Logical_Operator_out447_out1;

  Logical_Operator_out696_out1 <= Logical_Operator_out432_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out697_out1 <= Logical_Operator_out301_out1 XOR Logical_Operator_out317_out1;

  Logical_Operator_out698_out1 <= Logical_Operator_out302_out1 XOR Logical_Operator_out318_out1;

  Logical_Operator_out699_out1 <= Logical_Operator_out303_out1 XOR Logical_Operator_out319_out1;

  Logical_Operator_out700_out1 <= Logical_Operator_out304_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out701_out1 <= Logical_Operator_out175_out1 XOR Logical_Operator_out191_out1;

  Logical_Operator_out702_out1 <= Logical_Operator_out176_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out703_out1 <= Logical_Operator_out48_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out704_out1 <= in96 XOR in128;

  Logical_Operator_out705_out1 <= Logical_Operator_out577_out1 XOR Logical_Operator_out593_out1;

  Logical_Operator_out706_out1 <= Logical_Operator_out578_out1 XOR Logical_Operator_out594_out1;

  Logical_Operator_out707_out1 <= Logical_Operator_out579_out1 XOR Logical_Operator_out595_out1;

  Logical_Operator_out708_out1 <= Logical_Operator_out580_out1 XOR Logical_Operator_out596_out1;

  Logical_Operator_out709_out1 <= Logical_Operator_out581_out1 XOR Logical_Operator_out597_out1;

  Logical_Operator_out710_out1 <= Logical_Operator_out582_out1 XOR Logical_Operator_out598_out1;

  Logical_Operator_out711_out1 <= Logical_Operator_out583_out1 XOR Logical_Operator_out599_out1;

  Logical_Operator_out712_out1 <= Logical_Operator_out584_out1 XOR Logical_Operator_out600_out1;

  Logical_Operator_out713_out1 <= Logical_Operator_out585_out1 XOR Logical_Operator_out601_out1;

  Logical_Operator_out714_out1 <= Logical_Operator_out586_out1 XOR Logical_Operator_out602_out1;

  Logical_Operator_out715_out1 <= Logical_Operator_out587_out1 XOR Logical_Operator_out603_out1;

  Logical_Operator_out716_out1 <= Logical_Operator_out588_out1 XOR Logical_Operator_out604_out1;

  Logical_Operator_out717_out1 <= Logical_Operator_out589_out1 XOR Logical_Operator_out605_out1;

  Logical_Operator_out718_out1 <= Logical_Operator_out590_out1 XOR Logical_Operator_out606_out1;

  Logical_Operator_out719_out1 <= Logical_Operator_out591_out1 XOR Logical_Operator_out607_out1;

  Logical_Operator_out720_out1 <= Logical_Operator_out592_out1 XOR Logical_Operator_out608_out1;

  Logical_Operator_out721_out1 <= Logical_Operator_out457_out1 XOR Logical_Operator_out473_out1;

  Logical_Operator_out722_out1 <= Logical_Operator_out458_out1 XOR Logical_Operator_out474_out1;

  Logical_Operator_out723_out1 <= Logical_Operator_out459_out1 XOR Logical_Operator_out475_out1;

  Logical_Operator_out724_out1 <= Logical_Operator_out460_out1 XOR Logical_Operator_out476_out1;

  Logical_Operator_out725_out1 <= Logical_Operator_out461_out1 XOR Logical_Operator_out477_out1;

  Logical_Operator_out726_out1 <= Logical_Operator_out462_out1 XOR Logical_Operator_out478_out1;

  Logical_Operator_out727_out1 <= Logical_Operator_out463_out1 XOR Logical_Operator_out479_out1;

  Logical_Operator_out728_out1 <= Logical_Operator_out464_out1 XOR Logical_Operator_out480_out1;

  Logical_Operator_out729_out1 <= Logical_Operator_out333_out1 XOR Logical_Operator_out349_out1;

  Logical_Operator_out730_out1 <= Logical_Operator_out334_out1 XOR Logical_Operator_out350_out1;

  Logical_Operator_out731_out1 <= Logical_Operator_out335_out1 XOR Logical_Operator_out351_out1;

  Logical_Operator_out732_out1 <= Logical_Operator_out336_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out733_out1 <= Logical_Operator_out207_out1 XOR Logical_Operator_out223_out1;

  Logical_Operator_out734_out1 <= Logical_Operator_out208_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out735_out1 <= Logical_Operator_out80_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out736_out1 <= in160 XOR in192;

  Logical_Operator_out737_out1 <= Logical_Operator_out609_out1 XOR Logical_Operator_out625_out1;

  Logical_Operator_out738_out1 <= Logical_Operator_out610_out1 XOR Logical_Operator_out626_out1;

  Logical_Operator_out739_out1 <= Logical_Operator_out611_out1 XOR Logical_Operator_out627_out1;

  Logical_Operator_out740_out1 <= Logical_Operator_out612_out1 XOR Logical_Operator_out628_out1;

  Logical_Operator_out741_out1 <= Logical_Operator_out613_out1 XOR Logical_Operator_out629_out1;

  Logical_Operator_out742_out1 <= Logical_Operator_out614_out1 XOR Logical_Operator_out630_out1;

  Logical_Operator_out743_out1 <= Logical_Operator_out615_out1 XOR Logical_Operator_out631_out1;

  Logical_Operator_out744_out1 <= Logical_Operator_out616_out1 XOR Logical_Operator_out632_out1;

  Logical_Operator_out745_out1 <= Logical_Operator_out617_out1 XOR Logical_Operator_out633_out1;

  Logical_Operator_out746_out1 <= Logical_Operator_out618_out1 XOR Logical_Operator_out634_out1;

  Logical_Operator_out747_out1 <= Logical_Operator_out619_out1 XOR Logical_Operator_out635_out1;

  Logical_Operator_out748_out1 <= Logical_Operator_out620_out1 XOR Logical_Operator_out636_out1;

  Logical_Operator_out749_out1 <= Logical_Operator_out621_out1 XOR Logical_Operator_out637_out1;

  Logical_Operator_out750_out1 <= Logical_Operator_out622_out1 XOR Logical_Operator_out638_out1;

  Logical_Operator_out751_out1 <= Logical_Operator_out623_out1 XOR Logical_Operator_out639_out1;

  Logical_Operator_out752_out1 <= Logical_Operator_out624_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out753_out1 <= Logical_Operator_out489_out1 XOR Logical_Operator_out505_out1;

  Logical_Operator_out754_out1 <= Logical_Operator_out490_out1 XOR Logical_Operator_out506_out1;

  Logical_Operator_out755_out1 <= Logical_Operator_out491_out1 XOR Logical_Operator_out507_out1;

  Logical_Operator_out756_out1 <= Logical_Operator_out492_out1 XOR Logical_Operator_out508_out1;

  Logical_Operator_out757_out1 <= Logical_Operator_out493_out1 XOR Logical_Operator_out509_out1;

  Logical_Operator_out758_out1 <= Logical_Operator_out494_out1 XOR Logical_Operator_out510_out1;

  Logical_Operator_out759_out1 <= Logical_Operator_out495_out1 XOR Logical_Operator_out511_out1;

  Logical_Operator_out760_out1 <= Logical_Operator_out496_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out761_out1 <= Logical_Operator_out365_out1 XOR Logical_Operator_out381_out1;

  Logical_Operator_out762_out1 <= Logical_Operator_out366_out1 XOR Logical_Operator_out382_out1;

  Logical_Operator_out763_out1 <= Logical_Operator_out367_out1 XOR Logical_Operator_out383_out1;

  Logical_Operator_out764_out1 <= Logical_Operator_out368_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out765_out1 <= Logical_Operator_out239_out1 XOR Logical_Operator_out255_out1;

  Logical_Operator_out766_out1 <= Logical_Operator_out240_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out767_out1 <= Logical_Operator_out112_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out768_out1 <= in224 XOR in256;

  Logical_Operator_out769_out1 <= Logical_Operator_out641_out1 XOR Logical_Operator_out673_out1;

  Logical_Operator_out770_out1 <= Logical_Operator_out642_out1 XOR Logical_Operator_out674_out1;

  Logical_Operator_out771_out1 <= Logical_Operator_out643_out1 XOR Logical_Operator_out675_out1;

  Logical_Operator_out772_out1 <= Logical_Operator_out644_out1 XOR Logical_Operator_out676_out1;

  Logical_Operator_out773_out1 <= Logical_Operator_out645_out1 XOR Logical_Operator_out677_out1;

  Logical_Operator_out774_out1 <= Logical_Operator_out646_out1 XOR Logical_Operator_out678_out1;

  Logical_Operator_out775_out1 <= Logical_Operator_out647_out1 XOR Logical_Operator_out679_out1;

  Logical_Operator_out776_out1 <= Logical_Operator_out648_out1 XOR Logical_Operator_out680_out1;

  Logical_Operator_out777_out1 <= Logical_Operator_out649_out1 XOR Logical_Operator_out681_out1;

  Logical_Operator_out778_out1 <= Logical_Operator_out650_out1 XOR Logical_Operator_out682_out1;

  Logical_Operator_out779_out1 <= Logical_Operator_out651_out1 XOR Logical_Operator_out683_out1;

  Logical_Operator_out780_out1 <= Logical_Operator_out652_out1 XOR Logical_Operator_out684_out1;

  Logical_Operator_out781_out1 <= Logical_Operator_out653_out1 XOR Logical_Operator_out685_out1;

  Logical_Operator_out782_out1 <= Logical_Operator_out654_out1 XOR Logical_Operator_out686_out1;

  Logical_Operator_out783_out1 <= Logical_Operator_out655_out1 XOR Logical_Operator_out687_out1;

  Logical_Operator_out784_out1 <= Logical_Operator_out656_out1 XOR Logical_Operator_out688_out1;

  Logical_Operator_out785_out1 <= Logical_Operator_out657_out1 XOR Logical_Operator_out689_out1;

  Logical_Operator_out786_out1 <= Logical_Operator_out658_out1 XOR Logical_Operator_out690_out1;

  Logical_Operator_out787_out1 <= Logical_Operator_out659_out1 XOR Logical_Operator_out691_out1;

  Logical_Operator_out788_out1 <= Logical_Operator_out660_out1 XOR Logical_Operator_out692_out1;

  Logical_Operator_out789_out1 <= Logical_Operator_out661_out1 XOR Logical_Operator_out693_out1;

  Logical_Operator_out790_out1 <= Logical_Operator_out662_out1 XOR Logical_Operator_out694_out1;

  Logical_Operator_out791_out1 <= Logical_Operator_out663_out1 XOR Logical_Operator_out695_out1;

  Logical_Operator_out792_out1 <= Logical_Operator_out664_out1 XOR Logical_Operator_out696_out1;

  Logical_Operator_out793_out1 <= Logical_Operator_out665_out1 XOR Logical_Operator_out697_out1;

  Logical_Operator_out794_out1 <= Logical_Operator_out666_out1 XOR Logical_Operator_out698_out1;

  Logical_Operator_out795_out1 <= Logical_Operator_out667_out1 XOR Logical_Operator_out699_out1;

  Logical_Operator_out796_out1 <= Logical_Operator_out668_out1 XOR Logical_Operator_out700_out1;

  Logical_Operator_out797_out1 <= Logical_Operator_out669_out1 XOR Logical_Operator_out701_out1;

  Logical_Operator_out798_out1 <= Logical_Operator_out670_out1 XOR Logical_Operator_out702_out1;

  Logical_Operator_out799_out1 <= Logical_Operator_out671_out1 XOR Logical_Operator_out703_out1;

  Logical_Operator_out800_out1 <= Logical_Operator_out672_out1 XOR Logical_Operator_out704_out1;

  Logical_Operator_out801_out1 <= Logical_Operator_out529_out1 XOR Logical_Operator_out561_out1;

  Logical_Operator_out802_out1 <= Logical_Operator_out530_out1 XOR Logical_Operator_out562_out1;

  Logical_Operator_out803_out1 <= Logical_Operator_out531_out1 XOR Logical_Operator_out563_out1;

  Logical_Operator_out804_out1 <= Logical_Operator_out532_out1 XOR Logical_Operator_out564_out1;

  Logical_Operator_out805_out1 <= Logical_Operator_out533_out1 XOR Logical_Operator_out565_out1;

  Logical_Operator_out806_out1 <= Logical_Operator_out534_out1 XOR Logical_Operator_out566_out1;

  Logical_Operator_out807_out1 <= Logical_Operator_out535_out1 XOR Logical_Operator_out567_out1;

  Logical_Operator_out808_out1 <= Logical_Operator_out536_out1 XOR Logical_Operator_out568_out1;

  Logical_Operator_out809_out1 <= Logical_Operator_out537_out1 XOR Logical_Operator_out569_out1;

  Logical_Operator_out810_out1 <= Logical_Operator_out538_out1 XOR Logical_Operator_out570_out1;

  Logical_Operator_out811_out1 <= Logical_Operator_out539_out1 XOR Logical_Operator_out571_out1;

  Logical_Operator_out812_out1 <= Logical_Operator_out540_out1 XOR Logical_Operator_out572_out1;

  Logical_Operator_out813_out1 <= Logical_Operator_out541_out1 XOR Logical_Operator_out573_out1;

  Logical_Operator_out814_out1 <= Logical_Operator_out542_out1 XOR Logical_Operator_out574_out1;

  Logical_Operator_out815_out1 <= Logical_Operator_out543_out1 XOR Logical_Operator_out575_out1;

  Logical_Operator_out816_out1 <= Logical_Operator_out544_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out817_out1 <= Logical_Operator_out409_out1 XOR Logical_Operator_out441_out1;

  Logical_Operator_out818_out1 <= Logical_Operator_out410_out1 XOR Logical_Operator_out442_out1;

  Logical_Operator_out819_out1 <= Logical_Operator_out411_out1 XOR Logical_Operator_out443_out1;

  Logical_Operator_out820_out1 <= Logical_Operator_out412_out1 XOR Logical_Operator_out444_out1;

  Logical_Operator_out821_out1 <= Logical_Operator_out413_out1 XOR Logical_Operator_out445_out1;

  Logical_Operator_out822_out1 <= Logical_Operator_out414_out1 XOR Logical_Operator_out446_out1;

  Logical_Operator_out823_out1 <= Logical_Operator_out415_out1 XOR Logical_Operator_out447_out1;

  Logical_Operator_out824_out1 <= Logical_Operator_out416_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out825_out1 <= Logical_Operator_out285_out1 XOR Logical_Operator_out317_out1;

  Logical_Operator_out826_out1 <= Logical_Operator_out286_out1 XOR Logical_Operator_out318_out1;

  Logical_Operator_out827_out1 <= Logical_Operator_out287_out1 XOR Logical_Operator_out319_out1;

  Logical_Operator_out828_out1 <= Logical_Operator_out288_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out829_out1 <= Logical_Operator_out159_out1 XOR Logical_Operator_out191_out1;

  Logical_Operator_out830_out1 <= Logical_Operator_out160_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out831_out1 <= Logical_Operator_out32_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out832_out1 <= in64 XOR in128;

  Logical_Operator_out833_out1 <= Logical_Operator_out705_out1 XOR Logical_Operator_out737_out1;

  Logical_Operator_out834_out1 <= Logical_Operator_out706_out1 XOR Logical_Operator_out738_out1;

  Logical_Operator_out835_out1 <= Logical_Operator_out707_out1 XOR Logical_Operator_out739_out1;

  Logical_Operator_out836_out1 <= Logical_Operator_out708_out1 XOR Logical_Operator_out740_out1;

  Logical_Operator_out837_out1 <= Logical_Operator_out709_out1 XOR Logical_Operator_out741_out1;

  Logical_Operator_out838_out1 <= Logical_Operator_out710_out1 XOR Logical_Operator_out742_out1;

  Logical_Operator_out839_out1 <= Logical_Operator_out711_out1 XOR Logical_Operator_out743_out1;

  Logical_Operator_out840_out1 <= Logical_Operator_out712_out1 XOR Logical_Operator_out744_out1;

  Logical_Operator_out841_out1 <= Logical_Operator_out713_out1 XOR Logical_Operator_out745_out1;

  Logical_Operator_out842_out1 <= Logical_Operator_out714_out1 XOR Logical_Operator_out746_out1;

  Logical_Operator_out843_out1 <= Logical_Operator_out715_out1 XOR Logical_Operator_out747_out1;

  Logical_Operator_out844_out1 <= Logical_Operator_out716_out1 XOR Logical_Operator_out748_out1;

  Logical_Operator_out845_out1 <= Logical_Operator_out717_out1 XOR Logical_Operator_out749_out1;

  Logical_Operator_out846_out1 <= Logical_Operator_out718_out1 XOR Logical_Operator_out750_out1;

  Logical_Operator_out847_out1 <= Logical_Operator_out719_out1 XOR Logical_Operator_out751_out1;

  Logical_Operator_out848_out1 <= Logical_Operator_out720_out1 XOR Logical_Operator_out752_out1;

  Logical_Operator_out849_out1 <= Logical_Operator_out721_out1 XOR Logical_Operator_out753_out1;

  Logical_Operator_out850_out1 <= Logical_Operator_out722_out1 XOR Logical_Operator_out754_out1;

  Logical_Operator_out851_out1 <= Logical_Operator_out723_out1 XOR Logical_Operator_out755_out1;

  Logical_Operator_out852_out1 <= Logical_Operator_out724_out1 XOR Logical_Operator_out756_out1;

  Logical_Operator_out853_out1 <= Logical_Operator_out725_out1 XOR Logical_Operator_out757_out1;

  Logical_Operator_out854_out1 <= Logical_Operator_out726_out1 XOR Logical_Operator_out758_out1;

  Logical_Operator_out855_out1 <= Logical_Operator_out727_out1 XOR Logical_Operator_out759_out1;

  Logical_Operator_out856_out1 <= Logical_Operator_out728_out1 XOR Logical_Operator_out760_out1;

  Logical_Operator_out857_out1 <= Logical_Operator_out729_out1 XOR Logical_Operator_out761_out1;

  Logical_Operator_out858_out1 <= Logical_Operator_out730_out1 XOR Logical_Operator_out762_out1;

  Logical_Operator_out859_out1 <= Logical_Operator_out731_out1 XOR Logical_Operator_out763_out1;

  Logical_Operator_out860_out1 <= Logical_Operator_out732_out1 XOR Logical_Operator_out764_out1;

  Logical_Operator_out861_out1 <= Logical_Operator_out733_out1 XOR Logical_Operator_out765_out1;

  Logical_Operator_out862_out1 <= Logical_Operator_out734_out1 XOR Logical_Operator_out766_out1;

  Logical_Operator_out863_out1 <= Logical_Operator_out735_out1 XOR Logical_Operator_out767_out1;

  Logical_Operator_out864_out1 <= Logical_Operator_out736_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out865_out1 <= Logical_Operator_out593_out1 XOR Logical_Operator_out625_out1;

  Logical_Operator_out866_out1 <= Logical_Operator_out594_out1 XOR Logical_Operator_out626_out1;

  Logical_Operator_out867_out1 <= Logical_Operator_out595_out1 XOR Logical_Operator_out627_out1;

  Logical_Operator_out868_out1 <= Logical_Operator_out596_out1 XOR Logical_Operator_out628_out1;

  Logical_Operator_out869_out1 <= Logical_Operator_out597_out1 XOR Logical_Operator_out629_out1;

  Logical_Operator_out870_out1 <= Logical_Operator_out598_out1 XOR Logical_Operator_out630_out1;

  Logical_Operator_out871_out1 <= Logical_Operator_out599_out1 XOR Logical_Operator_out631_out1;

  Logical_Operator_out872_out1 <= Logical_Operator_out600_out1 XOR Logical_Operator_out632_out1;

  Logical_Operator_out873_out1 <= Logical_Operator_out601_out1 XOR Logical_Operator_out633_out1;

  Logical_Operator_out874_out1 <= Logical_Operator_out602_out1 XOR Logical_Operator_out634_out1;

  Logical_Operator_out875_out1 <= Logical_Operator_out603_out1 XOR Logical_Operator_out635_out1;

  Logical_Operator_out876_out1 <= Logical_Operator_out604_out1 XOR Logical_Operator_out636_out1;

  Logical_Operator_out877_out1 <= Logical_Operator_out605_out1 XOR Logical_Operator_out637_out1;

  Logical_Operator_out878_out1 <= Logical_Operator_out606_out1 XOR Logical_Operator_out638_out1;

  Logical_Operator_out879_out1 <= Logical_Operator_out607_out1 XOR Logical_Operator_out639_out1;

  Logical_Operator_out880_out1 <= Logical_Operator_out608_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out881_out1 <= Logical_Operator_out473_out1 XOR Logical_Operator_out505_out1;

  Logical_Operator_out882_out1 <= Logical_Operator_out474_out1 XOR Logical_Operator_out506_out1;

  Logical_Operator_out883_out1 <= Logical_Operator_out475_out1 XOR Logical_Operator_out507_out1;

  Logical_Operator_out884_out1 <= Logical_Operator_out476_out1 XOR Logical_Operator_out508_out1;

  Logical_Operator_out885_out1 <= Logical_Operator_out477_out1 XOR Logical_Operator_out509_out1;

  Logical_Operator_out886_out1 <= Logical_Operator_out478_out1 XOR Logical_Operator_out510_out1;

  Logical_Operator_out887_out1 <= Logical_Operator_out479_out1 XOR Logical_Operator_out511_out1;

  Logical_Operator_out888_out1 <= Logical_Operator_out480_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out889_out1 <= Logical_Operator_out349_out1 XOR Logical_Operator_out381_out1;

  Logical_Operator_out890_out1 <= Logical_Operator_out350_out1 XOR Logical_Operator_out382_out1;

  Logical_Operator_out891_out1 <= Logical_Operator_out351_out1 XOR Logical_Operator_out383_out1;

  Logical_Operator_out892_out1 <= Logical_Operator_out352_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out893_out1 <= Logical_Operator_out223_out1 XOR Logical_Operator_out255_out1;

  Logical_Operator_out894_out1 <= Logical_Operator_out224_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out895_out1 <= Logical_Operator_out96_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out896_out1 <= in192 XOR in256;

  Logical_Operator_out897_out1 <= Logical_Operator_out769_out1 XOR Logical_Operator_out833_out1;

  Logical_Operator_out898_out1 <= Logical_Operator_out770_out1 XOR Logical_Operator_out834_out1;

  Logical_Operator_out899_out1 <= Logical_Operator_out771_out1 XOR Logical_Operator_out835_out1;

  Logical_Operator_out900_out1 <= Logical_Operator_out772_out1 XOR Logical_Operator_out836_out1;

  Logical_Operator_out901_out1 <= Logical_Operator_out773_out1 XOR Logical_Operator_out837_out1;

  Logical_Operator_out902_out1 <= Logical_Operator_out774_out1 XOR Logical_Operator_out838_out1;

  Logical_Operator_out903_out1 <= Logical_Operator_out775_out1 XOR Logical_Operator_out839_out1;

  Logical_Operator_out904_out1 <= Logical_Operator_out776_out1 XOR Logical_Operator_out840_out1;

  Logical_Operator_out905_out1 <= Logical_Operator_out777_out1 XOR Logical_Operator_out841_out1;

  Logical_Operator_out906_out1 <= Logical_Operator_out778_out1 XOR Logical_Operator_out842_out1;

  Logical_Operator_out907_out1 <= Logical_Operator_out779_out1 XOR Logical_Operator_out843_out1;

  Logical_Operator_out908_out1 <= Logical_Operator_out780_out1 XOR Logical_Operator_out844_out1;

  Logical_Operator_out909_out1 <= Logical_Operator_out781_out1 XOR Logical_Operator_out845_out1;

  Logical_Operator_out910_out1 <= Logical_Operator_out782_out1 XOR Logical_Operator_out846_out1;

  Logical_Operator_out911_out1 <= Logical_Operator_out783_out1 XOR Logical_Operator_out847_out1;

  Logical_Operator_out912_out1 <= Logical_Operator_out784_out1 XOR Logical_Operator_out848_out1;

  Logical_Operator_out913_out1 <= Logical_Operator_out785_out1 XOR Logical_Operator_out849_out1;

  Logical_Operator_out914_out1 <= Logical_Operator_out786_out1 XOR Logical_Operator_out850_out1;

  Logical_Operator_out915_out1 <= Logical_Operator_out787_out1 XOR Logical_Operator_out851_out1;

  Logical_Operator_out916_out1 <= Logical_Operator_out788_out1 XOR Logical_Operator_out852_out1;

  Logical_Operator_out917_out1 <= Logical_Operator_out789_out1 XOR Logical_Operator_out853_out1;

  Logical_Operator_out918_out1 <= Logical_Operator_out790_out1 XOR Logical_Operator_out854_out1;

  Logical_Operator_out919_out1 <= Logical_Operator_out791_out1 XOR Logical_Operator_out855_out1;

  Logical_Operator_out920_out1 <= Logical_Operator_out792_out1 XOR Logical_Operator_out856_out1;

  Logical_Operator_out921_out1 <= Logical_Operator_out793_out1 XOR Logical_Operator_out857_out1;

  Logical_Operator_out922_out1 <= Logical_Operator_out794_out1 XOR Logical_Operator_out858_out1;

  Logical_Operator_out923_out1 <= Logical_Operator_out795_out1 XOR Logical_Operator_out859_out1;

  Logical_Operator_out924_out1 <= Logical_Operator_out796_out1 XOR Logical_Operator_out860_out1;

  Logical_Operator_out925_out1 <= Logical_Operator_out797_out1 XOR Logical_Operator_out861_out1;

  Logical_Operator_out926_out1 <= Logical_Operator_out798_out1 XOR Logical_Operator_out862_out1;

  Logical_Operator_out927_out1 <= Logical_Operator_out799_out1 XOR Logical_Operator_out863_out1;

  Logical_Operator_out928_out1 <= Logical_Operator_out800_out1 XOR Logical_Operator_out864_out1;

  Logical_Operator_out929_out1 <= Logical_Operator_out801_out1 XOR Logical_Operator_out865_out1;

  Logical_Operator_out930_out1 <= Logical_Operator_out802_out1 XOR Logical_Operator_out866_out1;

  Logical_Operator_out931_out1 <= Logical_Operator_out803_out1 XOR Logical_Operator_out867_out1;

  Logical_Operator_out932_out1 <= Logical_Operator_out804_out1 XOR Logical_Operator_out868_out1;

  Logical_Operator_out933_out1 <= Logical_Operator_out805_out1 XOR Logical_Operator_out869_out1;

  Logical_Operator_out934_out1 <= Logical_Operator_out806_out1 XOR Logical_Operator_out870_out1;

  Logical_Operator_out935_out1 <= Logical_Operator_out807_out1 XOR Logical_Operator_out871_out1;

  Logical_Operator_out936_out1 <= Logical_Operator_out808_out1 XOR Logical_Operator_out872_out1;

  Logical_Operator_out937_out1 <= Logical_Operator_out809_out1 XOR Logical_Operator_out873_out1;

  Logical_Operator_out938_out1 <= Logical_Operator_out810_out1 XOR Logical_Operator_out874_out1;

  Logical_Operator_out939_out1 <= Logical_Operator_out811_out1 XOR Logical_Operator_out875_out1;

  Logical_Operator_out940_out1 <= Logical_Operator_out812_out1 XOR Logical_Operator_out876_out1;

  Logical_Operator_out941_out1 <= Logical_Operator_out813_out1 XOR Logical_Operator_out877_out1;

  Logical_Operator_out942_out1 <= Logical_Operator_out814_out1 XOR Logical_Operator_out878_out1;

  Logical_Operator_out943_out1 <= Logical_Operator_out815_out1 XOR Logical_Operator_out879_out1;

  Logical_Operator_out944_out1 <= Logical_Operator_out816_out1 XOR Logical_Operator_out880_out1;

  Logical_Operator_out945_out1 <= Logical_Operator_out817_out1 XOR Logical_Operator_out881_out1;

  Logical_Operator_out946_out1 <= Logical_Operator_out818_out1 XOR Logical_Operator_out882_out1;

  Logical_Operator_out947_out1 <= Logical_Operator_out819_out1 XOR Logical_Operator_out883_out1;

  Logical_Operator_out948_out1 <= Logical_Operator_out820_out1 XOR Logical_Operator_out884_out1;

  Logical_Operator_out949_out1 <= Logical_Operator_out821_out1 XOR Logical_Operator_out885_out1;

  Logical_Operator_out950_out1 <= Logical_Operator_out822_out1 XOR Logical_Operator_out886_out1;

  Logical_Operator_out951_out1 <= Logical_Operator_out823_out1 XOR Logical_Operator_out887_out1;

  Logical_Operator_out952_out1 <= Logical_Operator_out824_out1 XOR Logical_Operator_out888_out1;

  Logical_Operator_out953_out1 <= Logical_Operator_out825_out1 XOR Logical_Operator_out889_out1;

  Logical_Operator_out954_out1 <= Logical_Operator_out826_out1 XOR Logical_Operator_out890_out1;

  Logical_Operator_out955_out1 <= Logical_Operator_out827_out1 XOR Logical_Operator_out891_out1;

  Logical_Operator_out956_out1 <= Logical_Operator_out828_out1 XOR Logical_Operator_out892_out1;

  Logical_Operator_out957_out1 <= Logical_Operator_out829_out1 XOR Logical_Operator_out893_out1;

  Logical_Operator_out958_out1 <= Logical_Operator_out830_out1 XOR Logical_Operator_out894_out1;

  Logical_Operator_out959_out1 <= Logical_Operator_out831_out1 XOR Logical_Operator_out895_out1;

  Logical_Operator_out960_out1 <= Logical_Operator_out832_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out961_out1 <= Logical_Operator_out673_out1 XOR Logical_Operator_out737_out1;

  Logical_Operator_out962_out1 <= Logical_Operator_out674_out1 XOR Logical_Operator_out738_out1;

  Logical_Operator_out963_out1 <= Logical_Operator_out675_out1 XOR Logical_Operator_out739_out1;

  Logical_Operator_out964_out1 <= Logical_Operator_out676_out1 XOR Logical_Operator_out740_out1;

  Logical_Operator_out965_out1 <= Logical_Operator_out677_out1 XOR Logical_Operator_out741_out1;

  Logical_Operator_out966_out1 <= Logical_Operator_out678_out1 XOR Logical_Operator_out742_out1;

  Logical_Operator_out967_out1 <= Logical_Operator_out679_out1 XOR Logical_Operator_out743_out1;

  Logical_Operator_out968_out1 <= Logical_Operator_out680_out1 XOR Logical_Operator_out744_out1;

  Logical_Operator_out969_out1 <= Logical_Operator_out681_out1 XOR Logical_Operator_out745_out1;

  Logical_Operator_out970_out1 <= Logical_Operator_out682_out1 XOR Logical_Operator_out746_out1;

  Logical_Operator_out971_out1 <= Logical_Operator_out683_out1 XOR Logical_Operator_out747_out1;

  Logical_Operator_out972_out1 <= Logical_Operator_out684_out1 XOR Logical_Operator_out748_out1;

  Logical_Operator_out973_out1 <= Logical_Operator_out685_out1 XOR Logical_Operator_out749_out1;

  Logical_Operator_out974_out1 <= Logical_Operator_out686_out1 XOR Logical_Operator_out750_out1;

  Logical_Operator_out975_out1 <= Logical_Operator_out687_out1 XOR Logical_Operator_out751_out1;

  Logical_Operator_out976_out1 <= Logical_Operator_out688_out1 XOR Logical_Operator_out752_out1;

  Logical_Operator_out977_out1 <= Logical_Operator_out689_out1 XOR Logical_Operator_out753_out1;

  Logical_Operator_out978_out1 <= Logical_Operator_out690_out1 XOR Logical_Operator_out754_out1;

  Logical_Operator_out979_out1 <= Logical_Operator_out691_out1 XOR Logical_Operator_out755_out1;

  Logical_Operator_out980_out1 <= Logical_Operator_out692_out1 XOR Logical_Operator_out756_out1;

  Logical_Operator_out981_out1 <= Logical_Operator_out693_out1 XOR Logical_Operator_out757_out1;

  Logical_Operator_out982_out1 <= Logical_Operator_out694_out1 XOR Logical_Operator_out758_out1;

  Logical_Operator_out983_out1 <= Logical_Operator_out695_out1 XOR Logical_Operator_out759_out1;

  Logical_Operator_out984_out1 <= Logical_Operator_out696_out1 XOR Logical_Operator_out760_out1;

  Logical_Operator_out985_out1 <= Logical_Operator_out697_out1 XOR Logical_Operator_out761_out1;

  Logical_Operator_out986_out1 <= Logical_Operator_out698_out1 XOR Logical_Operator_out762_out1;

  Logical_Operator_out987_out1 <= Logical_Operator_out699_out1 XOR Logical_Operator_out763_out1;

  Logical_Operator_out988_out1 <= Logical_Operator_out700_out1 XOR Logical_Operator_out764_out1;

  Logical_Operator_out989_out1 <= Logical_Operator_out701_out1 XOR Logical_Operator_out765_out1;

  Logical_Operator_out990_out1 <= Logical_Operator_out702_out1 XOR Logical_Operator_out766_out1;

  Logical_Operator_out991_out1 <= Logical_Operator_out703_out1 XOR Logical_Operator_out767_out1;

  Logical_Operator_out992_out1 <= Logical_Operator_out704_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out993_out1 <= Logical_Operator_out561_out1 XOR Logical_Operator_out625_out1;

  Logical_Operator_out994_out1 <= Logical_Operator_out562_out1 XOR Logical_Operator_out626_out1;

  Logical_Operator_out995_out1 <= Logical_Operator_out563_out1 XOR Logical_Operator_out627_out1;

  Logical_Operator_out996_out1 <= Logical_Operator_out564_out1 XOR Logical_Operator_out628_out1;

  Logical_Operator_out997_out1 <= Logical_Operator_out565_out1 XOR Logical_Operator_out629_out1;

  Logical_Operator_out998_out1 <= Logical_Operator_out566_out1 XOR Logical_Operator_out630_out1;

  Logical_Operator_out999_out1 <= Logical_Operator_out567_out1 XOR Logical_Operator_out631_out1;

  Logical_Operator_out1000_out1 <= Logical_Operator_out568_out1 XOR Logical_Operator_out632_out1;

  Logical_Operator_out1001_out1 <= Logical_Operator_out569_out1 XOR Logical_Operator_out633_out1;

  Logical_Operator_out1002_out1 <= Logical_Operator_out570_out1 XOR Logical_Operator_out634_out1;

  Logical_Operator_out1003_out1 <= Logical_Operator_out571_out1 XOR Logical_Operator_out635_out1;

  Logical_Operator_out1004_out1 <= Logical_Operator_out572_out1 XOR Logical_Operator_out636_out1;

  Logical_Operator_out1005_out1 <= Logical_Operator_out573_out1 XOR Logical_Operator_out637_out1;

  Logical_Operator_out1006_out1 <= Logical_Operator_out574_out1 XOR Logical_Operator_out638_out1;

  Logical_Operator_out1007_out1 <= Logical_Operator_out575_out1 XOR Logical_Operator_out639_out1;

  Logical_Operator_out1008_out1 <= Logical_Operator_out576_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out1009_out1 <= Logical_Operator_out441_out1 XOR Logical_Operator_out505_out1;

  Logical_Operator_out1010_out1 <= Logical_Operator_out442_out1 XOR Logical_Operator_out506_out1;

  Logical_Operator_out1011_out1 <= Logical_Operator_out443_out1 XOR Logical_Operator_out507_out1;

  Logical_Operator_out1012_out1 <= Logical_Operator_out444_out1 XOR Logical_Operator_out508_out1;

  Logical_Operator_out1013_out1 <= Logical_Operator_out445_out1 XOR Logical_Operator_out509_out1;

  Logical_Operator_out1014_out1 <= Logical_Operator_out446_out1 XOR Logical_Operator_out510_out1;

  Logical_Operator_out1015_out1 <= Logical_Operator_out447_out1 XOR Logical_Operator_out511_out1;

  Logical_Operator_out1016_out1 <= Logical_Operator_out448_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out1017_out1 <= Logical_Operator_out317_out1 XOR Logical_Operator_out381_out1;

  Logical_Operator_out1018_out1 <= Logical_Operator_out318_out1 XOR Logical_Operator_out382_out1;

  Logical_Operator_out1019_out1 <= Logical_Operator_out319_out1 XOR Logical_Operator_out383_out1;

  Logical_Operator_out1020_out1 <= Logical_Operator_out320_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out1021_out1 <= Logical_Operator_out191_out1 XOR Logical_Operator_out255_out1;

  Logical_Operator_out1022_out1 <= Logical_Operator_out192_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out1023_out1 <= Logical_Operator_out64_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out1024_out1 <= in128 XOR in256;

  out1 <= Logical_Operator_out897_out1;

  out2 <= Logical_Operator_out898_out1;

  out3 <= Logical_Operator_out899_out1;

  out4 <= Logical_Operator_out900_out1;

  out5 <= Logical_Operator_out901_out1;

  out6 <= Logical_Operator_out902_out1;

  out7 <= Logical_Operator_out903_out1;

  out8 <= Logical_Operator_out904_out1;

  out9 <= Logical_Operator_out905_out1;

  out10 <= Logical_Operator_out906_out1;

  out11 <= Logical_Operator_out907_out1;

  out12 <= Logical_Operator_out908_out1;

  out13 <= Logical_Operator_out909_out1;

  out14 <= Logical_Operator_out910_out1;

  out15 <= Logical_Operator_out911_out1;

  out16 <= Logical_Operator_out912_out1;

  out17 <= Logical_Operator_out913_out1;

  out18 <= Logical_Operator_out914_out1;

  out19 <= Logical_Operator_out915_out1;

  out20 <= Logical_Operator_out916_out1;

  out21 <= Logical_Operator_out917_out1;

  out22 <= Logical_Operator_out918_out1;

  out23 <= Logical_Operator_out919_out1;

  out24 <= Logical_Operator_out920_out1;

  out25 <= Logical_Operator_out921_out1;

  out26 <= Logical_Operator_out922_out1;

  out27 <= Logical_Operator_out923_out1;

  out28 <= Logical_Operator_out924_out1;

  out29 <= Logical_Operator_out925_out1;

  out30 <= Logical_Operator_out926_out1;

  out31 <= Logical_Operator_out927_out1;

  out32 <= Logical_Operator_out928_out1;

  out33 <= Logical_Operator_out929_out1;

  out34 <= Logical_Operator_out930_out1;

  out35 <= Logical_Operator_out931_out1;

  out36 <= Logical_Operator_out932_out1;

  out37 <= Logical_Operator_out933_out1;

  out38 <= Logical_Operator_out934_out1;

  out39 <= Logical_Operator_out935_out1;

  out40 <= Logical_Operator_out936_out1;

  out41 <= Logical_Operator_out937_out1;

  out42 <= Logical_Operator_out938_out1;

  out43 <= Logical_Operator_out939_out1;

  out44 <= Logical_Operator_out940_out1;

  out45 <= Logical_Operator_out941_out1;

  out46 <= Logical_Operator_out942_out1;

  out47 <= Logical_Operator_out943_out1;

  out48 <= Logical_Operator_out944_out1;

  out49 <= Logical_Operator_out945_out1;

  out50 <= Logical_Operator_out946_out1;

  out51 <= Logical_Operator_out947_out1;

  out52 <= Logical_Operator_out948_out1;

  out53 <= Logical_Operator_out949_out1;

  out54 <= Logical_Operator_out950_out1;

  out55 <= Logical_Operator_out951_out1;

  out56 <= Logical_Operator_out952_out1;

  out57 <= Logical_Operator_out953_out1;

  out58 <= Logical_Operator_out954_out1;

  out59 <= Logical_Operator_out955_out1;

  out60 <= Logical_Operator_out956_out1;

  out61 <= Logical_Operator_out957_out1;

  out62 <= Logical_Operator_out958_out1;

  out63 <= Logical_Operator_out959_out1;

  out64 <= Logical_Operator_out960_out1;

  out65 <= Logical_Operator_out961_out1;

  out66 <= Logical_Operator_out962_out1;

  out67 <= Logical_Operator_out963_out1;

  out68 <= Logical_Operator_out964_out1;

  out69 <= Logical_Operator_out965_out1;

  out70 <= Logical_Operator_out966_out1;

  out71 <= Logical_Operator_out967_out1;

  out72 <= Logical_Operator_out968_out1;

  out73 <= Logical_Operator_out969_out1;

  out74 <= Logical_Operator_out970_out1;

  out75 <= Logical_Operator_out971_out1;

  out76 <= Logical_Operator_out972_out1;

  out77 <= Logical_Operator_out973_out1;

  out78 <= Logical_Operator_out974_out1;

  out79 <= Logical_Operator_out975_out1;

  out80 <= Logical_Operator_out976_out1;

  out81 <= Logical_Operator_out977_out1;

  out82 <= Logical_Operator_out978_out1;

  out83 <= Logical_Operator_out979_out1;

  out84 <= Logical_Operator_out980_out1;

  out85 <= Logical_Operator_out981_out1;

  out86 <= Logical_Operator_out982_out1;

  out87 <= Logical_Operator_out983_out1;

  out88 <= Logical_Operator_out984_out1;

  out89 <= Logical_Operator_out985_out1;

  out90 <= Logical_Operator_out986_out1;

  out91 <= Logical_Operator_out987_out1;

  out92 <= Logical_Operator_out988_out1;

  out93 <= Logical_Operator_out989_out1;

  out94 <= Logical_Operator_out990_out1;

  out95 <= Logical_Operator_out991_out1;

  out96 <= Logical_Operator_out992_out1;

  out97 <= Logical_Operator_out993_out1;

  out98 <= Logical_Operator_out994_out1;

  out99 <= Logical_Operator_out995_out1;

  out100 <= Logical_Operator_out996_out1;

  out101 <= Logical_Operator_out997_out1;

  out102 <= Logical_Operator_out998_out1;

  out103 <= Logical_Operator_out999_out1;

  out104 <= Logical_Operator_out1000_out1;

  out105 <= Logical_Operator_out1001_out1;

  out106 <= Logical_Operator_out1002_out1;

  out107 <= Logical_Operator_out1003_out1;

  out108 <= Logical_Operator_out1004_out1;

  out109 <= Logical_Operator_out1005_out1;

  out110 <= Logical_Operator_out1006_out1;

  out111 <= Logical_Operator_out1007_out1;

  out112 <= Logical_Operator_out1008_out1;

  out113 <= Logical_Operator_out1009_out1;

  out114 <= Logical_Operator_out1010_out1;

  out115 <= Logical_Operator_out1011_out1;

  out116 <= Logical_Operator_out1012_out1;

  out117 <= Logical_Operator_out1013_out1;

  out118 <= Logical_Operator_out1014_out1;

  out119 <= Logical_Operator_out1015_out1;

  out120 <= Logical_Operator_out1016_out1;

  out121 <= Logical_Operator_out1017_out1;

  out122 <= Logical_Operator_out1018_out1;

  out123 <= Logical_Operator_out1019_out1;

  out124 <= Logical_Operator_out1020_out1;

  out125 <= Logical_Operator_out1021_out1;

  out126 <= Logical_Operator_out1022_out1;

  out127 <= Logical_Operator_out1023_out1;

  out128 <= Logical_Operator_out1024_out1;

  out129 <= Logical_Operator_out833_out1;

  out130 <= Logical_Operator_out834_out1;

  out131 <= Logical_Operator_out835_out1;

  out132 <= Logical_Operator_out836_out1;

  out133 <= Logical_Operator_out837_out1;

  out134 <= Logical_Operator_out838_out1;

  out135 <= Logical_Operator_out839_out1;

  out136 <= Logical_Operator_out840_out1;

  out137 <= Logical_Operator_out841_out1;

  out138 <= Logical_Operator_out842_out1;

  out139 <= Logical_Operator_out843_out1;

  out140 <= Logical_Operator_out844_out1;

  out141 <= Logical_Operator_out845_out1;

  out142 <= Logical_Operator_out846_out1;

  out143 <= Logical_Operator_out847_out1;

  out144 <= Logical_Operator_out848_out1;

  out145 <= Logical_Operator_out849_out1;

  out146 <= Logical_Operator_out850_out1;

  out147 <= Logical_Operator_out851_out1;

  out148 <= Logical_Operator_out852_out1;

  out149 <= Logical_Operator_out853_out1;

  out150 <= Logical_Operator_out854_out1;

  out151 <= Logical_Operator_out855_out1;

  out152 <= Logical_Operator_out856_out1;

  out153 <= Logical_Operator_out857_out1;

  out154 <= Logical_Operator_out858_out1;

  out155 <= Logical_Operator_out859_out1;

  out156 <= Logical_Operator_out860_out1;

  out157 <= Logical_Operator_out861_out1;

  out158 <= Logical_Operator_out862_out1;

  out159 <= Logical_Operator_out863_out1;

  out160 <= Logical_Operator_out864_out1;

  out161 <= Logical_Operator_out865_out1;

  out162 <= Logical_Operator_out866_out1;

  out163 <= Logical_Operator_out867_out1;

  out164 <= Logical_Operator_out868_out1;

  out165 <= Logical_Operator_out869_out1;

  out166 <= Logical_Operator_out870_out1;

  out167 <= Logical_Operator_out871_out1;

  out168 <= Logical_Operator_out872_out1;

  out169 <= Logical_Operator_out873_out1;

  out170 <= Logical_Operator_out874_out1;

  out171 <= Logical_Operator_out875_out1;

  out172 <= Logical_Operator_out876_out1;

  out173 <= Logical_Operator_out877_out1;

  out174 <= Logical_Operator_out878_out1;

  out175 <= Logical_Operator_out879_out1;

  out176 <= Logical_Operator_out880_out1;

  out177 <= Logical_Operator_out881_out1;

  out178 <= Logical_Operator_out882_out1;

  out179 <= Logical_Operator_out883_out1;

  out180 <= Logical_Operator_out884_out1;

  out181 <= Logical_Operator_out885_out1;

  out182 <= Logical_Operator_out886_out1;

  out183 <= Logical_Operator_out887_out1;

  out184 <= Logical_Operator_out888_out1;

  out185 <= Logical_Operator_out889_out1;

  out186 <= Logical_Operator_out890_out1;

  out187 <= Logical_Operator_out891_out1;

  out188 <= Logical_Operator_out892_out1;

  out189 <= Logical_Operator_out893_out1;

  out190 <= Logical_Operator_out894_out1;

  out191 <= Logical_Operator_out895_out1;

  out192 <= Logical_Operator_out896_out1;

  out193 <= Logical_Operator_out737_out1;

  out194 <= Logical_Operator_out738_out1;

  out195 <= Logical_Operator_out739_out1;

  out196 <= Logical_Operator_out740_out1;

  out197 <= Logical_Operator_out741_out1;

  out198 <= Logical_Operator_out742_out1;

  out199 <= Logical_Operator_out743_out1;

  out200 <= Logical_Operator_out744_out1;

  out201 <= Logical_Operator_out745_out1;

  out202 <= Logical_Operator_out746_out1;

  out203 <= Logical_Operator_out747_out1;

  out204 <= Logical_Operator_out748_out1;

  out205 <= Logical_Operator_out749_out1;

  out206 <= Logical_Operator_out750_out1;

  out207 <= Logical_Operator_out751_out1;

  out208 <= Logical_Operator_out752_out1;

  out209 <= Logical_Operator_out753_out1;

  out210 <= Logical_Operator_out754_out1;

  out211 <= Logical_Operator_out755_out1;

  out212 <= Logical_Operator_out756_out1;

  out213 <= Logical_Operator_out757_out1;

  out214 <= Logical_Operator_out758_out1;

  out215 <= Logical_Operator_out759_out1;

  out216 <= Logical_Operator_out760_out1;

  out217 <= Logical_Operator_out761_out1;

  out218 <= Logical_Operator_out762_out1;

  out219 <= Logical_Operator_out763_out1;

  out220 <= Logical_Operator_out764_out1;

  out221 <= Logical_Operator_out765_out1;

  out222 <= Logical_Operator_out766_out1;

  out223 <= Logical_Operator_out767_out1;

  out224 <= Logical_Operator_out768_out1;

  out225 <= Logical_Operator_out625_out1;

  out226 <= Logical_Operator_out626_out1;

  out227 <= Logical_Operator_out627_out1;

  out228 <= Logical_Operator_out628_out1;

  out229 <= Logical_Operator_out629_out1;

  out230 <= Logical_Operator_out630_out1;

  out231 <= Logical_Operator_out631_out1;

  out232 <= Logical_Operator_out632_out1;

  out233 <= Logical_Operator_out633_out1;

  out234 <= Logical_Operator_out634_out1;

  out235 <= Logical_Operator_out635_out1;

  out236 <= Logical_Operator_out636_out1;

  out237 <= Logical_Operator_out637_out1;

  out238 <= Logical_Operator_out638_out1;

  out239 <= Logical_Operator_out639_out1;

  out240 <= Logical_Operator_out640_out1;

  out241 <= Logical_Operator_out505_out1;

  out242 <= Logical_Operator_out506_out1;

  out243 <= Logical_Operator_out507_out1;

  out244 <= Logical_Operator_out508_out1;

  out245 <= Logical_Operator_out509_out1;

  out246 <= Logical_Operator_out510_out1;

  out247 <= Logical_Operator_out511_out1;

  out248 <= Logical_Operator_out512_out1;

  out249 <= Logical_Operator_out381_out1;

  out250 <= Logical_Operator_out382_out1;

  out251 <= Logical_Operator_out383_out1;

  out252 <= Logical_Operator_out384_out1;

  out253 <= Logical_Operator_out255_out1;

  out254 <= Logical_Operator_out256_out1;

  out255 <= Logical_Operator_out128_out1;

  out256 <= in256;

END rtl;
