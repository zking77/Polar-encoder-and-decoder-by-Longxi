LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY encoderN64 IS
PORT( 
	in1                               :   IN    std_logic;
	in2                               :   IN    std_logic;
	in3                               :   IN    std_logic;
	in4                               :   IN    std_logic;
	in5                               :   IN    std_logic;
	in6                               :   IN    std_logic;
	in7                               :   IN    std_logic;
	in8                               :   IN    std_logic;
	in9                               :   IN    std_logic;
	in10                               :   IN    std_logic;
	in11                               :   IN    std_logic;
	in12                               :   IN    std_logic;
	in13                               :   IN    std_logic;
	in14                               :   IN    std_logic;
	in15                               :   IN    std_logic;
	in16                               :   IN    std_logic;
	in17                               :   IN    std_logic;
	in18                               :   IN    std_logic;
	in19                               :   IN    std_logic;
	in20                               :   IN    std_logic;
	in21                               :   IN    std_logic;
	in22                               :   IN    std_logic;
	in23                               :   IN    std_logic;
	in24                               :   IN    std_logic;
	in25                               :   IN    std_logic;
	in26                               :   IN    std_logic;
	in27                               :   IN    std_logic;
	in28                               :   IN    std_logic;
	in29                               :   IN    std_logic;
	in30                               :   IN    std_logic;
	in31                               :   IN    std_logic;
	in32                               :   IN    std_logic;
	in33                               :   IN    std_logic;
	in34                               :   IN    std_logic;
	in35                               :   IN    std_logic;
	in36                               :   IN    std_logic;
	in37                               :   IN    std_logic;
	in38                               :   IN    std_logic;
	in39                               :   IN    std_logic;
	in40                               :   IN    std_logic;
	in41                               :   IN    std_logic;
	in42                               :   IN    std_logic;
	in43                               :   IN    std_logic;
	in44                               :   IN    std_logic;
	in45                               :   IN    std_logic;
	in46                               :   IN    std_logic;
	in47                               :   IN    std_logic;
	in48                               :   IN    std_logic;
	in49                               :   IN    std_logic;
	in50                               :   IN    std_logic;
	in51                               :   IN    std_logic;
	in52                               :   IN    std_logic;
	in53                               :   IN    std_logic;
	in54                               :   IN    std_logic;
	in55                               :   IN    std_logic;
	in56                               :   IN    std_logic;
	in57                               :   IN    std_logic;
	in58                               :   IN    std_logic;
	in59                               :   IN    std_logic;
	in60                               :   IN    std_logic;
	in61                               :   IN    std_logic;
	in62                               :   IN    std_logic;
	in63                               :   IN    std_logic;
	in64                               :   IN    std_logic;
	out1                               :   OUT    std_logic;
	out2                               :   OUT    std_logic;
	out3                               :   OUT    std_logic;
	out4                               :   OUT    std_logic;
	out5                               :   OUT    std_logic;
	out6                               :   OUT    std_logic;
	out7                               :   OUT    std_logic;
	out8                               :   OUT    std_logic;
	out9                               :   OUT    std_logic;
	out10                               :   OUT    std_logic;
	out11                               :   OUT    std_logic;
	out12                               :   OUT    std_logic;
	out13                               :   OUT    std_logic;
	out14                               :   OUT    std_logic;
	out15                               :   OUT    std_logic;
	out16                               :   OUT    std_logic;
	out17                               :   OUT    std_logic;
	out18                               :   OUT    std_logic;
	out19                               :   OUT    std_logic;
	out20                               :   OUT    std_logic;
	out21                               :   OUT    std_logic;
	out22                               :   OUT    std_logic;
	out23                               :   OUT    std_logic;
	out24                               :   OUT    std_logic;
	out25                               :   OUT    std_logic;
	out26                               :   OUT    std_logic;
	out27                               :   OUT    std_logic;
	out28                               :   OUT    std_logic;
	out29                               :   OUT    std_logic;
	out30                               :   OUT    std_logic;
	out31                               :   OUT    std_logic;
	out32                               :   OUT    std_logic;
	out33                               :   OUT    std_logic;
	out34                               :   OUT    std_logic;
	out35                               :   OUT    std_logic;
	out36                               :   OUT    std_logic;
	out37                               :   OUT    std_logic;
	out38                               :   OUT    std_logic;
	out39                               :   OUT    std_logic;
	out40                               :   OUT    std_logic;
	out41                               :   OUT    std_logic;
	out42                               :   OUT    std_logic;
	out43                               :   OUT    std_logic;
	out44                               :   OUT    std_logic;
	out45                               :   OUT    std_logic;
	out46                               :   OUT    std_logic;
	out47                               :   OUT    std_logic;
	out48                               :   OUT    std_logic;
	out49                               :   OUT    std_logic;
	out50                               :   OUT    std_logic;
	out51                               :   OUT    std_logic;
	out52                               :   OUT    std_logic;
	out53                               :   OUT    std_logic;
	out54                               :   OUT    std_logic;
	out55                               :   OUT    std_logic;
	out56                               :   OUT    std_logic;
	out57                               :   OUT    std_logic;
	out58                               :   OUT    std_logic;
	out59                               :   OUT    std_logic;
	out60                               :   OUT    std_logic;
	out61                               :   OUT    std_logic;
	out62                               :   OUT    std_logic;
	out63                               :   OUT    std_logic;
	out64                               :   OUT    std_logic
	);
END encoderN64;

ARCHITECTURE rtl OF encoderN64 IS

  SIGNAL Logical_Operator_out1_out1            : std_logic;
  SIGNAL Logical_Operator_out2_out1            : std_logic;
  SIGNAL Logical_Operator_out3_out1            : std_logic;
  SIGNAL Logical_Operator_out4_out1            : std_logic;
  SIGNAL Logical_Operator_out5_out1            : std_logic;
  SIGNAL Logical_Operator_out6_out1            : std_logic;
  SIGNAL Logical_Operator_out7_out1            : std_logic;
  SIGNAL Logical_Operator_out8_out1            : std_logic;
  SIGNAL Logical_Operator_out9_out1            : std_logic;
  SIGNAL Logical_Operator_out10_out1            : std_logic;
  SIGNAL Logical_Operator_out11_out1            : std_logic;
  SIGNAL Logical_Operator_out12_out1            : std_logic;
  SIGNAL Logical_Operator_out13_out1            : std_logic;
  SIGNAL Logical_Operator_out14_out1            : std_logic;
  SIGNAL Logical_Operator_out15_out1            : std_logic;
  SIGNAL Logical_Operator_out16_out1            : std_logic;
  SIGNAL Logical_Operator_out17_out1            : std_logic;
  SIGNAL Logical_Operator_out18_out1            : std_logic;
  SIGNAL Logical_Operator_out19_out1            : std_logic;
  SIGNAL Logical_Operator_out20_out1            : std_logic;
  SIGNAL Logical_Operator_out21_out1            : std_logic;
  SIGNAL Logical_Operator_out22_out1            : std_logic;
  SIGNAL Logical_Operator_out23_out1            : std_logic;
  SIGNAL Logical_Operator_out24_out1            : std_logic;
  SIGNAL Logical_Operator_out25_out1            : std_logic;
  SIGNAL Logical_Operator_out26_out1            : std_logic;
  SIGNAL Logical_Operator_out27_out1            : std_logic;
  SIGNAL Logical_Operator_out28_out1            : std_logic;
  SIGNAL Logical_Operator_out29_out1            : std_logic;
  SIGNAL Logical_Operator_out30_out1            : std_logic;
  SIGNAL Logical_Operator_out31_out1            : std_logic;
  SIGNAL Logical_Operator_out32_out1            : std_logic;
  SIGNAL Logical_Operator_out33_out1            : std_logic;
  SIGNAL Logical_Operator_out34_out1            : std_logic;
  SIGNAL Logical_Operator_out35_out1            : std_logic;
  SIGNAL Logical_Operator_out36_out1            : std_logic;
  SIGNAL Logical_Operator_out37_out1            : std_logic;
  SIGNAL Logical_Operator_out38_out1            : std_logic;
  SIGNAL Logical_Operator_out39_out1            : std_logic;
  SIGNAL Logical_Operator_out40_out1            : std_logic;
  SIGNAL Logical_Operator_out41_out1            : std_logic;
  SIGNAL Logical_Operator_out42_out1            : std_logic;
  SIGNAL Logical_Operator_out43_out1            : std_logic;
  SIGNAL Logical_Operator_out44_out1            : std_logic;
  SIGNAL Logical_Operator_out45_out1            : std_logic;
  SIGNAL Logical_Operator_out46_out1            : std_logic;
  SIGNAL Logical_Operator_out47_out1            : std_logic;
  SIGNAL Logical_Operator_out48_out1            : std_logic;
  SIGNAL Logical_Operator_out49_out1            : std_logic;
  SIGNAL Logical_Operator_out50_out1            : std_logic;
  SIGNAL Logical_Operator_out51_out1            : std_logic;
  SIGNAL Logical_Operator_out52_out1            : std_logic;
  SIGNAL Logical_Operator_out53_out1            : std_logic;
  SIGNAL Logical_Operator_out54_out1            : std_logic;
  SIGNAL Logical_Operator_out55_out1            : std_logic;
  SIGNAL Logical_Operator_out56_out1            : std_logic;
  SIGNAL Logical_Operator_out57_out1            : std_logic;
  SIGNAL Logical_Operator_out58_out1            : std_logic;
  SIGNAL Logical_Operator_out59_out1            : std_logic;
  SIGNAL Logical_Operator_out60_out1            : std_logic;
  SIGNAL Logical_Operator_out61_out1            : std_logic;
  SIGNAL Logical_Operator_out62_out1            : std_logic;
  SIGNAL Logical_Operator_out63_out1            : std_logic;
  SIGNAL Logical_Operator_out64_out1            : std_logic;
  SIGNAL Logical_Operator_out65_out1            : std_logic;
  SIGNAL Logical_Operator_out66_out1            : std_logic;
  SIGNAL Logical_Operator_out67_out1            : std_logic;
  SIGNAL Logical_Operator_out68_out1            : std_logic;
  SIGNAL Logical_Operator_out69_out1            : std_logic;
  SIGNAL Logical_Operator_out70_out1            : std_logic;
  SIGNAL Logical_Operator_out71_out1            : std_logic;
  SIGNAL Logical_Operator_out72_out1            : std_logic;
  SIGNAL Logical_Operator_out73_out1            : std_logic;
  SIGNAL Logical_Operator_out74_out1            : std_logic;
  SIGNAL Logical_Operator_out75_out1            : std_logic;
  SIGNAL Logical_Operator_out76_out1            : std_logic;
  SIGNAL Logical_Operator_out77_out1            : std_logic;
  SIGNAL Logical_Operator_out78_out1            : std_logic;
  SIGNAL Logical_Operator_out79_out1            : std_logic;
  SIGNAL Logical_Operator_out80_out1            : std_logic;
  SIGNAL Logical_Operator_out81_out1            : std_logic;
  SIGNAL Logical_Operator_out82_out1            : std_logic;
  SIGNAL Logical_Operator_out83_out1            : std_logic;
  SIGNAL Logical_Operator_out84_out1            : std_logic;
  SIGNAL Logical_Operator_out85_out1            : std_logic;
  SIGNAL Logical_Operator_out86_out1            : std_logic;
  SIGNAL Logical_Operator_out87_out1            : std_logic;
  SIGNAL Logical_Operator_out88_out1            : std_logic;
  SIGNAL Logical_Operator_out89_out1            : std_logic;
  SIGNAL Logical_Operator_out90_out1            : std_logic;
  SIGNAL Logical_Operator_out91_out1            : std_logic;
  SIGNAL Logical_Operator_out92_out1            : std_logic;
  SIGNAL Logical_Operator_out93_out1            : std_logic;
  SIGNAL Logical_Operator_out94_out1            : std_logic;
  SIGNAL Logical_Operator_out95_out1            : std_logic;
  SIGNAL Logical_Operator_out96_out1            : std_logic;
  SIGNAL Logical_Operator_out97_out1            : std_logic;
  SIGNAL Logical_Operator_out98_out1            : std_logic;
  SIGNAL Logical_Operator_out99_out1            : std_logic;
  SIGNAL Logical_Operator_out100_out1            : std_logic;
  SIGNAL Logical_Operator_out101_out1            : std_logic;
  SIGNAL Logical_Operator_out102_out1            : std_logic;
  SIGNAL Logical_Operator_out103_out1            : std_logic;
  SIGNAL Logical_Operator_out104_out1            : std_logic;
  SIGNAL Logical_Operator_out105_out1            : std_logic;
  SIGNAL Logical_Operator_out106_out1            : std_logic;
  SIGNAL Logical_Operator_out107_out1            : std_logic;
  SIGNAL Logical_Operator_out108_out1            : std_logic;
  SIGNAL Logical_Operator_out109_out1            : std_logic;
  SIGNAL Logical_Operator_out110_out1            : std_logic;
  SIGNAL Logical_Operator_out111_out1            : std_logic;
  SIGNAL Logical_Operator_out112_out1            : std_logic;
  SIGNAL Logical_Operator_out113_out1            : std_logic;
  SIGNAL Logical_Operator_out114_out1            : std_logic;
  SIGNAL Logical_Operator_out115_out1            : std_logic;
  SIGNAL Logical_Operator_out116_out1            : std_logic;
  SIGNAL Logical_Operator_out117_out1            : std_logic;
  SIGNAL Logical_Operator_out118_out1            : std_logic;
  SIGNAL Logical_Operator_out119_out1            : std_logic;
  SIGNAL Logical_Operator_out120_out1            : std_logic;
  SIGNAL Logical_Operator_out121_out1            : std_logic;
  SIGNAL Logical_Operator_out122_out1            : std_logic;
  SIGNAL Logical_Operator_out123_out1            : std_logic;
  SIGNAL Logical_Operator_out124_out1            : std_logic;
  SIGNAL Logical_Operator_out125_out1            : std_logic;
  SIGNAL Logical_Operator_out126_out1            : std_logic;
  SIGNAL Logical_Operator_out127_out1            : std_logic;
  SIGNAL Logical_Operator_out128_out1            : std_logic;
  SIGNAL Logical_Operator_out129_out1            : std_logic;
  SIGNAL Logical_Operator_out130_out1            : std_logic;
  SIGNAL Logical_Operator_out131_out1            : std_logic;
  SIGNAL Logical_Operator_out132_out1            : std_logic;
  SIGNAL Logical_Operator_out133_out1            : std_logic;
  SIGNAL Logical_Operator_out134_out1            : std_logic;
  SIGNAL Logical_Operator_out135_out1            : std_logic;
  SIGNAL Logical_Operator_out136_out1            : std_logic;
  SIGNAL Logical_Operator_out137_out1            : std_logic;
  SIGNAL Logical_Operator_out138_out1            : std_logic;
  SIGNAL Logical_Operator_out139_out1            : std_logic;
  SIGNAL Logical_Operator_out140_out1            : std_logic;
  SIGNAL Logical_Operator_out141_out1            : std_logic;
  SIGNAL Logical_Operator_out142_out1            : std_logic;
  SIGNAL Logical_Operator_out143_out1            : std_logic;
  SIGNAL Logical_Operator_out144_out1            : std_logic;
  SIGNAL Logical_Operator_out145_out1            : std_logic;
  SIGNAL Logical_Operator_out146_out1            : std_logic;
  SIGNAL Logical_Operator_out147_out1            : std_logic;
  SIGNAL Logical_Operator_out148_out1            : std_logic;
  SIGNAL Logical_Operator_out149_out1            : std_logic;
  SIGNAL Logical_Operator_out150_out1            : std_logic;
  SIGNAL Logical_Operator_out151_out1            : std_logic;
  SIGNAL Logical_Operator_out152_out1            : std_logic;
  SIGNAL Logical_Operator_out153_out1            : std_logic;
  SIGNAL Logical_Operator_out154_out1            : std_logic;
  SIGNAL Logical_Operator_out155_out1            : std_logic;
  SIGNAL Logical_Operator_out156_out1            : std_logic;
  SIGNAL Logical_Operator_out157_out1            : std_logic;
  SIGNAL Logical_Operator_out158_out1            : std_logic;
  SIGNAL Logical_Operator_out159_out1            : std_logic;
  SIGNAL Logical_Operator_out160_out1            : std_logic;
  SIGNAL Logical_Operator_out161_out1            : std_logic;
  SIGNAL Logical_Operator_out162_out1            : std_logic;
  SIGNAL Logical_Operator_out163_out1            : std_logic;
  SIGNAL Logical_Operator_out164_out1            : std_logic;
  SIGNAL Logical_Operator_out165_out1            : std_logic;
  SIGNAL Logical_Operator_out166_out1            : std_logic;
  SIGNAL Logical_Operator_out167_out1            : std_logic;
  SIGNAL Logical_Operator_out168_out1            : std_logic;
  SIGNAL Logical_Operator_out169_out1            : std_logic;
  SIGNAL Logical_Operator_out170_out1            : std_logic;
  SIGNAL Logical_Operator_out171_out1            : std_logic;
  SIGNAL Logical_Operator_out172_out1            : std_logic;
  SIGNAL Logical_Operator_out173_out1            : std_logic;
  SIGNAL Logical_Operator_out174_out1            : std_logic;
  SIGNAL Logical_Operator_out175_out1            : std_logic;
  SIGNAL Logical_Operator_out176_out1            : std_logic;
  SIGNAL Logical_Operator_out177_out1            : std_logic;
  SIGNAL Logical_Operator_out178_out1            : std_logic;
  SIGNAL Logical_Operator_out179_out1            : std_logic;
  SIGNAL Logical_Operator_out180_out1            : std_logic;
  SIGNAL Logical_Operator_out181_out1            : std_logic;
  SIGNAL Logical_Operator_out182_out1            : std_logic;
  SIGNAL Logical_Operator_out183_out1            : std_logic;
  SIGNAL Logical_Operator_out184_out1            : std_logic;
  SIGNAL Logical_Operator_out185_out1            : std_logic;
  SIGNAL Logical_Operator_out186_out1            : std_logic;
  SIGNAL Logical_Operator_out187_out1            : std_logic;
  SIGNAL Logical_Operator_out188_out1            : std_logic;
  SIGNAL Logical_Operator_out189_out1            : std_logic;
  SIGNAL Logical_Operator_out190_out1            : std_logic;
  SIGNAL Logical_Operator_out191_out1            : std_logic;
  SIGNAL Logical_Operator_out192_out1            : std_logic;

BEGIN

  Logical_Operator_out1_out1 <= in1 XOR in2;

  Logical_Operator_out2_out1 <= in3 XOR in4;

  Logical_Operator_out3_out1 <= in5 XOR in6;

  Logical_Operator_out4_out1 <= in7 XOR in8;

  Logical_Operator_out5_out1 <= in9 XOR in10;

  Logical_Operator_out6_out1 <= in11 XOR in12;

  Logical_Operator_out7_out1 <= in13 XOR in14;

  Logical_Operator_out8_out1 <= in15 XOR in16;

  Logical_Operator_out9_out1 <= in17 XOR in18;

  Logical_Operator_out10_out1 <= in19 XOR in20;

  Logical_Operator_out11_out1 <= in21 XOR in22;

  Logical_Operator_out12_out1 <= in23 XOR in24;

  Logical_Operator_out13_out1 <= in25 XOR in26;

  Logical_Operator_out14_out1 <= in27 XOR in28;

  Logical_Operator_out15_out1 <= in29 XOR in30;

  Logical_Operator_out16_out1 <= in31 XOR in32;

  Logical_Operator_out17_out1 <= in33 XOR in34;

  Logical_Operator_out18_out1 <= in35 XOR in36;

  Logical_Operator_out19_out1 <= in37 XOR in38;

  Logical_Operator_out20_out1 <= in39 XOR in40;

  Logical_Operator_out21_out1 <= in41 XOR in42;

  Logical_Operator_out22_out1 <= in43 XOR in44;

  Logical_Operator_out23_out1 <= in45 XOR in46;

  Logical_Operator_out24_out1 <= in47 XOR in48;

  Logical_Operator_out25_out1 <= in49 XOR in50;

  Logical_Operator_out26_out1 <= in51 XOR in52;

  Logical_Operator_out27_out1 <= in53 XOR in54;

  Logical_Operator_out28_out1 <= in55 XOR in56;

  Logical_Operator_out29_out1 <= in57 XOR in58;

  Logical_Operator_out30_out1 <= in59 XOR in60;

  Logical_Operator_out31_out1 <= in61 XOR in62;

  Logical_Operator_out32_out1 <= in63 XOR in64;

  Logical_Operator_out33_out1 <= Logical_Operator_out1_out1 XOR Logical_Operator_out2_out1;

  Logical_Operator_out34_out1 <= in2 XOR in4;

  Logical_Operator_out35_out1 <= Logical_Operator_out3_out1 XOR Logical_Operator_out4_out1;

  Logical_Operator_out36_out1 <= in6 XOR in8;

  Logical_Operator_out37_out1 <= Logical_Operator_out5_out1 XOR Logical_Operator_out6_out1;

  Logical_Operator_out38_out1 <= in10 XOR in12;

  Logical_Operator_out39_out1 <= Logical_Operator_out7_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out40_out1 <= in14 XOR in16;

  Logical_Operator_out41_out1 <= Logical_Operator_out9_out1 XOR Logical_Operator_out10_out1;

  Logical_Operator_out42_out1 <= in18 XOR in20;

  Logical_Operator_out43_out1 <= Logical_Operator_out11_out1 XOR Logical_Operator_out12_out1;

  Logical_Operator_out44_out1 <= in22 XOR in24;

  Logical_Operator_out45_out1 <= Logical_Operator_out13_out1 XOR Logical_Operator_out14_out1;

  Logical_Operator_out46_out1 <= in26 XOR in28;

  Logical_Operator_out47_out1 <= Logical_Operator_out15_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out48_out1 <= in30 XOR in32;

  Logical_Operator_out49_out1 <= Logical_Operator_out17_out1 XOR Logical_Operator_out18_out1;

  Logical_Operator_out50_out1 <= in34 XOR in36;

  Logical_Operator_out51_out1 <= Logical_Operator_out19_out1 XOR Logical_Operator_out20_out1;

  Logical_Operator_out52_out1 <= in38 XOR in40;

  Logical_Operator_out53_out1 <= Logical_Operator_out21_out1 XOR Logical_Operator_out22_out1;

  Logical_Operator_out54_out1 <= in42 XOR in44;

  Logical_Operator_out55_out1 <= Logical_Operator_out23_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out56_out1 <= in46 XOR in48;

  Logical_Operator_out57_out1 <= Logical_Operator_out25_out1 XOR Logical_Operator_out26_out1;

  Logical_Operator_out58_out1 <= in50 XOR in52;

  Logical_Operator_out59_out1 <= Logical_Operator_out27_out1 XOR Logical_Operator_out28_out1;

  Logical_Operator_out60_out1 <= in54 XOR in56;

  Logical_Operator_out61_out1 <= Logical_Operator_out29_out1 XOR Logical_Operator_out30_out1;

  Logical_Operator_out62_out1 <= in58 XOR in60;

  Logical_Operator_out63_out1 <= Logical_Operator_out31_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out64_out1 <= in62 XOR in64;

  Logical_Operator_out65_out1 <= Logical_Operator_out33_out1 XOR Logical_Operator_out35_out1;

  Logical_Operator_out66_out1 <= Logical_Operator_out34_out1 XOR Logical_Operator_out36_out1;

  Logical_Operator_out67_out1 <= Logical_Operator_out2_out1 XOR Logical_Operator_out4_out1;

  Logical_Operator_out68_out1 <= in4 XOR in8;

  Logical_Operator_out69_out1 <= Logical_Operator_out37_out1 XOR Logical_Operator_out39_out1;

  Logical_Operator_out70_out1 <= Logical_Operator_out38_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out71_out1 <= Logical_Operator_out6_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out72_out1 <= in12 XOR in16;

  Logical_Operator_out73_out1 <= Logical_Operator_out41_out1 XOR Logical_Operator_out43_out1;

  Logical_Operator_out74_out1 <= Logical_Operator_out42_out1 XOR Logical_Operator_out44_out1;

  Logical_Operator_out75_out1 <= Logical_Operator_out10_out1 XOR Logical_Operator_out12_out1;

  Logical_Operator_out76_out1 <= in20 XOR in24;

  Logical_Operator_out77_out1 <= Logical_Operator_out45_out1 XOR Logical_Operator_out47_out1;

  Logical_Operator_out78_out1 <= Logical_Operator_out46_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out79_out1 <= Logical_Operator_out14_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out80_out1 <= in28 XOR in32;

  Logical_Operator_out81_out1 <= Logical_Operator_out49_out1 XOR Logical_Operator_out51_out1;

  Logical_Operator_out82_out1 <= Logical_Operator_out50_out1 XOR Logical_Operator_out52_out1;

  Logical_Operator_out83_out1 <= Logical_Operator_out18_out1 XOR Logical_Operator_out20_out1;

  Logical_Operator_out84_out1 <= in36 XOR in40;

  Logical_Operator_out85_out1 <= Logical_Operator_out53_out1 XOR Logical_Operator_out55_out1;

  Logical_Operator_out86_out1 <= Logical_Operator_out54_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out87_out1 <= Logical_Operator_out22_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out88_out1 <= in44 XOR in48;

  Logical_Operator_out89_out1 <= Logical_Operator_out57_out1 XOR Logical_Operator_out59_out1;

  Logical_Operator_out90_out1 <= Logical_Operator_out58_out1 XOR Logical_Operator_out60_out1;

  Logical_Operator_out91_out1 <= Logical_Operator_out26_out1 XOR Logical_Operator_out28_out1;

  Logical_Operator_out92_out1 <= in52 XOR in56;

  Logical_Operator_out93_out1 <= Logical_Operator_out61_out1 XOR Logical_Operator_out63_out1;

  Logical_Operator_out94_out1 <= Logical_Operator_out62_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out95_out1 <= Logical_Operator_out30_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out96_out1 <= in60 XOR in64;

  Logical_Operator_out97_out1 <= Logical_Operator_out65_out1 XOR Logical_Operator_out69_out1;

  Logical_Operator_out98_out1 <= Logical_Operator_out66_out1 XOR Logical_Operator_out70_out1;

  Logical_Operator_out99_out1 <= Logical_Operator_out67_out1 XOR Logical_Operator_out71_out1;

  Logical_Operator_out100_out1 <= Logical_Operator_out68_out1 XOR Logical_Operator_out72_out1;

  Logical_Operator_out101_out1 <= Logical_Operator_out35_out1 XOR Logical_Operator_out39_out1;

  Logical_Operator_out102_out1 <= Logical_Operator_out36_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out103_out1 <= Logical_Operator_out4_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out104_out1 <= in8 XOR in16;

  Logical_Operator_out105_out1 <= Logical_Operator_out73_out1 XOR Logical_Operator_out77_out1;

  Logical_Operator_out106_out1 <= Logical_Operator_out74_out1 XOR Logical_Operator_out78_out1;

  Logical_Operator_out107_out1 <= Logical_Operator_out75_out1 XOR Logical_Operator_out79_out1;

  Logical_Operator_out108_out1 <= Logical_Operator_out76_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out109_out1 <= Logical_Operator_out43_out1 XOR Logical_Operator_out47_out1;

  Logical_Operator_out110_out1 <= Logical_Operator_out44_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out111_out1 <= Logical_Operator_out12_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out112_out1 <= in24 XOR in32;

  Logical_Operator_out113_out1 <= Logical_Operator_out81_out1 XOR Logical_Operator_out85_out1;

  Logical_Operator_out114_out1 <= Logical_Operator_out82_out1 XOR Logical_Operator_out86_out1;

  Logical_Operator_out115_out1 <= Logical_Operator_out83_out1 XOR Logical_Operator_out87_out1;

  Logical_Operator_out116_out1 <= Logical_Operator_out84_out1 XOR Logical_Operator_out88_out1;

  Logical_Operator_out117_out1 <= Logical_Operator_out51_out1 XOR Logical_Operator_out55_out1;

  Logical_Operator_out118_out1 <= Logical_Operator_out52_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out119_out1 <= Logical_Operator_out20_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out120_out1 <= in40 XOR in48;

  Logical_Operator_out121_out1 <= Logical_Operator_out89_out1 XOR Logical_Operator_out93_out1;

  Logical_Operator_out122_out1 <= Logical_Operator_out90_out1 XOR Logical_Operator_out94_out1;

  Logical_Operator_out123_out1 <= Logical_Operator_out91_out1 XOR Logical_Operator_out95_out1;

  Logical_Operator_out124_out1 <= Logical_Operator_out92_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out125_out1 <= Logical_Operator_out59_out1 XOR Logical_Operator_out63_out1;

  Logical_Operator_out126_out1 <= Logical_Operator_out60_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out127_out1 <= Logical_Operator_out28_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out128_out1 <= in56 XOR in64;

  Logical_Operator_out129_out1 <= Logical_Operator_out97_out1 XOR Logical_Operator_out105_out1;

  Logical_Operator_out130_out1 <= Logical_Operator_out98_out1 XOR Logical_Operator_out106_out1;

  Logical_Operator_out131_out1 <= Logical_Operator_out99_out1 XOR Logical_Operator_out107_out1;

  Logical_Operator_out132_out1 <= Logical_Operator_out100_out1 XOR Logical_Operator_out108_out1;

  Logical_Operator_out133_out1 <= Logical_Operator_out101_out1 XOR Logical_Operator_out109_out1;

  Logical_Operator_out134_out1 <= Logical_Operator_out102_out1 XOR Logical_Operator_out110_out1;

  Logical_Operator_out135_out1 <= Logical_Operator_out103_out1 XOR Logical_Operator_out111_out1;

  Logical_Operator_out136_out1 <= Logical_Operator_out104_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out137_out1 <= Logical_Operator_out69_out1 XOR Logical_Operator_out77_out1;

  Logical_Operator_out138_out1 <= Logical_Operator_out70_out1 XOR Logical_Operator_out78_out1;

  Logical_Operator_out139_out1 <= Logical_Operator_out71_out1 XOR Logical_Operator_out79_out1;

  Logical_Operator_out140_out1 <= Logical_Operator_out72_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out141_out1 <= Logical_Operator_out39_out1 XOR Logical_Operator_out47_out1;

  Logical_Operator_out142_out1 <= Logical_Operator_out40_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out143_out1 <= Logical_Operator_out8_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out144_out1 <= in16 XOR in32;

  Logical_Operator_out145_out1 <= Logical_Operator_out113_out1 XOR Logical_Operator_out121_out1;

  Logical_Operator_out146_out1 <= Logical_Operator_out114_out1 XOR Logical_Operator_out122_out1;

  Logical_Operator_out147_out1 <= Logical_Operator_out115_out1 XOR Logical_Operator_out123_out1;

  Logical_Operator_out148_out1 <= Logical_Operator_out116_out1 XOR Logical_Operator_out124_out1;

  Logical_Operator_out149_out1 <= Logical_Operator_out117_out1 XOR Logical_Operator_out125_out1;

  Logical_Operator_out150_out1 <= Logical_Operator_out118_out1 XOR Logical_Operator_out126_out1;

  Logical_Operator_out151_out1 <= Logical_Operator_out119_out1 XOR Logical_Operator_out127_out1;

  Logical_Operator_out152_out1 <= Logical_Operator_out120_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out153_out1 <= Logical_Operator_out85_out1 XOR Logical_Operator_out93_out1;

  Logical_Operator_out154_out1 <= Logical_Operator_out86_out1 XOR Logical_Operator_out94_out1;

  Logical_Operator_out155_out1 <= Logical_Operator_out87_out1 XOR Logical_Operator_out95_out1;

  Logical_Operator_out156_out1 <= Logical_Operator_out88_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out157_out1 <= Logical_Operator_out55_out1 XOR Logical_Operator_out63_out1;

  Logical_Operator_out158_out1 <= Logical_Operator_out56_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out159_out1 <= Logical_Operator_out24_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out160_out1 <= in48 XOR in64;

  Logical_Operator_out161_out1 <= Logical_Operator_out129_out1 XOR Logical_Operator_out145_out1;

  Logical_Operator_out162_out1 <= Logical_Operator_out130_out1 XOR Logical_Operator_out146_out1;

  Logical_Operator_out163_out1 <= Logical_Operator_out131_out1 XOR Logical_Operator_out147_out1;

  Logical_Operator_out164_out1 <= Logical_Operator_out132_out1 XOR Logical_Operator_out148_out1;

  Logical_Operator_out165_out1 <= Logical_Operator_out133_out1 XOR Logical_Operator_out149_out1;

  Logical_Operator_out166_out1 <= Logical_Operator_out134_out1 XOR Logical_Operator_out150_out1;

  Logical_Operator_out167_out1 <= Logical_Operator_out135_out1 XOR Logical_Operator_out151_out1;

  Logical_Operator_out168_out1 <= Logical_Operator_out136_out1 XOR Logical_Operator_out152_out1;

  Logical_Operator_out169_out1 <= Logical_Operator_out137_out1 XOR Logical_Operator_out153_out1;

  Logical_Operator_out170_out1 <= Logical_Operator_out138_out1 XOR Logical_Operator_out154_out1;

  Logical_Operator_out171_out1 <= Logical_Operator_out139_out1 XOR Logical_Operator_out155_out1;

  Logical_Operator_out172_out1 <= Logical_Operator_out140_out1 XOR Logical_Operator_out156_out1;

  Logical_Operator_out173_out1 <= Logical_Operator_out141_out1 XOR Logical_Operator_out157_out1;

  Logical_Operator_out174_out1 <= Logical_Operator_out142_out1 XOR Logical_Operator_out158_out1;

  Logical_Operator_out175_out1 <= Logical_Operator_out143_out1 XOR Logical_Operator_out159_out1;

  Logical_Operator_out176_out1 <= Logical_Operator_out144_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out177_out1 <= Logical_Operator_out105_out1 XOR Logical_Operator_out121_out1;

  Logical_Operator_out178_out1 <= Logical_Operator_out106_out1 XOR Logical_Operator_out122_out1;

  Logical_Operator_out179_out1 <= Logical_Operator_out107_out1 XOR Logical_Operator_out123_out1;

  Logical_Operator_out180_out1 <= Logical_Operator_out108_out1 XOR Logical_Operator_out124_out1;

  Logical_Operator_out181_out1 <= Logical_Operator_out109_out1 XOR Logical_Operator_out125_out1;

  Logical_Operator_out182_out1 <= Logical_Operator_out110_out1 XOR Logical_Operator_out126_out1;

  Logical_Operator_out183_out1 <= Logical_Operator_out111_out1 XOR Logical_Operator_out127_out1;

  Logical_Operator_out184_out1 <= Logical_Operator_out112_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out185_out1 <= Logical_Operator_out77_out1 XOR Logical_Operator_out93_out1;

  Logical_Operator_out186_out1 <= Logical_Operator_out78_out1 XOR Logical_Operator_out94_out1;

  Logical_Operator_out187_out1 <= Logical_Operator_out79_out1 XOR Logical_Operator_out95_out1;

  Logical_Operator_out188_out1 <= Logical_Operator_out80_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out189_out1 <= Logical_Operator_out47_out1 XOR Logical_Operator_out63_out1;

  Logical_Operator_out190_out1 <= Logical_Operator_out48_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out191_out1 <= Logical_Operator_out16_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out192_out1 <= in32 XOR in64;

  out1 <= Logical_Operator_out161_out1;

  out2 <= Logical_Operator_out162_out1;

  out3 <= Logical_Operator_out163_out1;

  out4 <= Logical_Operator_out164_out1;

  out5 <= Logical_Operator_out165_out1;

  out6 <= Logical_Operator_out166_out1;

  out7 <= Logical_Operator_out167_out1;

  out8 <= Logical_Operator_out168_out1;

  out9 <= Logical_Operator_out169_out1;

  out10 <= Logical_Operator_out170_out1;

  out11 <= Logical_Operator_out171_out1;

  out12 <= Logical_Operator_out172_out1;

  out13 <= Logical_Operator_out173_out1;

  out14 <= Logical_Operator_out174_out1;

  out15 <= Logical_Operator_out175_out1;

  out16 <= Logical_Operator_out176_out1;

  out17 <= Logical_Operator_out177_out1;

  out18 <= Logical_Operator_out178_out1;

  out19 <= Logical_Operator_out179_out1;

  out20 <= Logical_Operator_out180_out1;

  out21 <= Logical_Operator_out181_out1;

  out22 <= Logical_Operator_out182_out1;

  out23 <= Logical_Operator_out183_out1;

  out24 <= Logical_Operator_out184_out1;

  out25 <= Logical_Operator_out185_out1;

  out26 <= Logical_Operator_out186_out1;

  out27 <= Logical_Operator_out187_out1;

  out28 <= Logical_Operator_out188_out1;

  out29 <= Logical_Operator_out189_out1;

  out30 <= Logical_Operator_out190_out1;

  out31 <= Logical_Operator_out191_out1;

  out32 <= Logical_Operator_out192_out1;

  out33 <= Logical_Operator_out145_out1;

  out34 <= Logical_Operator_out146_out1;

  out35 <= Logical_Operator_out147_out1;

  out36 <= Logical_Operator_out148_out1;

  out37 <= Logical_Operator_out149_out1;

  out38 <= Logical_Operator_out150_out1;

  out39 <= Logical_Operator_out151_out1;

  out40 <= Logical_Operator_out152_out1;

  out41 <= Logical_Operator_out153_out1;

  out42 <= Logical_Operator_out154_out1;

  out43 <= Logical_Operator_out155_out1;

  out44 <= Logical_Operator_out156_out1;

  out45 <= Logical_Operator_out157_out1;

  out46 <= Logical_Operator_out158_out1;

  out47 <= Logical_Operator_out159_out1;

  out48 <= Logical_Operator_out160_out1;

  out49 <= Logical_Operator_out121_out1;

  out50 <= Logical_Operator_out122_out1;

  out51 <= Logical_Operator_out123_out1;

  out52 <= Logical_Operator_out124_out1;

  out53 <= Logical_Operator_out125_out1;

  out54 <= Logical_Operator_out126_out1;

  out55 <= Logical_Operator_out127_out1;

  out56 <= Logical_Operator_out128_out1;

  out57 <= Logical_Operator_out93_out1;

  out58 <= Logical_Operator_out94_out1;

  out59 <= Logical_Operator_out95_out1;

  out60 <= Logical_Operator_out96_out1;

  out61 <= Logical_Operator_out63_out1;

  out62 <= Logical_Operator_out64_out1;

  out63 <= Logical_Operator_out32_out1;

  out64 <= in64;

END rtl;
