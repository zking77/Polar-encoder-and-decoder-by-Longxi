LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY encoderN512 IS
PORT( 
	in1                               :   IN    std_logic;
	in2                               :   IN    std_logic;
	in3                               :   IN    std_logic;
	in4                               :   IN    std_logic;
	in5                               :   IN    std_logic;
	in6                               :   IN    std_logic;
	in7                               :   IN    std_logic;
	in8                               :   IN    std_logic;
	in9                               :   IN    std_logic;
	in10                               :   IN    std_logic;
	in11                               :   IN    std_logic;
	in12                               :   IN    std_logic;
	in13                               :   IN    std_logic;
	in14                               :   IN    std_logic;
	in15                               :   IN    std_logic;
	in16                               :   IN    std_logic;
	in17                               :   IN    std_logic;
	in18                               :   IN    std_logic;
	in19                               :   IN    std_logic;
	in20                               :   IN    std_logic;
	in21                               :   IN    std_logic;
	in22                               :   IN    std_logic;
	in23                               :   IN    std_logic;
	in24                               :   IN    std_logic;
	in25                               :   IN    std_logic;
	in26                               :   IN    std_logic;
	in27                               :   IN    std_logic;
	in28                               :   IN    std_logic;
	in29                               :   IN    std_logic;
	in30                               :   IN    std_logic;
	in31                               :   IN    std_logic;
	in32                               :   IN    std_logic;
	in33                               :   IN    std_logic;
	in34                               :   IN    std_logic;
	in35                               :   IN    std_logic;
	in36                               :   IN    std_logic;
	in37                               :   IN    std_logic;
	in38                               :   IN    std_logic;
	in39                               :   IN    std_logic;
	in40                               :   IN    std_logic;
	in41                               :   IN    std_logic;
	in42                               :   IN    std_logic;
	in43                               :   IN    std_logic;
	in44                               :   IN    std_logic;
	in45                               :   IN    std_logic;
	in46                               :   IN    std_logic;
	in47                               :   IN    std_logic;
	in48                               :   IN    std_logic;
	in49                               :   IN    std_logic;
	in50                               :   IN    std_logic;
	in51                               :   IN    std_logic;
	in52                               :   IN    std_logic;
	in53                               :   IN    std_logic;
	in54                               :   IN    std_logic;
	in55                               :   IN    std_logic;
	in56                               :   IN    std_logic;
	in57                               :   IN    std_logic;
	in58                               :   IN    std_logic;
	in59                               :   IN    std_logic;
	in60                               :   IN    std_logic;
	in61                               :   IN    std_logic;
	in62                               :   IN    std_logic;
	in63                               :   IN    std_logic;
	in64                               :   IN    std_logic;
	in65                               :   IN    std_logic;
	in66                               :   IN    std_logic;
	in67                               :   IN    std_logic;
	in68                               :   IN    std_logic;
	in69                               :   IN    std_logic;
	in70                               :   IN    std_logic;
	in71                               :   IN    std_logic;
	in72                               :   IN    std_logic;
	in73                               :   IN    std_logic;
	in74                               :   IN    std_logic;
	in75                               :   IN    std_logic;
	in76                               :   IN    std_logic;
	in77                               :   IN    std_logic;
	in78                               :   IN    std_logic;
	in79                               :   IN    std_logic;
	in80                               :   IN    std_logic;
	in81                               :   IN    std_logic;
	in82                               :   IN    std_logic;
	in83                               :   IN    std_logic;
	in84                               :   IN    std_logic;
	in85                               :   IN    std_logic;
	in86                               :   IN    std_logic;
	in87                               :   IN    std_logic;
	in88                               :   IN    std_logic;
	in89                               :   IN    std_logic;
	in90                               :   IN    std_logic;
	in91                               :   IN    std_logic;
	in92                               :   IN    std_logic;
	in93                               :   IN    std_logic;
	in94                               :   IN    std_logic;
	in95                               :   IN    std_logic;
	in96                               :   IN    std_logic;
	in97                               :   IN    std_logic;
	in98                               :   IN    std_logic;
	in99                               :   IN    std_logic;
	in100                               :   IN    std_logic;
	in101                               :   IN    std_logic;
	in102                               :   IN    std_logic;
	in103                               :   IN    std_logic;
	in104                               :   IN    std_logic;
	in105                               :   IN    std_logic;
	in106                               :   IN    std_logic;
	in107                               :   IN    std_logic;
	in108                               :   IN    std_logic;
	in109                               :   IN    std_logic;
	in110                               :   IN    std_logic;
	in111                               :   IN    std_logic;
	in112                               :   IN    std_logic;
	in113                               :   IN    std_logic;
	in114                               :   IN    std_logic;
	in115                               :   IN    std_logic;
	in116                               :   IN    std_logic;
	in117                               :   IN    std_logic;
	in118                               :   IN    std_logic;
	in119                               :   IN    std_logic;
	in120                               :   IN    std_logic;
	in121                               :   IN    std_logic;
	in122                               :   IN    std_logic;
	in123                               :   IN    std_logic;
	in124                               :   IN    std_logic;
	in125                               :   IN    std_logic;
	in126                               :   IN    std_logic;
	in127                               :   IN    std_logic;
	in128                               :   IN    std_logic;
	in129                               :   IN    std_logic;
	in130                               :   IN    std_logic;
	in131                               :   IN    std_logic;
	in132                               :   IN    std_logic;
	in133                               :   IN    std_logic;
	in134                               :   IN    std_logic;
	in135                               :   IN    std_logic;
	in136                               :   IN    std_logic;
	in137                               :   IN    std_logic;
	in138                               :   IN    std_logic;
	in139                               :   IN    std_logic;
	in140                               :   IN    std_logic;
	in141                               :   IN    std_logic;
	in142                               :   IN    std_logic;
	in143                               :   IN    std_logic;
	in144                               :   IN    std_logic;
	in145                               :   IN    std_logic;
	in146                               :   IN    std_logic;
	in147                               :   IN    std_logic;
	in148                               :   IN    std_logic;
	in149                               :   IN    std_logic;
	in150                               :   IN    std_logic;
	in151                               :   IN    std_logic;
	in152                               :   IN    std_logic;
	in153                               :   IN    std_logic;
	in154                               :   IN    std_logic;
	in155                               :   IN    std_logic;
	in156                               :   IN    std_logic;
	in157                               :   IN    std_logic;
	in158                               :   IN    std_logic;
	in159                               :   IN    std_logic;
	in160                               :   IN    std_logic;
	in161                               :   IN    std_logic;
	in162                               :   IN    std_logic;
	in163                               :   IN    std_logic;
	in164                               :   IN    std_logic;
	in165                               :   IN    std_logic;
	in166                               :   IN    std_logic;
	in167                               :   IN    std_logic;
	in168                               :   IN    std_logic;
	in169                               :   IN    std_logic;
	in170                               :   IN    std_logic;
	in171                               :   IN    std_logic;
	in172                               :   IN    std_logic;
	in173                               :   IN    std_logic;
	in174                               :   IN    std_logic;
	in175                               :   IN    std_logic;
	in176                               :   IN    std_logic;
	in177                               :   IN    std_logic;
	in178                               :   IN    std_logic;
	in179                               :   IN    std_logic;
	in180                               :   IN    std_logic;
	in181                               :   IN    std_logic;
	in182                               :   IN    std_logic;
	in183                               :   IN    std_logic;
	in184                               :   IN    std_logic;
	in185                               :   IN    std_logic;
	in186                               :   IN    std_logic;
	in187                               :   IN    std_logic;
	in188                               :   IN    std_logic;
	in189                               :   IN    std_logic;
	in190                               :   IN    std_logic;
	in191                               :   IN    std_logic;
	in192                               :   IN    std_logic;
	in193                               :   IN    std_logic;
	in194                               :   IN    std_logic;
	in195                               :   IN    std_logic;
	in196                               :   IN    std_logic;
	in197                               :   IN    std_logic;
	in198                               :   IN    std_logic;
	in199                               :   IN    std_logic;
	in200                               :   IN    std_logic;
	in201                               :   IN    std_logic;
	in202                               :   IN    std_logic;
	in203                               :   IN    std_logic;
	in204                               :   IN    std_logic;
	in205                               :   IN    std_logic;
	in206                               :   IN    std_logic;
	in207                               :   IN    std_logic;
	in208                               :   IN    std_logic;
	in209                               :   IN    std_logic;
	in210                               :   IN    std_logic;
	in211                               :   IN    std_logic;
	in212                               :   IN    std_logic;
	in213                               :   IN    std_logic;
	in214                               :   IN    std_logic;
	in215                               :   IN    std_logic;
	in216                               :   IN    std_logic;
	in217                               :   IN    std_logic;
	in218                               :   IN    std_logic;
	in219                               :   IN    std_logic;
	in220                               :   IN    std_logic;
	in221                               :   IN    std_logic;
	in222                               :   IN    std_logic;
	in223                               :   IN    std_logic;
	in224                               :   IN    std_logic;
	in225                               :   IN    std_logic;
	in226                               :   IN    std_logic;
	in227                               :   IN    std_logic;
	in228                               :   IN    std_logic;
	in229                               :   IN    std_logic;
	in230                               :   IN    std_logic;
	in231                               :   IN    std_logic;
	in232                               :   IN    std_logic;
	in233                               :   IN    std_logic;
	in234                               :   IN    std_logic;
	in235                               :   IN    std_logic;
	in236                               :   IN    std_logic;
	in237                               :   IN    std_logic;
	in238                               :   IN    std_logic;
	in239                               :   IN    std_logic;
	in240                               :   IN    std_logic;
	in241                               :   IN    std_logic;
	in242                               :   IN    std_logic;
	in243                               :   IN    std_logic;
	in244                               :   IN    std_logic;
	in245                               :   IN    std_logic;
	in246                               :   IN    std_logic;
	in247                               :   IN    std_logic;
	in248                               :   IN    std_logic;
	in249                               :   IN    std_logic;
	in250                               :   IN    std_logic;
	in251                               :   IN    std_logic;
	in252                               :   IN    std_logic;
	in253                               :   IN    std_logic;
	in254                               :   IN    std_logic;
	in255                               :   IN    std_logic;
	in256                               :   IN    std_logic;
	in257                               :   IN    std_logic;
	in258                               :   IN    std_logic;
	in259                               :   IN    std_logic;
	in260                               :   IN    std_logic;
	in261                               :   IN    std_logic;
	in262                               :   IN    std_logic;
	in263                               :   IN    std_logic;
	in264                               :   IN    std_logic;
	in265                               :   IN    std_logic;
	in266                               :   IN    std_logic;
	in267                               :   IN    std_logic;
	in268                               :   IN    std_logic;
	in269                               :   IN    std_logic;
	in270                               :   IN    std_logic;
	in271                               :   IN    std_logic;
	in272                               :   IN    std_logic;
	in273                               :   IN    std_logic;
	in274                               :   IN    std_logic;
	in275                               :   IN    std_logic;
	in276                               :   IN    std_logic;
	in277                               :   IN    std_logic;
	in278                               :   IN    std_logic;
	in279                               :   IN    std_logic;
	in280                               :   IN    std_logic;
	in281                               :   IN    std_logic;
	in282                               :   IN    std_logic;
	in283                               :   IN    std_logic;
	in284                               :   IN    std_logic;
	in285                               :   IN    std_logic;
	in286                               :   IN    std_logic;
	in287                               :   IN    std_logic;
	in288                               :   IN    std_logic;
	in289                               :   IN    std_logic;
	in290                               :   IN    std_logic;
	in291                               :   IN    std_logic;
	in292                               :   IN    std_logic;
	in293                               :   IN    std_logic;
	in294                               :   IN    std_logic;
	in295                               :   IN    std_logic;
	in296                               :   IN    std_logic;
	in297                               :   IN    std_logic;
	in298                               :   IN    std_logic;
	in299                               :   IN    std_logic;
	in300                               :   IN    std_logic;
	in301                               :   IN    std_logic;
	in302                               :   IN    std_logic;
	in303                               :   IN    std_logic;
	in304                               :   IN    std_logic;
	in305                               :   IN    std_logic;
	in306                               :   IN    std_logic;
	in307                               :   IN    std_logic;
	in308                               :   IN    std_logic;
	in309                               :   IN    std_logic;
	in310                               :   IN    std_logic;
	in311                               :   IN    std_logic;
	in312                               :   IN    std_logic;
	in313                               :   IN    std_logic;
	in314                               :   IN    std_logic;
	in315                               :   IN    std_logic;
	in316                               :   IN    std_logic;
	in317                               :   IN    std_logic;
	in318                               :   IN    std_logic;
	in319                               :   IN    std_logic;
	in320                               :   IN    std_logic;
	in321                               :   IN    std_logic;
	in322                               :   IN    std_logic;
	in323                               :   IN    std_logic;
	in324                               :   IN    std_logic;
	in325                               :   IN    std_logic;
	in326                               :   IN    std_logic;
	in327                               :   IN    std_logic;
	in328                               :   IN    std_logic;
	in329                               :   IN    std_logic;
	in330                               :   IN    std_logic;
	in331                               :   IN    std_logic;
	in332                               :   IN    std_logic;
	in333                               :   IN    std_logic;
	in334                               :   IN    std_logic;
	in335                               :   IN    std_logic;
	in336                               :   IN    std_logic;
	in337                               :   IN    std_logic;
	in338                               :   IN    std_logic;
	in339                               :   IN    std_logic;
	in340                               :   IN    std_logic;
	in341                               :   IN    std_logic;
	in342                               :   IN    std_logic;
	in343                               :   IN    std_logic;
	in344                               :   IN    std_logic;
	in345                               :   IN    std_logic;
	in346                               :   IN    std_logic;
	in347                               :   IN    std_logic;
	in348                               :   IN    std_logic;
	in349                               :   IN    std_logic;
	in350                               :   IN    std_logic;
	in351                               :   IN    std_logic;
	in352                               :   IN    std_logic;
	in353                               :   IN    std_logic;
	in354                               :   IN    std_logic;
	in355                               :   IN    std_logic;
	in356                               :   IN    std_logic;
	in357                               :   IN    std_logic;
	in358                               :   IN    std_logic;
	in359                               :   IN    std_logic;
	in360                               :   IN    std_logic;
	in361                               :   IN    std_logic;
	in362                               :   IN    std_logic;
	in363                               :   IN    std_logic;
	in364                               :   IN    std_logic;
	in365                               :   IN    std_logic;
	in366                               :   IN    std_logic;
	in367                               :   IN    std_logic;
	in368                               :   IN    std_logic;
	in369                               :   IN    std_logic;
	in370                               :   IN    std_logic;
	in371                               :   IN    std_logic;
	in372                               :   IN    std_logic;
	in373                               :   IN    std_logic;
	in374                               :   IN    std_logic;
	in375                               :   IN    std_logic;
	in376                               :   IN    std_logic;
	in377                               :   IN    std_logic;
	in378                               :   IN    std_logic;
	in379                               :   IN    std_logic;
	in380                               :   IN    std_logic;
	in381                               :   IN    std_logic;
	in382                               :   IN    std_logic;
	in383                               :   IN    std_logic;
	in384                               :   IN    std_logic;
	in385                               :   IN    std_logic;
	in386                               :   IN    std_logic;
	in387                               :   IN    std_logic;
	in388                               :   IN    std_logic;
	in389                               :   IN    std_logic;
	in390                               :   IN    std_logic;
	in391                               :   IN    std_logic;
	in392                               :   IN    std_logic;
	in393                               :   IN    std_logic;
	in394                               :   IN    std_logic;
	in395                               :   IN    std_logic;
	in396                               :   IN    std_logic;
	in397                               :   IN    std_logic;
	in398                               :   IN    std_logic;
	in399                               :   IN    std_logic;
	in400                               :   IN    std_logic;
	in401                               :   IN    std_logic;
	in402                               :   IN    std_logic;
	in403                               :   IN    std_logic;
	in404                               :   IN    std_logic;
	in405                               :   IN    std_logic;
	in406                               :   IN    std_logic;
	in407                               :   IN    std_logic;
	in408                               :   IN    std_logic;
	in409                               :   IN    std_logic;
	in410                               :   IN    std_logic;
	in411                               :   IN    std_logic;
	in412                               :   IN    std_logic;
	in413                               :   IN    std_logic;
	in414                               :   IN    std_logic;
	in415                               :   IN    std_logic;
	in416                               :   IN    std_logic;
	in417                               :   IN    std_logic;
	in418                               :   IN    std_logic;
	in419                               :   IN    std_logic;
	in420                               :   IN    std_logic;
	in421                               :   IN    std_logic;
	in422                               :   IN    std_logic;
	in423                               :   IN    std_logic;
	in424                               :   IN    std_logic;
	in425                               :   IN    std_logic;
	in426                               :   IN    std_logic;
	in427                               :   IN    std_logic;
	in428                               :   IN    std_logic;
	in429                               :   IN    std_logic;
	in430                               :   IN    std_logic;
	in431                               :   IN    std_logic;
	in432                               :   IN    std_logic;
	in433                               :   IN    std_logic;
	in434                               :   IN    std_logic;
	in435                               :   IN    std_logic;
	in436                               :   IN    std_logic;
	in437                               :   IN    std_logic;
	in438                               :   IN    std_logic;
	in439                               :   IN    std_logic;
	in440                               :   IN    std_logic;
	in441                               :   IN    std_logic;
	in442                               :   IN    std_logic;
	in443                               :   IN    std_logic;
	in444                               :   IN    std_logic;
	in445                               :   IN    std_logic;
	in446                               :   IN    std_logic;
	in447                               :   IN    std_logic;
	in448                               :   IN    std_logic;
	in449                               :   IN    std_logic;
	in450                               :   IN    std_logic;
	in451                               :   IN    std_logic;
	in452                               :   IN    std_logic;
	in453                               :   IN    std_logic;
	in454                               :   IN    std_logic;
	in455                               :   IN    std_logic;
	in456                               :   IN    std_logic;
	in457                               :   IN    std_logic;
	in458                               :   IN    std_logic;
	in459                               :   IN    std_logic;
	in460                               :   IN    std_logic;
	in461                               :   IN    std_logic;
	in462                               :   IN    std_logic;
	in463                               :   IN    std_logic;
	in464                               :   IN    std_logic;
	in465                               :   IN    std_logic;
	in466                               :   IN    std_logic;
	in467                               :   IN    std_logic;
	in468                               :   IN    std_logic;
	in469                               :   IN    std_logic;
	in470                               :   IN    std_logic;
	in471                               :   IN    std_logic;
	in472                               :   IN    std_logic;
	in473                               :   IN    std_logic;
	in474                               :   IN    std_logic;
	in475                               :   IN    std_logic;
	in476                               :   IN    std_logic;
	in477                               :   IN    std_logic;
	in478                               :   IN    std_logic;
	in479                               :   IN    std_logic;
	in480                               :   IN    std_logic;
	in481                               :   IN    std_logic;
	in482                               :   IN    std_logic;
	in483                               :   IN    std_logic;
	in484                               :   IN    std_logic;
	in485                               :   IN    std_logic;
	in486                               :   IN    std_logic;
	in487                               :   IN    std_logic;
	in488                               :   IN    std_logic;
	in489                               :   IN    std_logic;
	in490                               :   IN    std_logic;
	in491                               :   IN    std_logic;
	in492                               :   IN    std_logic;
	in493                               :   IN    std_logic;
	in494                               :   IN    std_logic;
	in495                               :   IN    std_logic;
	in496                               :   IN    std_logic;
	in497                               :   IN    std_logic;
	in498                               :   IN    std_logic;
	in499                               :   IN    std_logic;
	in500                               :   IN    std_logic;
	in501                               :   IN    std_logic;
	in502                               :   IN    std_logic;
	in503                               :   IN    std_logic;
	in504                               :   IN    std_logic;
	in505                               :   IN    std_logic;
	in506                               :   IN    std_logic;
	in507                               :   IN    std_logic;
	in508                               :   IN    std_logic;
	in509                               :   IN    std_logic;
	in510                               :   IN    std_logic;
	in511                               :   IN    std_logic;
	in512                               :   IN    std_logic;
	out1                               :   OUT    std_logic;
	out2                               :   OUT    std_logic;
	out3                               :   OUT    std_logic;
	out4                               :   OUT    std_logic;
	out5                               :   OUT    std_logic;
	out6                               :   OUT    std_logic;
	out7                               :   OUT    std_logic;
	out8                               :   OUT    std_logic;
	out9                               :   OUT    std_logic;
	out10                               :   OUT    std_logic;
	out11                               :   OUT    std_logic;
	out12                               :   OUT    std_logic;
	out13                               :   OUT    std_logic;
	out14                               :   OUT    std_logic;
	out15                               :   OUT    std_logic;
	out16                               :   OUT    std_logic;
	out17                               :   OUT    std_logic;
	out18                               :   OUT    std_logic;
	out19                               :   OUT    std_logic;
	out20                               :   OUT    std_logic;
	out21                               :   OUT    std_logic;
	out22                               :   OUT    std_logic;
	out23                               :   OUT    std_logic;
	out24                               :   OUT    std_logic;
	out25                               :   OUT    std_logic;
	out26                               :   OUT    std_logic;
	out27                               :   OUT    std_logic;
	out28                               :   OUT    std_logic;
	out29                               :   OUT    std_logic;
	out30                               :   OUT    std_logic;
	out31                               :   OUT    std_logic;
	out32                               :   OUT    std_logic;
	out33                               :   OUT    std_logic;
	out34                               :   OUT    std_logic;
	out35                               :   OUT    std_logic;
	out36                               :   OUT    std_logic;
	out37                               :   OUT    std_logic;
	out38                               :   OUT    std_logic;
	out39                               :   OUT    std_logic;
	out40                               :   OUT    std_logic;
	out41                               :   OUT    std_logic;
	out42                               :   OUT    std_logic;
	out43                               :   OUT    std_logic;
	out44                               :   OUT    std_logic;
	out45                               :   OUT    std_logic;
	out46                               :   OUT    std_logic;
	out47                               :   OUT    std_logic;
	out48                               :   OUT    std_logic;
	out49                               :   OUT    std_logic;
	out50                               :   OUT    std_logic;
	out51                               :   OUT    std_logic;
	out52                               :   OUT    std_logic;
	out53                               :   OUT    std_logic;
	out54                               :   OUT    std_logic;
	out55                               :   OUT    std_logic;
	out56                               :   OUT    std_logic;
	out57                               :   OUT    std_logic;
	out58                               :   OUT    std_logic;
	out59                               :   OUT    std_logic;
	out60                               :   OUT    std_logic;
	out61                               :   OUT    std_logic;
	out62                               :   OUT    std_logic;
	out63                               :   OUT    std_logic;
	out64                               :   OUT    std_logic;
	out65                               :   OUT    std_logic;
	out66                               :   OUT    std_logic;
	out67                               :   OUT    std_logic;
	out68                               :   OUT    std_logic;
	out69                               :   OUT    std_logic;
	out70                               :   OUT    std_logic;
	out71                               :   OUT    std_logic;
	out72                               :   OUT    std_logic;
	out73                               :   OUT    std_logic;
	out74                               :   OUT    std_logic;
	out75                               :   OUT    std_logic;
	out76                               :   OUT    std_logic;
	out77                               :   OUT    std_logic;
	out78                               :   OUT    std_logic;
	out79                               :   OUT    std_logic;
	out80                               :   OUT    std_logic;
	out81                               :   OUT    std_logic;
	out82                               :   OUT    std_logic;
	out83                               :   OUT    std_logic;
	out84                               :   OUT    std_logic;
	out85                               :   OUT    std_logic;
	out86                               :   OUT    std_logic;
	out87                               :   OUT    std_logic;
	out88                               :   OUT    std_logic;
	out89                               :   OUT    std_logic;
	out90                               :   OUT    std_logic;
	out91                               :   OUT    std_logic;
	out92                               :   OUT    std_logic;
	out93                               :   OUT    std_logic;
	out94                               :   OUT    std_logic;
	out95                               :   OUT    std_logic;
	out96                               :   OUT    std_logic;
	out97                               :   OUT    std_logic;
	out98                               :   OUT    std_logic;
	out99                               :   OUT    std_logic;
	out100                               :   OUT    std_logic;
	out101                               :   OUT    std_logic;
	out102                               :   OUT    std_logic;
	out103                               :   OUT    std_logic;
	out104                               :   OUT    std_logic;
	out105                               :   OUT    std_logic;
	out106                               :   OUT    std_logic;
	out107                               :   OUT    std_logic;
	out108                               :   OUT    std_logic;
	out109                               :   OUT    std_logic;
	out110                               :   OUT    std_logic;
	out111                               :   OUT    std_logic;
	out112                               :   OUT    std_logic;
	out113                               :   OUT    std_logic;
	out114                               :   OUT    std_logic;
	out115                               :   OUT    std_logic;
	out116                               :   OUT    std_logic;
	out117                               :   OUT    std_logic;
	out118                               :   OUT    std_logic;
	out119                               :   OUT    std_logic;
	out120                               :   OUT    std_logic;
	out121                               :   OUT    std_logic;
	out122                               :   OUT    std_logic;
	out123                               :   OUT    std_logic;
	out124                               :   OUT    std_logic;
	out125                               :   OUT    std_logic;
	out126                               :   OUT    std_logic;
	out127                               :   OUT    std_logic;
	out128                               :   OUT    std_logic;
	out129                               :   OUT    std_logic;
	out130                               :   OUT    std_logic;
	out131                               :   OUT    std_logic;
	out132                               :   OUT    std_logic;
	out133                               :   OUT    std_logic;
	out134                               :   OUT    std_logic;
	out135                               :   OUT    std_logic;
	out136                               :   OUT    std_logic;
	out137                               :   OUT    std_logic;
	out138                               :   OUT    std_logic;
	out139                               :   OUT    std_logic;
	out140                               :   OUT    std_logic;
	out141                               :   OUT    std_logic;
	out142                               :   OUT    std_logic;
	out143                               :   OUT    std_logic;
	out144                               :   OUT    std_logic;
	out145                               :   OUT    std_logic;
	out146                               :   OUT    std_logic;
	out147                               :   OUT    std_logic;
	out148                               :   OUT    std_logic;
	out149                               :   OUT    std_logic;
	out150                               :   OUT    std_logic;
	out151                               :   OUT    std_logic;
	out152                               :   OUT    std_logic;
	out153                               :   OUT    std_logic;
	out154                               :   OUT    std_logic;
	out155                               :   OUT    std_logic;
	out156                               :   OUT    std_logic;
	out157                               :   OUT    std_logic;
	out158                               :   OUT    std_logic;
	out159                               :   OUT    std_logic;
	out160                               :   OUT    std_logic;
	out161                               :   OUT    std_logic;
	out162                               :   OUT    std_logic;
	out163                               :   OUT    std_logic;
	out164                               :   OUT    std_logic;
	out165                               :   OUT    std_logic;
	out166                               :   OUT    std_logic;
	out167                               :   OUT    std_logic;
	out168                               :   OUT    std_logic;
	out169                               :   OUT    std_logic;
	out170                               :   OUT    std_logic;
	out171                               :   OUT    std_logic;
	out172                               :   OUT    std_logic;
	out173                               :   OUT    std_logic;
	out174                               :   OUT    std_logic;
	out175                               :   OUT    std_logic;
	out176                               :   OUT    std_logic;
	out177                               :   OUT    std_logic;
	out178                               :   OUT    std_logic;
	out179                               :   OUT    std_logic;
	out180                               :   OUT    std_logic;
	out181                               :   OUT    std_logic;
	out182                               :   OUT    std_logic;
	out183                               :   OUT    std_logic;
	out184                               :   OUT    std_logic;
	out185                               :   OUT    std_logic;
	out186                               :   OUT    std_logic;
	out187                               :   OUT    std_logic;
	out188                               :   OUT    std_logic;
	out189                               :   OUT    std_logic;
	out190                               :   OUT    std_logic;
	out191                               :   OUT    std_logic;
	out192                               :   OUT    std_logic;
	out193                               :   OUT    std_logic;
	out194                               :   OUT    std_logic;
	out195                               :   OUT    std_logic;
	out196                               :   OUT    std_logic;
	out197                               :   OUT    std_logic;
	out198                               :   OUT    std_logic;
	out199                               :   OUT    std_logic;
	out200                               :   OUT    std_logic;
	out201                               :   OUT    std_logic;
	out202                               :   OUT    std_logic;
	out203                               :   OUT    std_logic;
	out204                               :   OUT    std_logic;
	out205                               :   OUT    std_logic;
	out206                               :   OUT    std_logic;
	out207                               :   OUT    std_logic;
	out208                               :   OUT    std_logic;
	out209                               :   OUT    std_logic;
	out210                               :   OUT    std_logic;
	out211                               :   OUT    std_logic;
	out212                               :   OUT    std_logic;
	out213                               :   OUT    std_logic;
	out214                               :   OUT    std_logic;
	out215                               :   OUT    std_logic;
	out216                               :   OUT    std_logic;
	out217                               :   OUT    std_logic;
	out218                               :   OUT    std_logic;
	out219                               :   OUT    std_logic;
	out220                               :   OUT    std_logic;
	out221                               :   OUT    std_logic;
	out222                               :   OUT    std_logic;
	out223                               :   OUT    std_logic;
	out224                               :   OUT    std_logic;
	out225                               :   OUT    std_logic;
	out226                               :   OUT    std_logic;
	out227                               :   OUT    std_logic;
	out228                               :   OUT    std_logic;
	out229                               :   OUT    std_logic;
	out230                               :   OUT    std_logic;
	out231                               :   OUT    std_logic;
	out232                               :   OUT    std_logic;
	out233                               :   OUT    std_logic;
	out234                               :   OUT    std_logic;
	out235                               :   OUT    std_logic;
	out236                               :   OUT    std_logic;
	out237                               :   OUT    std_logic;
	out238                               :   OUT    std_logic;
	out239                               :   OUT    std_logic;
	out240                               :   OUT    std_logic;
	out241                               :   OUT    std_logic;
	out242                               :   OUT    std_logic;
	out243                               :   OUT    std_logic;
	out244                               :   OUT    std_logic;
	out245                               :   OUT    std_logic;
	out246                               :   OUT    std_logic;
	out247                               :   OUT    std_logic;
	out248                               :   OUT    std_logic;
	out249                               :   OUT    std_logic;
	out250                               :   OUT    std_logic;
	out251                               :   OUT    std_logic;
	out252                               :   OUT    std_logic;
	out253                               :   OUT    std_logic;
	out254                               :   OUT    std_logic;
	out255                               :   OUT    std_logic;
	out256                               :   OUT    std_logic;
	out257                               :   OUT    std_logic;
	out258                               :   OUT    std_logic;
	out259                               :   OUT    std_logic;
	out260                               :   OUT    std_logic;
	out261                               :   OUT    std_logic;
	out262                               :   OUT    std_logic;
	out263                               :   OUT    std_logic;
	out264                               :   OUT    std_logic;
	out265                               :   OUT    std_logic;
	out266                               :   OUT    std_logic;
	out267                               :   OUT    std_logic;
	out268                               :   OUT    std_logic;
	out269                               :   OUT    std_logic;
	out270                               :   OUT    std_logic;
	out271                               :   OUT    std_logic;
	out272                               :   OUT    std_logic;
	out273                               :   OUT    std_logic;
	out274                               :   OUT    std_logic;
	out275                               :   OUT    std_logic;
	out276                               :   OUT    std_logic;
	out277                               :   OUT    std_logic;
	out278                               :   OUT    std_logic;
	out279                               :   OUT    std_logic;
	out280                               :   OUT    std_logic;
	out281                               :   OUT    std_logic;
	out282                               :   OUT    std_logic;
	out283                               :   OUT    std_logic;
	out284                               :   OUT    std_logic;
	out285                               :   OUT    std_logic;
	out286                               :   OUT    std_logic;
	out287                               :   OUT    std_logic;
	out288                               :   OUT    std_logic;
	out289                               :   OUT    std_logic;
	out290                               :   OUT    std_logic;
	out291                               :   OUT    std_logic;
	out292                               :   OUT    std_logic;
	out293                               :   OUT    std_logic;
	out294                               :   OUT    std_logic;
	out295                               :   OUT    std_logic;
	out296                               :   OUT    std_logic;
	out297                               :   OUT    std_logic;
	out298                               :   OUT    std_logic;
	out299                               :   OUT    std_logic;
	out300                               :   OUT    std_logic;
	out301                               :   OUT    std_logic;
	out302                               :   OUT    std_logic;
	out303                               :   OUT    std_logic;
	out304                               :   OUT    std_logic;
	out305                               :   OUT    std_logic;
	out306                               :   OUT    std_logic;
	out307                               :   OUT    std_logic;
	out308                               :   OUT    std_logic;
	out309                               :   OUT    std_logic;
	out310                               :   OUT    std_logic;
	out311                               :   OUT    std_logic;
	out312                               :   OUT    std_logic;
	out313                               :   OUT    std_logic;
	out314                               :   OUT    std_logic;
	out315                               :   OUT    std_logic;
	out316                               :   OUT    std_logic;
	out317                               :   OUT    std_logic;
	out318                               :   OUT    std_logic;
	out319                               :   OUT    std_logic;
	out320                               :   OUT    std_logic;
	out321                               :   OUT    std_logic;
	out322                               :   OUT    std_logic;
	out323                               :   OUT    std_logic;
	out324                               :   OUT    std_logic;
	out325                               :   OUT    std_logic;
	out326                               :   OUT    std_logic;
	out327                               :   OUT    std_logic;
	out328                               :   OUT    std_logic;
	out329                               :   OUT    std_logic;
	out330                               :   OUT    std_logic;
	out331                               :   OUT    std_logic;
	out332                               :   OUT    std_logic;
	out333                               :   OUT    std_logic;
	out334                               :   OUT    std_logic;
	out335                               :   OUT    std_logic;
	out336                               :   OUT    std_logic;
	out337                               :   OUT    std_logic;
	out338                               :   OUT    std_logic;
	out339                               :   OUT    std_logic;
	out340                               :   OUT    std_logic;
	out341                               :   OUT    std_logic;
	out342                               :   OUT    std_logic;
	out343                               :   OUT    std_logic;
	out344                               :   OUT    std_logic;
	out345                               :   OUT    std_logic;
	out346                               :   OUT    std_logic;
	out347                               :   OUT    std_logic;
	out348                               :   OUT    std_logic;
	out349                               :   OUT    std_logic;
	out350                               :   OUT    std_logic;
	out351                               :   OUT    std_logic;
	out352                               :   OUT    std_logic;
	out353                               :   OUT    std_logic;
	out354                               :   OUT    std_logic;
	out355                               :   OUT    std_logic;
	out356                               :   OUT    std_logic;
	out357                               :   OUT    std_logic;
	out358                               :   OUT    std_logic;
	out359                               :   OUT    std_logic;
	out360                               :   OUT    std_logic;
	out361                               :   OUT    std_logic;
	out362                               :   OUT    std_logic;
	out363                               :   OUT    std_logic;
	out364                               :   OUT    std_logic;
	out365                               :   OUT    std_logic;
	out366                               :   OUT    std_logic;
	out367                               :   OUT    std_logic;
	out368                               :   OUT    std_logic;
	out369                               :   OUT    std_logic;
	out370                               :   OUT    std_logic;
	out371                               :   OUT    std_logic;
	out372                               :   OUT    std_logic;
	out373                               :   OUT    std_logic;
	out374                               :   OUT    std_logic;
	out375                               :   OUT    std_logic;
	out376                               :   OUT    std_logic;
	out377                               :   OUT    std_logic;
	out378                               :   OUT    std_logic;
	out379                               :   OUT    std_logic;
	out380                               :   OUT    std_logic;
	out381                               :   OUT    std_logic;
	out382                               :   OUT    std_logic;
	out383                               :   OUT    std_logic;
	out384                               :   OUT    std_logic;
	out385                               :   OUT    std_logic;
	out386                               :   OUT    std_logic;
	out387                               :   OUT    std_logic;
	out388                               :   OUT    std_logic;
	out389                               :   OUT    std_logic;
	out390                               :   OUT    std_logic;
	out391                               :   OUT    std_logic;
	out392                               :   OUT    std_logic;
	out393                               :   OUT    std_logic;
	out394                               :   OUT    std_logic;
	out395                               :   OUT    std_logic;
	out396                               :   OUT    std_logic;
	out397                               :   OUT    std_logic;
	out398                               :   OUT    std_logic;
	out399                               :   OUT    std_logic;
	out400                               :   OUT    std_logic;
	out401                               :   OUT    std_logic;
	out402                               :   OUT    std_logic;
	out403                               :   OUT    std_logic;
	out404                               :   OUT    std_logic;
	out405                               :   OUT    std_logic;
	out406                               :   OUT    std_logic;
	out407                               :   OUT    std_logic;
	out408                               :   OUT    std_logic;
	out409                               :   OUT    std_logic;
	out410                               :   OUT    std_logic;
	out411                               :   OUT    std_logic;
	out412                               :   OUT    std_logic;
	out413                               :   OUT    std_logic;
	out414                               :   OUT    std_logic;
	out415                               :   OUT    std_logic;
	out416                               :   OUT    std_logic;
	out417                               :   OUT    std_logic;
	out418                               :   OUT    std_logic;
	out419                               :   OUT    std_logic;
	out420                               :   OUT    std_logic;
	out421                               :   OUT    std_logic;
	out422                               :   OUT    std_logic;
	out423                               :   OUT    std_logic;
	out424                               :   OUT    std_logic;
	out425                               :   OUT    std_logic;
	out426                               :   OUT    std_logic;
	out427                               :   OUT    std_logic;
	out428                               :   OUT    std_logic;
	out429                               :   OUT    std_logic;
	out430                               :   OUT    std_logic;
	out431                               :   OUT    std_logic;
	out432                               :   OUT    std_logic;
	out433                               :   OUT    std_logic;
	out434                               :   OUT    std_logic;
	out435                               :   OUT    std_logic;
	out436                               :   OUT    std_logic;
	out437                               :   OUT    std_logic;
	out438                               :   OUT    std_logic;
	out439                               :   OUT    std_logic;
	out440                               :   OUT    std_logic;
	out441                               :   OUT    std_logic;
	out442                               :   OUT    std_logic;
	out443                               :   OUT    std_logic;
	out444                               :   OUT    std_logic;
	out445                               :   OUT    std_logic;
	out446                               :   OUT    std_logic;
	out447                               :   OUT    std_logic;
	out448                               :   OUT    std_logic;
	out449                               :   OUT    std_logic;
	out450                               :   OUT    std_logic;
	out451                               :   OUT    std_logic;
	out452                               :   OUT    std_logic;
	out453                               :   OUT    std_logic;
	out454                               :   OUT    std_logic;
	out455                               :   OUT    std_logic;
	out456                               :   OUT    std_logic;
	out457                               :   OUT    std_logic;
	out458                               :   OUT    std_logic;
	out459                               :   OUT    std_logic;
	out460                               :   OUT    std_logic;
	out461                               :   OUT    std_logic;
	out462                               :   OUT    std_logic;
	out463                               :   OUT    std_logic;
	out464                               :   OUT    std_logic;
	out465                               :   OUT    std_logic;
	out466                               :   OUT    std_logic;
	out467                               :   OUT    std_logic;
	out468                               :   OUT    std_logic;
	out469                               :   OUT    std_logic;
	out470                               :   OUT    std_logic;
	out471                               :   OUT    std_logic;
	out472                               :   OUT    std_logic;
	out473                               :   OUT    std_logic;
	out474                               :   OUT    std_logic;
	out475                               :   OUT    std_logic;
	out476                               :   OUT    std_logic;
	out477                               :   OUT    std_logic;
	out478                               :   OUT    std_logic;
	out479                               :   OUT    std_logic;
	out480                               :   OUT    std_logic;
	out481                               :   OUT    std_logic;
	out482                               :   OUT    std_logic;
	out483                               :   OUT    std_logic;
	out484                               :   OUT    std_logic;
	out485                               :   OUT    std_logic;
	out486                               :   OUT    std_logic;
	out487                               :   OUT    std_logic;
	out488                               :   OUT    std_logic;
	out489                               :   OUT    std_logic;
	out490                               :   OUT    std_logic;
	out491                               :   OUT    std_logic;
	out492                               :   OUT    std_logic;
	out493                               :   OUT    std_logic;
	out494                               :   OUT    std_logic;
	out495                               :   OUT    std_logic;
	out496                               :   OUT    std_logic;
	out497                               :   OUT    std_logic;
	out498                               :   OUT    std_logic;
	out499                               :   OUT    std_logic;
	out500                               :   OUT    std_logic;
	out501                               :   OUT    std_logic;
	out502                               :   OUT    std_logic;
	out503                               :   OUT    std_logic;
	out504                               :   OUT    std_logic;
	out505                               :   OUT    std_logic;
	out506                               :   OUT    std_logic;
	out507                               :   OUT    std_logic;
	out508                               :   OUT    std_logic;
	out509                               :   OUT    std_logic;
	out510                               :   OUT    std_logic;
	out511                               :   OUT    std_logic;
	out512                               :   OUT    std_logic
	);
END encoderN512;

ARCHITECTURE rtl OF encoderN512 IS

  SIGNAL Logical_Operator_out1_out1            : std_logic;
  SIGNAL Logical_Operator_out2_out1            : std_logic;
  SIGNAL Logical_Operator_out3_out1            : std_logic;
  SIGNAL Logical_Operator_out4_out1            : std_logic;
  SIGNAL Logical_Operator_out5_out1            : std_logic;
  SIGNAL Logical_Operator_out6_out1            : std_logic;
  SIGNAL Logical_Operator_out7_out1            : std_logic;
  SIGNAL Logical_Operator_out8_out1            : std_logic;
  SIGNAL Logical_Operator_out9_out1            : std_logic;
  SIGNAL Logical_Operator_out10_out1            : std_logic;
  SIGNAL Logical_Operator_out11_out1            : std_logic;
  SIGNAL Logical_Operator_out12_out1            : std_logic;
  SIGNAL Logical_Operator_out13_out1            : std_logic;
  SIGNAL Logical_Operator_out14_out1            : std_logic;
  SIGNAL Logical_Operator_out15_out1            : std_logic;
  SIGNAL Logical_Operator_out16_out1            : std_logic;
  SIGNAL Logical_Operator_out17_out1            : std_logic;
  SIGNAL Logical_Operator_out18_out1            : std_logic;
  SIGNAL Logical_Operator_out19_out1            : std_logic;
  SIGNAL Logical_Operator_out20_out1            : std_logic;
  SIGNAL Logical_Operator_out21_out1            : std_logic;
  SIGNAL Logical_Operator_out22_out1            : std_logic;
  SIGNAL Logical_Operator_out23_out1            : std_logic;
  SIGNAL Logical_Operator_out24_out1            : std_logic;
  SIGNAL Logical_Operator_out25_out1            : std_logic;
  SIGNAL Logical_Operator_out26_out1            : std_logic;
  SIGNAL Logical_Operator_out27_out1            : std_logic;
  SIGNAL Logical_Operator_out28_out1            : std_logic;
  SIGNAL Logical_Operator_out29_out1            : std_logic;
  SIGNAL Logical_Operator_out30_out1            : std_logic;
  SIGNAL Logical_Operator_out31_out1            : std_logic;
  SIGNAL Logical_Operator_out32_out1            : std_logic;
  SIGNAL Logical_Operator_out33_out1            : std_logic;
  SIGNAL Logical_Operator_out34_out1            : std_logic;
  SIGNAL Logical_Operator_out35_out1            : std_logic;
  SIGNAL Logical_Operator_out36_out1            : std_logic;
  SIGNAL Logical_Operator_out37_out1            : std_logic;
  SIGNAL Logical_Operator_out38_out1            : std_logic;
  SIGNAL Logical_Operator_out39_out1            : std_logic;
  SIGNAL Logical_Operator_out40_out1            : std_logic;
  SIGNAL Logical_Operator_out41_out1            : std_logic;
  SIGNAL Logical_Operator_out42_out1            : std_logic;
  SIGNAL Logical_Operator_out43_out1            : std_logic;
  SIGNAL Logical_Operator_out44_out1            : std_logic;
  SIGNAL Logical_Operator_out45_out1            : std_logic;
  SIGNAL Logical_Operator_out46_out1            : std_logic;
  SIGNAL Logical_Operator_out47_out1            : std_logic;
  SIGNAL Logical_Operator_out48_out1            : std_logic;
  SIGNAL Logical_Operator_out49_out1            : std_logic;
  SIGNAL Logical_Operator_out50_out1            : std_logic;
  SIGNAL Logical_Operator_out51_out1            : std_logic;
  SIGNAL Logical_Operator_out52_out1            : std_logic;
  SIGNAL Logical_Operator_out53_out1            : std_logic;
  SIGNAL Logical_Operator_out54_out1            : std_logic;
  SIGNAL Logical_Operator_out55_out1            : std_logic;
  SIGNAL Logical_Operator_out56_out1            : std_logic;
  SIGNAL Logical_Operator_out57_out1            : std_logic;
  SIGNAL Logical_Operator_out58_out1            : std_logic;
  SIGNAL Logical_Operator_out59_out1            : std_logic;
  SIGNAL Logical_Operator_out60_out1            : std_logic;
  SIGNAL Logical_Operator_out61_out1            : std_logic;
  SIGNAL Logical_Operator_out62_out1            : std_logic;
  SIGNAL Logical_Operator_out63_out1            : std_logic;
  SIGNAL Logical_Operator_out64_out1            : std_logic;
  SIGNAL Logical_Operator_out65_out1            : std_logic;
  SIGNAL Logical_Operator_out66_out1            : std_logic;
  SIGNAL Logical_Operator_out67_out1            : std_logic;
  SIGNAL Logical_Operator_out68_out1            : std_logic;
  SIGNAL Logical_Operator_out69_out1            : std_logic;
  SIGNAL Logical_Operator_out70_out1            : std_logic;
  SIGNAL Logical_Operator_out71_out1            : std_logic;
  SIGNAL Logical_Operator_out72_out1            : std_logic;
  SIGNAL Logical_Operator_out73_out1            : std_logic;
  SIGNAL Logical_Operator_out74_out1            : std_logic;
  SIGNAL Logical_Operator_out75_out1            : std_logic;
  SIGNAL Logical_Operator_out76_out1            : std_logic;
  SIGNAL Logical_Operator_out77_out1            : std_logic;
  SIGNAL Logical_Operator_out78_out1            : std_logic;
  SIGNAL Logical_Operator_out79_out1            : std_logic;
  SIGNAL Logical_Operator_out80_out1            : std_logic;
  SIGNAL Logical_Operator_out81_out1            : std_logic;
  SIGNAL Logical_Operator_out82_out1            : std_logic;
  SIGNAL Logical_Operator_out83_out1            : std_logic;
  SIGNAL Logical_Operator_out84_out1            : std_logic;
  SIGNAL Logical_Operator_out85_out1            : std_logic;
  SIGNAL Logical_Operator_out86_out1            : std_logic;
  SIGNAL Logical_Operator_out87_out1            : std_logic;
  SIGNAL Logical_Operator_out88_out1            : std_logic;
  SIGNAL Logical_Operator_out89_out1            : std_logic;
  SIGNAL Logical_Operator_out90_out1            : std_logic;
  SIGNAL Logical_Operator_out91_out1            : std_logic;
  SIGNAL Logical_Operator_out92_out1            : std_logic;
  SIGNAL Logical_Operator_out93_out1            : std_logic;
  SIGNAL Logical_Operator_out94_out1            : std_logic;
  SIGNAL Logical_Operator_out95_out1            : std_logic;
  SIGNAL Logical_Operator_out96_out1            : std_logic;
  SIGNAL Logical_Operator_out97_out1            : std_logic;
  SIGNAL Logical_Operator_out98_out1            : std_logic;
  SIGNAL Logical_Operator_out99_out1            : std_logic;
  SIGNAL Logical_Operator_out100_out1            : std_logic;
  SIGNAL Logical_Operator_out101_out1            : std_logic;
  SIGNAL Logical_Operator_out102_out1            : std_logic;
  SIGNAL Logical_Operator_out103_out1            : std_logic;
  SIGNAL Logical_Operator_out104_out1            : std_logic;
  SIGNAL Logical_Operator_out105_out1            : std_logic;
  SIGNAL Logical_Operator_out106_out1            : std_logic;
  SIGNAL Logical_Operator_out107_out1            : std_logic;
  SIGNAL Logical_Operator_out108_out1            : std_logic;
  SIGNAL Logical_Operator_out109_out1            : std_logic;
  SIGNAL Logical_Operator_out110_out1            : std_logic;
  SIGNAL Logical_Operator_out111_out1            : std_logic;
  SIGNAL Logical_Operator_out112_out1            : std_logic;
  SIGNAL Logical_Operator_out113_out1            : std_logic;
  SIGNAL Logical_Operator_out114_out1            : std_logic;
  SIGNAL Logical_Operator_out115_out1            : std_logic;
  SIGNAL Logical_Operator_out116_out1            : std_logic;
  SIGNAL Logical_Operator_out117_out1            : std_logic;
  SIGNAL Logical_Operator_out118_out1            : std_logic;
  SIGNAL Logical_Operator_out119_out1            : std_logic;
  SIGNAL Logical_Operator_out120_out1            : std_logic;
  SIGNAL Logical_Operator_out121_out1            : std_logic;
  SIGNAL Logical_Operator_out122_out1            : std_logic;
  SIGNAL Logical_Operator_out123_out1            : std_logic;
  SIGNAL Logical_Operator_out124_out1            : std_logic;
  SIGNAL Logical_Operator_out125_out1            : std_logic;
  SIGNAL Logical_Operator_out126_out1            : std_logic;
  SIGNAL Logical_Operator_out127_out1            : std_logic;
  SIGNAL Logical_Operator_out128_out1            : std_logic;
  SIGNAL Logical_Operator_out129_out1            : std_logic;
  SIGNAL Logical_Operator_out130_out1            : std_logic;
  SIGNAL Logical_Operator_out131_out1            : std_logic;
  SIGNAL Logical_Operator_out132_out1            : std_logic;
  SIGNAL Logical_Operator_out133_out1            : std_logic;
  SIGNAL Logical_Operator_out134_out1            : std_logic;
  SIGNAL Logical_Operator_out135_out1            : std_logic;
  SIGNAL Logical_Operator_out136_out1            : std_logic;
  SIGNAL Logical_Operator_out137_out1            : std_logic;
  SIGNAL Logical_Operator_out138_out1            : std_logic;
  SIGNAL Logical_Operator_out139_out1            : std_logic;
  SIGNAL Logical_Operator_out140_out1            : std_logic;
  SIGNAL Logical_Operator_out141_out1            : std_logic;
  SIGNAL Logical_Operator_out142_out1            : std_logic;
  SIGNAL Logical_Operator_out143_out1            : std_logic;
  SIGNAL Logical_Operator_out144_out1            : std_logic;
  SIGNAL Logical_Operator_out145_out1            : std_logic;
  SIGNAL Logical_Operator_out146_out1            : std_logic;
  SIGNAL Logical_Operator_out147_out1            : std_logic;
  SIGNAL Logical_Operator_out148_out1            : std_logic;
  SIGNAL Logical_Operator_out149_out1            : std_logic;
  SIGNAL Logical_Operator_out150_out1            : std_logic;
  SIGNAL Logical_Operator_out151_out1            : std_logic;
  SIGNAL Logical_Operator_out152_out1            : std_logic;
  SIGNAL Logical_Operator_out153_out1            : std_logic;
  SIGNAL Logical_Operator_out154_out1            : std_logic;
  SIGNAL Logical_Operator_out155_out1            : std_logic;
  SIGNAL Logical_Operator_out156_out1            : std_logic;
  SIGNAL Logical_Operator_out157_out1            : std_logic;
  SIGNAL Logical_Operator_out158_out1            : std_logic;
  SIGNAL Logical_Operator_out159_out1            : std_logic;
  SIGNAL Logical_Operator_out160_out1            : std_logic;
  SIGNAL Logical_Operator_out161_out1            : std_logic;
  SIGNAL Logical_Operator_out162_out1            : std_logic;
  SIGNAL Logical_Operator_out163_out1            : std_logic;
  SIGNAL Logical_Operator_out164_out1            : std_logic;
  SIGNAL Logical_Operator_out165_out1            : std_logic;
  SIGNAL Logical_Operator_out166_out1            : std_logic;
  SIGNAL Logical_Operator_out167_out1            : std_logic;
  SIGNAL Logical_Operator_out168_out1            : std_logic;
  SIGNAL Logical_Operator_out169_out1            : std_logic;
  SIGNAL Logical_Operator_out170_out1            : std_logic;
  SIGNAL Logical_Operator_out171_out1            : std_logic;
  SIGNAL Logical_Operator_out172_out1            : std_logic;
  SIGNAL Logical_Operator_out173_out1            : std_logic;
  SIGNAL Logical_Operator_out174_out1            : std_logic;
  SIGNAL Logical_Operator_out175_out1            : std_logic;
  SIGNAL Logical_Operator_out176_out1            : std_logic;
  SIGNAL Logical_Operator_out177_out1            : std_logic;
  SIGNAL Logical_Operator_out178_out1            : std_logic;
  SIGNAL Logical_Operator_out179_out1            : std_logic;
  SIGNAL Logical_Operator_out180_out1            : std_logic;
  SIGNAL Logical_Operator_out181_out1            : std_logic;
  SIGNAL Logical_Operator_out182_out1            : std_logic;
  SIGNAL Logical_Operator_out183_out1            : std_logic;
  SIGNAL Logical_Operator_out184_out1            : std_logic;
  SIGNAL Logical_Operator_out185_out1            : std_logic;
  SIGNAL Logical_Operator_out186_out1            : std_logic;
  SIGNAL Logical_Operator_out187_out1            : std_logic;
  SIGNAL Logical_Operator_out188_out1            : std_logic;
  SIGNAL Logical_Operator_out189_out1            : std_logic;
  SIGNAL Logical_Operator_out190_out1            : std_logic;
  SIGNAL Logical_Operator_out191_out1            : std_logic;
  SIGNAL Logical_Operator_out192_out1            : std_logic;
  SIGNAL Logical_Operator_out193_out1            : std_logic;
  SIGNAL Logical_Operator_out194_out1            : std_logic;
  SIGNAL Logical_Operator_out195_out1            : std_logic;
  SIGNAL Logical_Operator_out196_out1            : std_logic;
  SIGNAL Logical_Operator_out197_out1            : std_logic;
  SIGNAL Logical_Operator_out198_out1            : std_logic;
  SIGNAL Logical_Operator_out199_out1            : std_logic;
  SIGNAL Logical_Operator_out200_out1            : std_logic;
  SIGNAL Logical_Operator_out201_out1            : std_logic;
  SIGNAL Logical_Operator_out202_out1            : std_logic;
  SIGNAL Logical_Operator_out203_out1            : std_logic;
  SIGNAL Logical_Operator_out204_out1            : std_logic;
  SIGNAL Logical_Operator_out205_out1            : std_logic;
  SIGNAL Logical_Operator_out206_out1            : std_logic;
  SIGNAL Logical_Operator_out207_out1            : std_logic;
  SIGNAL Logical_Operator_out208_out1            : std_logic;
  SIGNAL Logical_Operator_out209_out1            : std_logic;
  SIGNAL Logical_Operator_out210_out1            : std_logic;
  SIGNAL Logical_Operator_out211_out1            : std_logic;
  SIGNAL Logical_Operator_out212_out1            : std_logic;
  SIGNAL Logical_Operator_out213_out1            : std_logic;
  SIGNAL Logical_Operator_out214_out1            : std_logic;
  SIGNAL Logical_Operator_out215_out1            : std_logic;
  SIGNAL Logical_Operator_out216_out1            : std_logic;
  SIGNAL Logical_Operator_out217_out1            : std_logic;
  SIGNAL Logical_Operator_out218_out1            : std_logic;
  SIGNAL Logical_Operator_out219_out1            : std_logic;
  SIGNAL Logical_Operator_out220_out1            : std_logic;
  SIGNAL Logical_Operator_out221_out1            : std_logic;
  SIGNAL Logical_Operator_out222_out1            : std_logic;
  SIGNAL Logical_Operator_out223_out1            : std_logic;
  SIGNAL Logical_Operator_out224_out1            : std_logic;
  SIGNAL Logical_Operator_out225_out1            : std_logic;
  SIGNAL Logical_Operator_out226_out1            : std_logic;
  SIGNAL Logical_Operator_out227_out1            : std_logic;
  SIGNAL Logical_Operator_out228_out1            : std_logic;
  SIGNAL Logical_Operator_out229_out1            : std_logic;
  SIGNAL Logical_Operator_out230_out1            : std_logic;
  SIGNAL Logical_Operator_out231_out1            : std_logic;
  SIGNAL Logical_Operator_out232_out1            : std_logic;
  SIGNAL Logical_Operator_out233_out1            : std_logic;
  SIGNAL Logical_Operator_out234_out1            : std_logic;
  SIGNAL Logical_Operator_out235_out1            : std_logic;
  SIGNAL Logical_Operator_out236_out1            : std_logic;
  SIGNAL Logical_Operator_out237_out1            : std_logic;
  SIGNAL Logical_Operator_out238_out1            : std_logic;
  SIGNAL Logical_Operator_out239_out1            : std_logic;
  SIGNAL Logical_Operator_out240_out1            : std_logic;
  SIGNAL Logical_Operator_out241_out1            : std_logic;
  SIGNAL Logical_Operator_out242_out1            : std_logic;
  SIGNAL Logical_Operator_out243_out1            : std_logic;
  SIGNAL Logical_Operator_out244_out1            : std_logic;
  SIGNAL Logical_Operator_out245_out1            : std_logic;
  SIGNAL Logical_Operator_out246_out1            : std_logic;
  SIGNAL Logical_Operator_out247_out1            : std_logic;
  SIGNAL Logical_Operator_out248_out1            : std_logic;
  SIGNAL Logical_Operator_out249_out1            : std_logic;
  SIGNAL Logical_Operator_out250_out1            : std_logic;
  SIGNAL Logical_Operator_out251_out1            : std_logic;
  SIGNAL Logical_Operator_out252_out1            : std_logic;
  SIGNAL Logical_Operator_out253_out1            : std_logic;
  SIGNAL Logical_Operator_out254_out1            : std_logic;
  SIGNAL Logical_Operator_out255_out1            : std_logic;
  SIGNAL Logical_Operator_out256_out1            : std_logic;
  SIGNAL Logical_Operator_out257_out1            : std_logic;
  SIGNAL Logical_Operator_out258_out1            : std_logic;
  SIGNAL Logical_Operator_out259_out1            : std_logic;
  SIGNAL Logical_Operator_out260_out1            : std_logic;
  SIGNAL Logical_Operator_out261_out1            : std_logic;
  SIGNAL Logical_Operator_out262_out1            : std_logic;
  SIGNAL Logical_Operator_out263_out1            : std_logic;
  SIGNAL Logical_Operator_out264_out1            : std_logic;
  SIGNAL Logical_Operator_out265_out1            : std_logic;
  SIGNAL Logical_Operator_out266_out1            : std_logic;
  SIGNAL Logical_Operator_out267_out1            : std_logic;
  SIGNAL Logical_Operator_out268_out1            : std_logic;
  SIGNAL Logical_Operator_out269_out1            : std_logic;
  SIGNAL Logical_Operator_out270_out1            : std_logic;
  SIGNAL Logical_Operator_out271_out1            : std_logic;
  SIGNAL Logical_Operator_out272_out1            : std_logic;
  SIGNAL Logical_Operator_out273_out1            : std_logic;
  SIGNAL Logical_Operator_out274_out1            : std_logic;
  SIGNAL Logical_Operator_out275_out1            : std_logic;
  SIGNAL Logical_Operator_out276_out1            : std_logic;
  SIGNAL Logical_Operator_out277_out1            : std_logic;
  SIGNAL Logical_Operator_out278_out1            : std_logic;
  SIGNAL Logical_Operator_out279_out1            : std_logic;
  SIGNAL Logical_Operator_out280_out1            : std_logic;
  SIGNAL Logical_Operator_out281_out1            : std_logic;
  SIGNAL Logical_Operator_out282_out1            : std_logic;
  SIGNAL Logical_Operator_out283_out1            : std_logic;
  SIGNAL Logical_Operator_out284_out1            : std_logic;
  SIGNAL Logical_Operator_out285_out1            : std_logic;
  SIGNAL Logical_Operator_out286_out1            : std_logic;
  SIGNAL Logical_Operator_out287_out1            : std_logic;
  SIGNAL Logical_Operator_out288_out1            : std_logic;
  SIGNAL Logical_Operator_out289_out1            : std_logic;
  SIGNAL Logical_Operator_out290_out1            : std_logic;
  SIGNAL Logical_Operator_out291_out1            : std_logic;
  SIGNAL Logical_Operator_out292_out1            : std_logic;
  SIGNAL Logical_Operator_out293_out1            : std_logic;
  SIGNAL Logical_Operator_out294_out1            : std_logic;
  SIGNAL Logical_Operator_out295_out1            : std_logic;
  SIGNAL Logical_Operator_out296_out1            : std_logic;
  SIGNAL Logical_Operator_out297_out1            : std_logic;
  SIGNAL Logical_Operator_out298_out1            : std_logic;
  SIGNAL Logical_Operator_out299_out1            : std_logic;
  SIGNAL Logical_Operator_out300_out1            : std_logic;
  SIGNAL Logical_Operator_out301_out1            : std_logic;
  SIGNAL Logical_Operator_out302_out1            : std_logic;
  SIGNAL Logical_Operator_out303_out1            : std_logic;
  SIGNAL Logical_Operator_out304_out1            : std_logic;
  SIGNAL Logical_Operator_out305_out1            : std_logic;
  SIGNAL Logical_Operator_out306_out1            : std_logic;
  SIGNAL Logical_Operator_out307_out1            : std_logic;
  SIGNAL Logical_Operator_out308_out1            : std_logic;
  SIGNAL Logical_Operator_out309_out1            : std_logic;
  SIGNAL Logical_Operator_out310_out1            : std_logic;
  SIGNAL Logical_Operator_out311_out1            : std_logic;
  SIGNAL Logical_Operator_out312_out1            : std_logic;
  SIGNAL Logical_Operator_out313_out1            : std_logic;
  SIGNAL Logical_Operator_out314_out1            : std_logic;
  SIGNAL Logical_Operator_out315_out1            : std_logic;
  SIGNAL Logical_Operator_out316_out1            : std_logic;
  SIGNAL Logical_Operator_out317_out1            : std_logic;
  SIGNAL Logical_Operator_out318_out1            : std_logic;
  SIGNAL Logical_Operator_out319_out1            : std_logic;
  SIGNAL Logical_Operator_out320_out1            : std_logic;
  SIGNAL Logical_Operator_out321_out1            : std_logic;
  SIGNAL Logical_Operator_out322_out1            : std_logic;
  SIGNAL Logical_Operator_out323_out1            : std_logic;
  SIGNAL Logical_Operator_out324_out1            : std_logic;
  SIGNAL Logical_Operator_out325_out1            : std_logic;
  SIGNAL Logical_Operator_out326_out1            : std_logic;
  SIGNAL Logical_Operator_out327_out1            : std_logic;
  SIGNAL Logical_Operator_out328_out1            : std_logic;
  SIGNAL Logical_Operator_out329_out1            : std_logic;
  SIGNAL Logical_Operator_out330_out1            : std_logic;
  SIGNAL Logical_Operator_out331_out1            : std_logic;
  SIGNAL Logical_Operator_out332_out1            : std_logic;
  SIGNAL Logical_Operator_out333_out1            : std_logic;
  SIGNAL Logical_Operator_out334_out1            : std_logic;
  SIGNAL Logical_Operator_out335_out1            : std_logic;
  SIGNAL Logical_Operator_out336_out1            : std_logic;
  SIGNAL Logical_Operator_out337_out1            : std_logic;
  SIGNAL Logical_Operator_out338_out1            : std_logic;
  SIGNAL Logical_Operator_out339_out1            : std_logic;
  SIGNAL Logical_Operator_out340_out1            : std_logic;
  SIGNAL Logical_Operator_out341_out1            : std_logic;
  SIGNAL Logical_Operator_out342_out1            : std_logic;
  SIGNAL Logical_Operator_out343_out1            : std_logic;
  SIGNAL Logical_Operator_out344_out1            : std_logic;
  SIGNAL Logical_Operator_out345_out1            : std_logic;
  SIGNAL Logical_Operator_out346_out1            : std_logic;
  SIGNAL Logical_Operator_out347_out1            : std_logic;
  SIGNAL Logical_Operator_out348_out1            : std_logic;
  SIGNAL Logical_Operator_out349_out1            : std_logic;
  SIGNAL Logical_Operator_out350_out1            : std_logic;
  SIGNAL Logical_Operator_out351_out1            : std_logic;
  SIGNAL Logical_Operator_out352_out1            : std_logic;
  SIGNAL Logical_Operator_out353_out1            : std_logic;
  SIGNAL Logical_Operator_out354_out1            : std_logic;
  SIGNAL Logical_Operator_out355_out1            : std_logic;
  SIGNAL Logical_Operator_out356_out1            : std_logic;
  SIGNAL Logical_Operator_out357_out1            : std_logic;
  SIGNAL Logical_Operator_out358_out1            : std_logic;
  SIGNAL Logical_Operator_out359_out1            : std_logic;
  SIGNAL Logical_Operator_out360_out1            : std_logic;
  SIGNAL Logical_Operator_out361_out1            : std_logic;
  SIGNAL Logical_Operator_out362_out1            : std_logic;
  SIGNAL Logical_Operator_out363_out1            : std_logic;
  SIGNAL Logical_Operator_out364_out1            : std_logic;
  SIGNAL Logical_Operator_out365_out1            : std_logic;
  SIGNAL Logical_Operator_out366_out1            : std_logic;
  SIGNAL Logical_Operator_out367_out1            : std_logic;
  SIGNAL Logical_Operator_out368_out1            : std_logic;
  SIGNAL Logical_Operator_out369_out1            : std_logic;
  SIGNAL Logical_Operator_out370_out1            : std_logic;
  SIGNAL Logical_Operator_out371_out1            : std_logic;
  SIGNAL Logical_Operator_out372_out1            : std_logic;
  SIGNAL Logical_Operator_out373_out1            : std_logic;
  SIGNAL Logical_Operator_out374_out1            : std_logic;
  SIGNAL Logical_Operator_out375_out1            : std_logic;
  SIGNAL Logical_Operator_out376_out1            : std_logic;
  SIGNAL Logical_Operator_out377_out1            : std_logic;
  SIGNAL Logical_Operator_out378_out1            : std_logic;
  SIGNAL Logical_Operator_out379_out1            : std_logic;
  SIGNAL Logical_Operator_out380_out1            : std_logic;
  SIGNAL Logical_Operator_out381_out1            : std_logic;
  SIGNAL Logical_Operator_out382_out1            : std_logic;
  SIGNAL Logical_Operator_out383_out1            : std_logic;
  SIGNAL Logical_Operator_out384_out1            : std_logic;
  SIGNAL Logical_Operator_out385_out1            : std_logic;
  SIGNAL Logical_Operator_out386_out1            : std_logic;
  SIGNAL Logical_Operator_out387_out1            : std_logic;
  SIGNAL Logical_Operator_out388_out1            : std_logic;
  SIGNAL Logical_Operator_out389_out1            : std_logic;
  SIGNAL Logical_Operator_out390_out1            : std_logic;
  SIGNAL Logical_Operator_out391_out1            : std_logic;
  SIGNAL Logical_Operator_out392_out1            : std_logic;
  SIGNAL Logical_Operator_out393_out1            : std_logic;
  SIGNAL Logical_Operator_out394_out1            : std_logic;
  SIGNAL Logical_Operator_out395_out1            : std_logic;
  SIGNAL Logical_Operator_out396_out1            : std_logic;
  SIGNAL Logical_Operator_out397_out1            : std_logic;
  SIGNAL Logical_Operator_out398_out1            : std_logic;
  SIGNAL Logical_Operator_out399_out1            : std_logic;
  SIGNAL Logical_Operator_out400_out1            : std_logic;
  SIGNAL Logical_Operator_out401_out1            : std_logic;
  SIGNAL Logical_Operator_out402_out1            : std_logic;
  SIGNAL Logical_Operator_out403_out1            : std_logic;
  SIGNAL Logical_Operator_out404_out1            : std_logic;
  SIGNAL Logical_Operator_out405_out1            : std_logic;
  SIGNAL Logical_Operator_out406_out1            : std_logic;
  SIGNAL Logical_Operator_out407_out1            : std_logic;
  SIGNAL Logical_Operator_out408_out1            : std_logic;
  SIGNAL Logical_Operator_out409_out1            : std_logic;
  SIGNAL Logical_Operator_out410_out1            : std_logic;
  SIGNAL Logical_Operator_out411_out1            : std_logic;
  SIGNAL Logical_Operator_out412_out1            : std_logic;
  SIGNAL Logical_Operator_out413_out1            : std_logic;
  SIGNAL Logical_Operator_out414_out1            : std_logic;
  SIGNAL Logical_Operator_out415_out1            : std_logic;
  SIGNAL Logical_Operator_out416_out1            : std_logic;
  SIGNAL Logical_Operator_out417_out1            : std_logic;
  SIGNAL Logical_Operator_out418_out1            : std_logic;
  SIGNAL Logical_Operator_out419_out1            : std_logic;
  SIGNAL Logical_Operator_out420_out1            : std_logic;
  SIGNAL Logical_Operator_out421_out1            : std_logic;
  SIGNAL Logical_Operator_out422_out1            : std_logic;
  SIGNAL Logical_Operator_out423_out1            : std_logic;
  SIGNAL Logical_Operator_out424_out1            : std_logic;
  SIGNAL Logical_Operator_out425_out1            : std_logic;
  SIGNAL Logical_Operator_out426_out1            : std_logic;
  SIGNAL Logical_Operator_out427_out1            : std_logic;
  SIGNAL Logical_Operator_out428_out1            : std_logic;
  SIGNAL Logical_Operator_out429_out1            : std_logic;
  SIGNAL Logical_Operator_out430_out1            : std_logic;
  SIGNAL Logical_Operator_out431_out1            : std_logic;
  SIGNAL Logical_Operator_out432_out1            : std_logic;
  SIGNAL Logical_Operator_out433_out1            : std_logic;
  SIGNAL Logical_Operator_out434_out1            : std_logic;
  SIGNAL Logical_Operator_out435_out1            : std_logic;
  SIGNAL Logical_Operator_out436_out1            : std_logic;
  SIGNAL Logical_Operator_out437_out1            : std_logic;
  SIGNAL Logical_Operator_out438_out1            : std_logic;
  SIGNAL Logical_Operator_out439_out1            : std_logic;
  SIGNAL Logical_Operator_out440_out1            : std_logic;
  SIGNAL Logical_Operator_out441_out1            : std_logic;
  SIGNAL Logical_Operator_out442_out1            : std_logic;
  SIGNAL Logical_Operator_out443_out1            : std_logic;
  SIGNAL Logical_Operator_out444_out1            : std_logic;
  SIGNAL Logical_Operator_out445_out1            : std_logic;
  SIGNAL Logical_Operator_out446_out1            : std_logic;
  SIGNAL Logical_Operator_out447_out1            : std_logic;
  SIGNAL Logical_Operator_out448_out1            : std_logic;
  SIGNAL Logical_Operator_out449_out1            : std_logic;
  SIGNAL Logical_Operator_out450_out1            : std_logic;
  SIGNAL Logical_Operator_out451_out1            : std_logic;
  SIGNAL Logical_Operator_out452_out1            : std_logic;
  SIGNAL Logical_Operator_out453_out1            : std_logic;
  SIGNAL Logical_Operator_out454_out1            : std_logic;
  SIGNAL Logical_Operator_out455_out1            : std_logic;
  SIGNAL Logical_Operator_out456_out1            : std_logic;
  SIGNAL Logical_Operator_out457_out1            : std_logic;
  SIGNAL Logical_Operator_out458_out1            : std_logic;
  SIGNAL Logical_Operator_out459_out1            : std_logic;
  SIGNAL Logical_Operator_out460_out1            : std_logic;
  SIGNAL Logical_Operator_out461_out1            : std_logic;
  SIGNAL Logical_Operator_out462_out1            : std_logic;
  SIGNAL Logical_Operator_out463_out1            : std_logic;
  SIGNAL Logical_Operator_out464_out1            : std_logic;
  SIGNAL Logical_Operator_out465_out1            : std_logic;
  SIGNAL Logical_Operator_out466_out1            : std_logic;
  SIGNAL Logical_Operator_out467_out1            : std_logic;
  SIGNAL Logical_Operator_out468_out1            : std_logic;
  SIGNAL Logical_Operator_out469_out1            : std_logic;
  SIGNAL Logical_Operator_out470_out1            : std_logic;
  SIGNAL Logical_Operator_out471_out1            : std_logic;
  SIGNAL Logical_Operator_out472_out1            : std_logic;
  SIGNAL Logical_Operator_out473_out1            : std_logic;
  SIGNAL Logical_Operator_out474_out1            : std_logic;
  SIGNAL Logical_Operator_out475_out1            : std_logic;
  SIGNAL Logical_Operator_out476_out1            : std_logic;
  SIGNAL Logical_Operator_out477_out1            : std_logic;
  SIGNAL Logical_Operator_out478_out1            : std_logic;
  SIGNAL Logical_Operator_out479_out1            : std_logic;
  SIGNAL Logical_Operator_out480_out1            : std_logic;
  SIGNAL Logical_Operator_out481_out1            : std_logic;
  SIGNAL Logical_Operator_out482_out1            : std_logic;
  SIGNAL Logical_Operator_out483_out1            : std_logic;
  SIGNAL Logical_Operator_out484_out1            : std_logic;
  SIGNAL Logical_Operator_out485_out1            : std_logic;
  SIGNAL Logical_Operator_out486_out1            : std_logic;
  SIGNAL Logical_Operator_out487_out1            : std_logic;
  SIGNAL Logical_Operator_out488_out1            : std_logic;
  SIGNAL Logical_Operator_out489_out1            : std_logic;
  SIGNAL Logical_Operator_out490_out1            : std_logic;
  SIGNAL Logical_Operator_out491_out1            : std_logic;
  SIGNAL Logical_Operator_out492_out1            : std_logic;
  SIGNAL Logical_Operator_out493_out1            : std_logic;
  SIGNAL Logical_Operator_out494_out1            : std_logic;
  SIGNAL Logical_Operator_out495_out1            : std_logic;
  SIGNAL Logical_Operator_out496_out1            : std_logic;
  SIGNAL Logical_Operator_out497_out1            : std_logic;
  SIGNAL Logical_Operator_out498_out1            : std_logic;
  SIGNAL Logical_Operator_out499_out1            : std_logic;
  SIGNAL Logical_Operator_out500_out1            : std_logic;
  SIGNAL Logical_Operator_out501_out1            : std_logic;
  SIGNAL Logical_Operator_out502_out1            : std_logic;
  SIGNAL Logical_Operator_out503_out1            : std_logic;
  SIGNAL Logical_Operator_out504_out1            : std_logic;
  SIGNAL Logical_Operator_out505_out1            : std_logic;
  SIGNAL Logical_Operator_out506_out1            : std_logic;
  SIGNAL Logical_Operator_out507_out1            : std_logic;
  SIGNAL Logical_Operator_out508_out1            : std_logic;
  SIGNAL Logical_Operator_out509_out1            : std_logic;
  SIGNAL Logical_Operator_out510_out1            : std_logic;
  SIGNAL Logical_Operator_out511_out1            : std_logic;
  SIGNAL Logical_Operator_out512_out1            : std_logic;
  SIGNAL Logical_Operator_out513_out1            : std_logic;
  SIGNAL Logical_Operator_out514_out1            : std_logic;
  SIGNAL Logical_Operator_out515_out1            : std_logic;
  SIGNAL Logical_Operator_out516_out1            : std_logic;
  SIGNAL Logical_Operator_out517_out1            : std_logic;
  SIGNAL Logical_Operator_out518_out1            : std_logic;
  SIGNAL Logical_Operator_out519_out1            : std_logic;
  SIGNAL Logical_Operator_out520_out1            : std_logic;
  SIGNAL Logical_Operator_out521_out1            : std_logic;
  SIGNAL Logical_Operator_out522_out1            : std_logic;
  SIGNAL Logical_Operator_out523_out1            : std_logic;
  SIGNAL Logical_Operator_out524_out1            : std_logic;
  SIGNAL Logical_Operator_out525_out1            : std_logic;
  SIGNAL Logical_Operator_out526_out1            : std_logic;
  SIGNAL Logical_Operator_out527_out1            : std_logic;
  SIGNAL Logical_Operator_out528_out1            : std_logic;
  SIGNAL Logical_Operator_out529_out1            : std_logic;
  SIGNAL Logical_Operator_out530_out1            : std_logic;
  SIGNAL Logical_Operator_out531_out1            : std_logic;
  SIGNAL Logical_Operator_out532_out1            : std_logic;
  SIGNAL Logical_Operator_out533_out1            : std_logic;
  SIGNAL Logical_Operator_out534_out1            : std_logic;
  SIGNAL Logical_Operator_out535_out1            : std_logic;
  SIGNAL Logical_Operator_out536_out1            : std_logic;
  SIGNAL Logical_Operator_out537_out1            : std_logic;
  SIGNAL Logical_Operator_out538_out1            : std_logic;
  SIGNAL Logical_Operator_out539_out1            : std_logic;
  SIGNAL Logical_Operator_out540_out1            : std_logic;
  SIGNAL Logical_Operator_out541_out1            : std_logic;
  SIGNAL Logical_Operator_out542_out1            : std_logic;
  SIGNAL Logical_Operator_out543_out1            : std_logic;
  SIGNAL Logical_Operator_out544_out1            : std_logic;
  SIGNAL Logical_Operator_out545_out1            : std_logic;
  SIGNAL Logical_Operator_out546_out1            : std_logic;
  SIGNAL Logical_Operator_out547_out1            : std_logic;
  SIGNAL Logical_Operator_out548_out1            : std_logic;
  SIGNAL Logical_Operator_out549_out1            : std_logic;
  SIGNAL Logical_Operator_out550_out1            : std_logic;
  SIGNAL Logical_Operator_out551_out1            : std_logic;
  SIGNAL Logical_Operator_out552_out1            : std_logic;
  SIGNAL Logical_Operator_out553_out1            : std_logic;
  SIGNAL Logical_Operator_out554_out1            : std_logic;
  SIGNAL Logical_Operator_out555_out1            : std_logic;
  SIGNAL Logical_Operator_out556_out1            : std_logic;
  SIGNAL Logical_Operator_out557_out1            : std_logic;
  SIGNAL Logical_Operator_out558_out1            : std_logic;
  SIGNAL Logical_Operator_out559_out1            : std_logic;
  SIGNAL Logical_Operator_out560_out1            : std_logic;
  SIGNAL Logical_Operator_out561_out1            : std_logic;
  SIGNAL Logical_Operator_out562_out1            : std_logic;
  SIGNAL Logical_Operator_out563_out1            : std_logic;
  SIGNAL Logical_Operator_out564_out1            : std_logic;
  SIGNAL Logical_Operator_out565_out1            : std_logic;
  SIGNAL Logical_Operator_out566_out1            : std_logic;
  SIGNAL Logical_Operator_out567_out1            : std_logic;
  SIGNAL Logical_Operator_out568_out1            : std_logic;
  SIGNAL Logical_Operator_out569_out1            : std_logic;
  SIGNAL Logical_Operator_out570_out1            : std_logic;
  SIGNAL Logical_Operator_out571_out1            : std_logic;
  SIGNAL Logical_Operator_out572_out1            : std_logic;
  SIGNAL Logical_Operator_out573_out1            : std_logic;
  SIGNAL Logical_Operator_out574_out1            : std_logic;
  SIGNAL Logical_Operator_out575_out1            : std_logic;
  SIGNAL Logical_Operator_out576_out1            : std_logic;
  SIGNAL Logical_Operator_out577_out1            : std_logic;
  SIGNAL Logical_Operator_out578_out1            : std_logic;
  SIGNAL Logical_Operator_out579_out1            : std_logic;
  SIGNAL Logical_Operator_out580_out1            : std_logic;
  SIGNAL Logical_Operator_out581_out1            : std_logic;
  SIGNAL Logical_Operator_out582_out1            : std_logic;
  SIGNAL Logical_Operator_out583_out1            : std_logic;
  SIGNAL Logical_Operator_out584_out1            : std_logic;
  SIGNAL Logical_Operator_out585_out1            : std_logic;
  SIGNAL Logical_Operator_out586_out1            : std_logic;
  SIGNAL Logical_Operator_out587_out1            : std_logic;
  SIGNAL Logical_Operator_out588_out1            : std_logic;
  SIGNAL Logical_Operator_out589_out1            : std_logic;
  SIGNAL Logical_Operator_out590_out1            : std_logic;
  SIGNAL Logical_Operator_out591_out1            : std_logic;
  SIGNAL Logical_Operator_out592_out1            : std_logic;
  SIGNAL Logical_Operator_out593_out1            : std_logic;
  SIGNAL Logical_Operator_out594_out1            : std_logic;
  SIGNAL Logical_Operator_out595_out1            : std_logic;
  SIGNAL Logical_Operator_out596_out1            : std_logic;
  SIGNAL Logical_Operator_out597_out1            : std_logic;
  SIGNAL Logical_Operator_out598_out1            : std_logic;
  SIGNAL Logical_Operator_out599_out1            : std_logic;
  SIGNAL Logical_Operator_out600_out1            : std_logic;
  SIGNAL Logical_Operator_out601_out1            : std_logic;
  SIGNAL Logical_Operator_out602_out1            : std_logic;
  SIGNAL Logical_Operator_out603_out1            : std_logic;
  SIGNAL Logical_Operator_out604_out1            : std_logic;
  SIGNAL Logical_Operator_out605_out1            : std_logic;
  SIGNAL Logical_Operator_out606_out1            : std_logic;
  SIGNAL Logical_Operator_out607_out1            : std_logic;
  SIGNAL Logical_Operator_out608_out1            : std_logic;
  SIGNAL Logical_Operator_out609_out1            : std_logic;
  SIGNAL Logical_Operator_out610_out1            : std_logic;
  SIGNAL Logical_Operator_out611_out1            : std_logic;
  SIGNAL Logical_Operator_out612_out1            : std_logic;
  SIGNAL Logical_Operator_out613_out1            : std_logic;
  SIGNAL Logical_Operator_out614_out1            : std_logic;
  SIGNAL Logical_Operator_out615_out1            : std_logic;
  SIGNAL Logical_Operator_out616_out1            : std_logic;
  SIGNAL Logical_Operator_out617_out1            : std_logic;
  SIGNAL Logical_Operator_out618_out1            : std_logic;
  SIGNAL Logical_Operator_out619_out1            : std_logic;
  SIGNAL Logical_Operator_out620_out1            : std_logic;
  SIGNAL Logical_Operator_out621_out1            : std_logic;
  SIGNAL Logical_Operator_out622_out1            : std_logic;
  SIGNAL Logical_Operator_out623_out1            : std_logic;
  SIGNAL Logical_Operator_out624_out1            : std_logic;
  SIGNAL Logical_Operator_out625_out1            : std_logic;
  SIGNAL Logical_Operator_out626_out1            : std_logic;
  SIGNAL Logical_Operator_out627_out1            : std_logic;
  SIGNAL Logical_Operator_out628_out1            : std_logic;
  SIGNAL Logical_Operator_out629_out1            : std_logic;
  SIGNAL Logical_Operator_out630_out1            : std_logic;
  SIGNAL Logical_Operator_out631_out1            : std_logic;
  SIGNAL Logical_Operator_out632_out1            : std_logic;
  SIGNAL Logical_Operator_out633_out1            : std_logic;
  SIGNAL Logical_Operator_out634_out1            : std_logic;
  SIGNAL Logical_Operator_out635_out1            : std_logic;
  SIGNAL Logical_Operator_out636_out1            : std_logic;
  SIGNAL Logical_Operator_out637_out1            : std_logic;
  SIGNAL Logical_Operator_out638_out1            : std_logic;
  SIGNAL Logical_Operator_out639_out1            : std_logic;
  SIGNAL Logical_Operator_out640_out1            : std_logic;
  SIGNAL Logical_Operator_out641_out1            : std_logic;
  SIGNAL Logical_Operator_out642_out1            : std_logic;
  SIGNAL Logical_Operator_out643_out1            : std_logic;
  SIGNAL Logical_Operator_out644_out1            : std_logic;
  SIGNAL Logical_Operator_out645_out1            : std_logic;
  SIGNAL Logical_Operator_out646_out1            : std_logic;
  SIGNAL Logical_Operator_out647_out1            : std_logic;
  SIGNAL Logical_Operator_out648_out1            : std_logic;
  SIGNAL Logical_Operator_out649_out1            : std_logic;
  SIGNAL Logical_Operator_out650_out1            : std_logic;
  SIGNAL Logical_Operator_out651_out1            : std_logic;
  SIGNAL Logical_Operator_out652_out1            : std_logic;
  SIGNAL Logical_Operator_out653_out1            : std_logic;
  SIGNAL Logical_Operator_out654_out1            : std_logic;
  SIGNAL Logical_Operator_out655_out1            : std_logic;
  SIGNAL Logical_Operator_out656_out1            : std_logic;
  SIGNAL Logical_Operator_out657_out1            : std_logic;
  SIGNAL Logical_Operator_out658_out1            : std_logic;
  SIGNAL Logical_Operator_out659_out1            : std_logic;
  SIGNAL Logical_Operator_out660_out1            : std_logic;
  SIGNAL Logical_Operator_out661_out1            : std_logic;
  SIGNAL Logical_Operator_out662_out1            : std_logic;
  SIGNAL Logical_Operator_out663_out1            : std_logic;
  SIGNAL Logical_Operator_out664_out1            : std_logic;
  SIGNAL Logical_Operator_out665_out1            : std_logic;
  SIGNAL Logical_Operator_out666_out1            : std_logic;
  SIGNAL Logical_Operator_out667_out1            : std_logic;
  SIGNAL Logical_Operator_out668_out1            : std_logic;
  SIGNAL Logical_Operator_out669_out1            : std_logic;
  SIGNAL Logical_Operator_out670_out1            : std_logic;
  SIGNAL Logical_Operator_out671_out1            : std_logic;
  SIGNAL Logical_Operator_out672_out1            : std_logic;
  SIGNAL Logical_Operator_out673_out1            : std_logic;
  SIGNAL Logical_Operator_out674_out1            : std_logic;
  SIGNAL Logical_Operator_out675_out1            : std_logic;
  SIGNAL Logical_Operator_out676_out1            : std_logic;
  SIGNAL Logical_Operator_out677_out1            : std_logic;
  SIGNAL Logical_Operator_out678_out1            : std_logic;
  SIGNAL Logical_Operator_out679_out1            : std_logic;
  SIGNAL Logical_Operator_out680_out1            : std_logic;
  SIGNAL Logical_Operator_out681_out1            : std_logic;
  SIGNAL Logical_Operator_out682_out1            : std_logic;
  SIGNAL Logical_Operator_out683_out1            : std_logic;
  SIGNAL Logical_Operator_out684_out1            : std_logic;
  SIGNAL Logical_Operator_out685_out1            : std_logic;
  SIGNAL Logical_Operator_out686_out1            : std_logic;
  SIGNAL Logical_Operator_out687_out1            : std_logic;
  SIGNAL Logical_Operator_out688_out1            : std_logic;
  SIGNAL Logical_Operator_out689_out1            : std_logic;
  SIGNAL Logical_Operator_out690_out1            : std_logic;
  SIGNAL Logical_Operator_out691_out1            : std_logic;
  SIGNAL Logical_Operator_out692_out1            : std_logic;
  SIGNAL Logical_Operator_out693_out1            : std_logic;
  SIGNAL Logical_Operator_out694_out1            : std_logic;
  SIGNAL Logical_Operator_out695_out1            : std_logic;
  SIGNAL Logical_Operator_out696_out1            : std_logic;
  SIGNAL Logical_Operator_out697_out1            : std_logic;
  SIGNAL Logical_Operator_out698_out1            : std_logic;
  SIGNAL Logical_Operator_out699_out1            : std_logic;
  SIGNAL Logical_Operator_out700_out1            : std_logic;
  SIGNAL Logical_Operator_out701_out1            : std_logic;
  SIGNAL Logical_Operator_out702_out1            : std_logic;
  SIGNAL Logical_Operator_out703_out1            : std_logic;
  SIGNAL Logical_Operator_out704_out1            : std_logic;
  SIGNAL Logical_Operator_out705_out1            : std_logic;
  SIGNAL Logical_Operator_out706_out1            : std_logic;
  SIGNAL Logical_Operator_out707_out1            : std_logic;
  SIGNAL Logical_Operator_out708_out1            : std_logic;
  SIGNAL Logical_Operator_out709_out1            : std_logic;
  SIGNAL Logical_Operator_out710_out1            : std_logic;
  SIGNAL Logical_Operator_out711_out1            : std_logic;
  SIGNAL Logical_Operator_out712_out1            : std_logic;
  SIGNAL Logical_Operator_out713_out1            : std_logic;
  SIGNAL Logical_Operator_out714_out1            : std_logic;
  SIGNAL Logical_Operator_out715_out1            : std_logic;
  SIGNAL Logical_Operator_out716_out1            : std_logic;
  SIGNAL Logical_Operator_out717_out1            : std_logic;
  SIGNAL Logical_Operator_out718_out1            : std_logic;
  SIGNAL Logical_Operator_out719_out1            : std_logic;
  SIGNAL Logical_Operator_out720_out1            : std_logic;
  SIGNAL Logical_Operator_out721_out1            : std_logic;
  SIGNAL Logical_Operator_out722_out1            : std_logic;
  SIGNAL Logical_Operator_out723_out1            : std_logic;
  SIGNAL Logical_Operator_out724_out1            : std_logic;
  SIGNAL Logical_Operator_out725_out1            : std_logic;
  SIGNAL Logical_Operator_out726_out1            : std_logic;
  SIGNAL Logical_Operator_out727_out1            : std_logic;
  SIGNAL Logical_Operator_out728_out1            : std_logic;
  SIGNAL Logical_Operator_out729_out1            : std_logic;
  SIGNAL Logical_Operator_out730_out1            : std_logic;
  SIGNAL Logical_Operator_out731_out1            : std_logic;
  SIGNAL Logical_Operator_out732_out1            : std_logic;
  SIGNAL Logical_Operator_out733_out1            : std_logic;
  SIGNAL Logical_Operator_out734_out1            : std_logic;
  SIGNAL Logical_Operator_out735_out1            : std_logic;
  SIGNAL Logical_Operator_out736_out1            : std_logic;
  SIGNAL Logical_Operator_out737_out1            : std_logic;
  SIGNAL Logical_Operator_out738_out1            : std_logic;
  SIGNAL Logical_Operator_out739_out1            : std_logic;
  SIGNAL Logical_Operator_out740_out1            : std_logic;
  SIGNAL Logical_Operator_out741_out1            : std_logic;
  SIGNAL Logical_Operator_out742_out1            : std_logic;
  SIGNAL Logical_Operator_out743_out1            : std_logic;
  SIGNAL Logical_Operator_out744_out1            : std_logic;
  SIGNAL Logical_Operator_out745_out1            : std_logic;
  SIGNAL Logical_Operator_out746_out1            : std_logic;
  SIGNAL Logical_Operator_out747_out1            : std_logic;
  SIGNAL Logical_Operator_out748_out1            : std_logic;
  SIGNAL Logical_Operator_out749_out1            : std_logic;
  SIGNAL Logical_Operator_out750_out1            : std_logic;
  SIGNAL Logical_Operator_out751_out1            : std_logic;
  SIGNAL Logical_Operator_out752_out1            : std_logic;
  SIGNAL Logical_Operator_out753_out1            : std_logic;
  SIGNAL Logical_Operator_out754_out1            : std_logic;
  SIGNAL Logical_Operator_out755_out1            : std_logic;
  SIGNAL Logical_Operator_out756_out1            : std_logic;
  SIGNAL Logical_Operator_out757_out1            : std_logic;
  SIGNAL Logical_Operator_out758_out1            : std_logic;
  SIGNAL Logical_Operator_out759_out1            : std_logic;
  SIGNAL Logical_Operator_out760_out1            : std_logic;
  SIGNAL Logical_Operator_out761_out1            : std_logic;
  SIGNAL Logical_Operator_out762_out1            : std_logic;
  SIGNAL Logical_Operator_out763_out1            : std_logic;
  SIGNAL Logical_Operator_out764_out1            : std_logic;
  SIGNAL Logical_Operator_out765_out1            : std_logic;
  SIGNAL Logical_Operator_out766_out1            : std_logic;
  SIGNAL Logical_Operator_out767_out1            : std_logic;
  SIGNAL Logical_Operator_out768_out1            : std_logic;
  SIGNAL Logical_Operator_out769_out1            : std_logic;
  SIGNAL Logical_Operator_out770_out1            : std_logic;
  SIGNAL Logical_Operator_out771_out1            : std_logic;
  SIGNAL Logical_Operator_out772_out1            : std_logic;
  SIGNAL Logical_Operator_out773_out1            : std_logic;
  SIGNAL Logical_Operator_out774_out1            : std_logic;
  SIGNAL Logical_Operator_out775_out1            : std_logic;
  SIGNAL Logical_Operator_out776_out1            : std_logic;
  SIGNAL Logical_Operator_out777_out1            : std_logic;
  SIGNAL Logical_Operator_out778_out1            : std_logic;
  SIGNAL Logical_Operator_out779_out1            : std_logic;
  SIGNAL Logical_Operator_out780_out1            : std_logic;
  SIGNAL Logical_Operator_out781_out1            : std_logic;
  SIGNAL Logical_Operator_out782_out1            : std_logic;
  SIGNAL Logical_Operator_out783_out1            : std_logic;
  SIGNAL Logical_Operator_out784_out1            : std_logic;
  SIGNAL Logical_Operator_out785_out1            : std_logic;
  SIGNAL Logical_Operator_out786_out1            : std_logic;
  SIGNAL Logical_Operator_out787_out1            : std_logic;
  SIGNAL Logical_Operator_out788_out1            : std_logic;
  SIGNAL Logical_Operator_out789_out1            : std_logic;
  SIGNAL Logical_Operator_out790_out1            : std_logic;
  SIGNAL Logical_Operator_out791_out1            : std_logic;
  SIGNAL Logical_Operator_out792_out1            : std_logic;
  SIGNAL Logical_Operator_out793_out1            : std_logic;
  SIGNAL Logical_Operator_out794_out1            : std_logic;
  SIGNAL Logical_Operator_out795_out1            : std_logic;
  SIGNAL Logical_Operator_out796_out1            : std_logic;
  SIGNAL Logical_Operator_out797_out1            : std_logic;
  SIGNAL Logical_Operator_out798_out1            : std_logic;
  SIGNAL Logical_Operator_out799_out1            : std_logic;
  SIGNAL Logical_Operator_out800_out1            : std_logic;
  SIGNAL Logical_Operator_out801_out1            : std_logic;
  SIGNAL Logical_Operator_out802_out1            : std_logic;
  SIGNAL Logical_Operator_out803_out1            : std_logic;
  SIGNAL Logical_Operator_out804_out1            : std_logic;
  SIGNAL Logical_Operator_out805_out1            : std_logic;
  SIGNAL Logical_Operator_out806_out1            : std_logic;
  SIGNAL Logical_Operator_out807_out1            : std_logic;
  SIGNAL Logical_Operator_out808_out1            : std_logic;
  SIGNAL Logical_Operator_out809_out1            : std_logic;
  SIGNAL Logical_Operator_out810_out1            : std_logic;
  SIGNAL Logical_Operator_out811_out1            : std_logic;
  SIGNAL Logical_Operator_out812_out1            : std_logic;
  SIGNAL Logical_Operator_out813_out1            : std_logic;
  SIGNAL Logical_Operator_out814_out1            : std_logic;
  SIGNAL Logical_Operator_out815_out1            : std_logic;
  SIGNAL Logical_Operator_out816_out1            : std_logic;
  SIGNAL Logical_Operator_out817_out1            : std_logic;
  SIGNAL Logical_Operator_out818_out1            : std_logic;
  SIGNAL Logical_Operator_out819_out1            : std_logic;
  SIGNAL Logical_Operator_out820_out1            : std_logic;
  SIGNAL Logical_Operator_out821_out1            : std_logic;
  SIGNAL Logical_Operator_out822_out1            : std_logic;
  SIGNAL Logical_Operator_out823_out1            : std_logic;
  SIGNAL Logical_Operator_out824_out1            : std_logic;
  SIGNAL Logical_Operator_out825_out1            : std_logic;
  SIGNAL Logical_Operator_out826_out1            : std_logic;
  SIGNAL Logical_Operator_out827_out1            : std_logic;
  SIGNAL Logical_Operator_out828_out1            : std_logic;
  SIGNAL Logical_Operator_out829_out1            : std_logic;
  SIGNAL Logical_Operator_out830_out1            : std_logic;
  SIGNAL Logical_Operator_out831_out1            : std_logic;
  SIGNAL Logical_Operator_out832_out1            : std_logic;
  SIGNAL Logical_Operator_out833_out1            : std_logic;
  SIGNAL Logical_Operator_out834_out1            : std_logic;
  SIGNAL Logical_Operator_out835_out1            : std_logic;
  SIGNAL Logical_Operator_out836_out1            : std_logic;
  SIGNAL Logical_Operator_out837_out1            : std_logic;
  SIGNAL Logical_Operator_out838_out1            : std_logic;
  SIGNAL Logical_Operator_out839_out1            : std_logic;
  SIGNAL Logical_Operator_out840_out1            : std_logic;
  SIGNAL Logical_Operator_out841_out1            : std_logic;
  SIGNAL Logical_Operator_out842_out1            : std_logic;
  SIGNAL Logical_Operator_out843_out1            : std_logic;
  SIGNAL Logical_Operator_out844_out1            : std_logic;
  SIGNAL Logical_Operator_out845_out1            : std_logic;
  SIGNAL Logical_Operator_out846_out1            : std_logic;
  SIGNAL Logical_Operator_out847_out1            : std_logic;
  SIGNAL Logical_Operator_out848_out1            : std_logic;
  SIGNAL Logical_Operator_out849_out1            : std_logic;
  SIGNAL Logical_Operator_out850_out1            : std_logic;
  SIGNAL Logical_Operator_out851_out1            : std_logic;
  SIGNAL Logical_Operator_out852_out1            : std_logic;
  SIGNAL Logical_Operator_out853_out1            : std_logic;
  SIGNAL Logical_Operator_out854_out1            : std_logic;
  SIGNAL Logical_Operator_out855_out1            : std_logic;
  SIGNAL Logical_Operator_out856_out1            : std_logic;
  SIGNAL Logical_Operator_out857_out1            : std_logic;
  SIGNAL Logical_Operator_out858_out1            : std_logic;
  SIGNAL Logical_Operator_out859_out1            : std_logic;
  SIGNAL Logical_Operator_out860_out1            : std_logic;
  SIGNAL Logical_Operator_out861_out1            : std_logic;
  SIGNAL Logical_Operator_out862_out1            : std_logic;
  SIGNAL Logical_Operator_out863_out1            : std_logic;
  SIGNAL Logical_Operator_out864_out1            : std_logic;
  SIGNAL Logical_Operator_out865_out1            : std_logic;
  SIGNAL Logical_Operator_out866_out1            : std_logic;
  SIGNAL Logical_Operator_out867_out1            : std_logic;
  SIGNAL Logical_Operator_out868_out1            : std_logic;
  SIGNAL Logical_Operator_out869_out1            : std_logic;
  SIGNAL Logical_Operator_out870_out1            : std_logic;
  SIGNAL Logical_Operator_out871_out1            : std_logic;
  SIGNAL Logical_Operator_out872_out1            : std_logic;
  SIGNAL Logical_Operator_out873_out1            : std_logic;
  SIGNAL Logical_Operator_out874_out1            : std_logic;
  SIGNAL Logical_Operator_out875_out1            : std_logic;
  SIGNAL Logical_Operator_out876_out1            : std_logic;
  SIGNAL Logical_Operator_out877_out1            : std_logic;
  SIGNAL Logical_Operator_out878_out1            : std_logic;
  SIGNAL Logical_Operator_out879_out1            : std_logic;
  SIGNAL Logical_Operator_out880_out1            : std_logic;
  SIGNAL Logical_Operator_out881_out1            : std_logic;
  SIGNAL Logical_Operator_out882_out1            : std_logic;
  SIGNAL Logical_Operator_out883_out1            : std_logic;
  SIGNAL Logical_Operator_out884_out1            : std_logic;
  SIGNAL Logical_Operator_out885_out1            : std_logic;
  SIGNAL Logical_Operator_out886_out1            : std_logic;
  SIGNAL Logical_Operator_out887_out1            : std_logic;
  SIGNAL Logical_Operator_out888_out1            : std_logic;
  SIGNAL Logical_Operator_out889_out1            : std_logic;
  SIGNAL Logical_Operator_out890_out1            : std_logic;
  SIGNAL Logical_Operator_out891_out1            : std_logic;
  SIGNAL Logical_Operator_out892_out1            : std_logic;
  SIGNAL Logical_Operator_out893_out1            : std_logic;
  SIGNAL Logical_Operator_out894_out1            : std_logic;
  SIGNAL Logical_Operator_out895_out1            : std_logic;
  SIGNAL Logical_Operator_out896_out1            : std_logic;
  SIGNAL Logical_Operator_out897_out1            : std_logic;
  SIGNAL Logical_Operator_out898_out1            : std_logic;
  SIGNAL Logical_Operator_out899_out1            : std_logic;
  SIGNAL Logical_Operator_out900_out1            : std_logic;
  SIGNAL Logical_Operator_out901_out1            : std_logic;
  SIGNAL Logical_Operator_out902_out1            : std_logic;
  SIGNAL Logical_Operator_out903_out1            : std_logic;
  SIGNAL Logical_Operator_out904_out1            : std_logic;
  SIGNAL Logical_Operator_out905_out1            : std_logic;
  SIGNAL Logical_Operator_out906_out1            : std_logic;
  SIGNAL Logical_Operator_out907_out1            : std_logic;
  SIGNAL Logical_Operator_out908_out1            : std_logic;
  SIGNAL Logical_Operator_out909_out1            : std_logic;
  SIGNAL Logical_Operator_out910_out1            : std_logic;
  SIGNAL Logical_Operator_out911_out1            : std_logic;
  SIGNAL Logical_Operator_out912_out1            : std_logic;
  SIGNAL Logical_Operator_out913_out1            : std_logic;
  SIGNAL Logical_Operator_out914_out1            : std_logic;
  SIGNAL Logical_Operator_out915_out1            : std_logic;
  SIGNAL Logical_Operator_out916_out1            : std_logic;
  SIGNAL Logical_Operator_out917_out1            : std_logic;
  SIGNAL Logical_Operator_out918_out1            : std_logic;
  SIGNAL Logical_Operator_out919_out1            : std_logic;
  SIGNAL Logical_Operator_out920_out1            : std_logic;
  SIGNAL Logical_Operator_out921_out1            : std_logic;
  SIGNAL Logical_Operator_out922_out1            : std_logic;
  SIGNAL Logical_Operator_out923_out1            : std_logic;
  SIGNAL Logical_Operator_out924_out1            : std_logic;
  SIGNAL Logical_Operator_out925_out1            : std_logic;
  SIGNAL Logical_Operator_out926_out1            : std_logic;
  SIGNAL Logical_Operator_out927_out1            : std_logic;
  SIGNAL Logical_Operator_out928_out1            : std_logic;
  SIGNAL Logical_Operator_out929_out1            : std_logic;
  SIGNAL Logical_Operator_out930_out1            : std_logic;
  SIGNAL Logical_Operator_out931_out1            : std_logic;
  SIGNAL Logical_Operator_out932_out1            : std_logic;
  SIGNAL Logical_Operator_out933_out1            : std_logic;
  SIGNAL Logical_Operator_out934_out1            : std_logic;
  SIGNAL Logical_Operator_out935_out1            : std_logic;
  SIGNAL Logical_Operator_out936_out1            : std_logic;
  SIGNAL Logical_Operator_out937_out1            : std_logic;
  SIGNAL Logical_Operator_out938_out1            : std_logic;
  SIGNAL Logical_Operator_out939_out1            : std_logic;
  SIGNAL Logical_Operator_out940_out1            : std_logic;
  SIGNAL Logical_Operator_out941_out1            : std_logic;
  SIGNAL Logical_Operator_out942_out1            : std_logic;
  SIGNAL Logical_Operator_out943_out1            : std_logic;
  SIGNAL Logical_Operator_out944_out1            : std_logic;
  SIGNAL Logical_Operator_out945_out1            : std_logic;
  SIGNAL Logical_Operator_out946_out1            : std_logic;
  SIGNAL Logical_Operator_out947_out1            : std_logic;
  SIGNAL Logical_Operator_out948_out1            : std_logic;
  SIGNAL Logical_Operator_out949_out1            : std_logic;
  SIGNAL Logical_Operator_out950_out1            : std_logic;
  SIGNAL Logical_Operator_out951_out1            : std_logic;
  SIGNAL Logical_Operator_out952_out1            : std_logic;
  SIGNAL Logical_Operator_out953_out1            : std_logic;
  SIGNAL Logical_Operator_out954_out1            : std_logic;
  SIGNAL Logical_Operator_out955_out1            : std_logic;
  SIGNAL Logical_Operator_out956_out1            : std_logic;
  SIGNAL Logical_Operator_out957_out1            : std_logic;
  SIGNAL Logical_Operator_out958_out1            : std_logic;
  SIGNAL Logical_Operator_out959_out1            : std_logic;
  SIGNAL Logical_Operator_out960_out1            : std_logic;
  SIGNAL Logical_Operator_out961_out1            : std_logic;
  SIGNAL Logical_Operator_out962_out1            : std_logic;
  SIGNAL Logical_Operator_out963_out1            : std_logic;
  SIGNAL Logical_Operator_out964_out1            : std_logic;
  SIGNAL Logical_Operator_out965_out1            : std_logic;
  SIGNAL Logical_Operator_out966_out1            : std_logic;
  SIGNAL Logical_Operator_out967_out1            : std_logic;
  SIGNAL Logical_Operator_out968_out1            : std_logic;
  SIGNAL Logical_Operator_out969_out1            : std_logic;
  SIGNAL Logical_Operator_out970_out1            : std_logic;
  SIGNAL Logical_Operator_out971_out1            : std_logic;
  SIGNAL Logical_Operator_out972_out1            : std_logic;
  SIGNAL Logical_Operator_out973_out1            : std_logic;
  SIGNAL Logical_Operator_out974_out1            : std_logic;
  SIGNAL Logical_Operator_out975_out1            : std_logic;
  SIGNAL Logical_Operator_out976_out1            : std_logic;
  SIGNAL Logical_Operator_out977_out1            : std_logic;
  SIGNAL Logical_Operator_out978_out1            : std_logic;
  SIGNAL Logical_Operator_out979_out1            : std_logic;
  SIGNAL Logical_Operator_out980_out1            : std_logic;
  SIGNAL Logical_Operator_out981_out1            : std_logic;
  SIGNAL Logical_Operator_out982_out1            : std_logic;
  SIGNAL Logical_Operator_out983_out1            : std_logic;
  SIGNAL Logical_Operator_out984_out1            : std_logic;
  SIGNAL Logical_Operator_out985_out1            : std_logic;
  SIGNAL Logical_Operator_out986_out1            : std_logic;
  SIGNAL Logical_Operator_out987_out1            : std_logic;
  SIGNAL Logical_Operator_out988_out1            : std_logic;
  SIGNAL Logical_Operator_out989_out1            : std_logic;
  SIGNAL Logical_Operator_out990_out1            : std_logic;
  SIGNAL Logical_Operator_out991_out1            : std_logic;
  SIGNAL Logical_Operator_out992_out1            : std_logic;
  SIGNAL Logical_Operator_out993_out1            : std_logic;
  SIGNAL Logical_Operator_out994_out1            : std_logic;
  SIGNAL Logical_Operator_out995_out1            : std_logic;
  SIGNAL Logical_Operator_out996_out1            : std_logic;
  SIGNAL Logical_Operator_out997_out1            : std_logic;
  SIGNAL Logical_Operator_out998_out1            : std_logic;
  SIGNAL Logical_Operator_out999_out1            : std_logic;
  SIGNAL Logical_Operator_out1000_out1            : std_logic;
  SIGNAL Logical_Operator_out1001_out1            : std_logic;
  SIGNAL Logical_Operator_out1002_out1            : std_logic;
  SIGNAL Logical_Operator_out1003_out1            : std_logic;
  SIGNAL Logical_Operator_out1004_out1            : std_logic;
  SIGNAL Logical_Operator_out1005_out1            : std_logic;
  SIGNAL Logical_Operator_out1006_out1            : std_logic;
  SIGNAL Logical_Operator_out1007_out1            : std_logic;
  SIGNAL Logical_Operator_out1008_out1            : std_logic;
  SIGNAL Logical_Operator_out1009_out1            : std_logic;
  SIGNAL Logical_Operator_out1010_out1            : std_logic;
  SIGNAL Logical_Operator_out1011_out1            : std_logic;
  SIGNAL Logical_Operator_out1012_out1            : std_logic;
  SIGNAL Logical_Operator_out1013_out1            : std_logic;
  SIGNAL Logical_Operator_out1014_out1            : std_logic;
  SIGNAL Logical_Operator_out1015_out1            : std_logic;
  SIGNAL Logical_Operator_out1016_out1            : std_logic;
  SIGNAL Logical_Operator_out1017_out1            : std_logic;
  SIGNAL Logical_Operator_out1018_out1            : std_logic;
  SIGNAL Logical_Operator_out1019_out1            : std_logic;
  SIGNAL Logical_Operator_out1020_out1            : std_logic;
  SIGNAL Logical_Operator_out1021_out1            : std_logic;
  SIGNAL Logical_Operator_out1022_out1            : std_logic;
  SIGNAL Logical_Operator_out1023_out1            : std_logic;
  SIGNAL Logical_Operator_out1024_out1            : std_logic;
  SIGNAL Logical_Operator_out1025_out1            : std_logic;
  SIGNAL Logical_Operator_out1026_out1            : std_logic;
  SIGNAL Logical_Operator_out1027_out1            : std_logic;
  SIGNAL Logical_Operator_out1028_out1            : std_logic;
  SIGNAL Logical_Operator_out1029_out1            : std_logic;
  SIGNAL Logical_Operator_out1030_out1            : std_logic;
  SIGNAL Logical_Operator_out1031_out1            : std_logic;
  SIGNAL Logical_Operator_out1032_out1            : std_logic;
  SIGNAL Logical_Operator_out1033_out1            : std_logic;
  SIGNAL Logical_Operator_out1034_out1            : std_logic;
  SIGNAL Logical_Operator_out1035_out1            : std_logic;
  SIGNAL Logical_Operator_out1036_out1            : std_logic;
  SIGNAL Logical_Operator_out1037_out1            : std_logic;
  SIGNAL Logical_Operator_out1038_out1            : std_logic;
  SIGNAL Logical_Operator_out1039_out1            : std_logic;
  SIGNAL Logical_Operator_out1040_out1            : std_logic;
  SIGNAL Logical_Operator_out1041_out1            : std_logic;
  SIGNAL Logical_Operator_out1042_out1            : std_logic;
  SIGNAL Logical_Operator_out1043_out1            : std_logic;
  SIGNAL Logical_Operator_out1044_out1            : std_logic;
  SIGNAL Logical_Operator_out1045_out1            : std_logic;
  SIGNAL Logical_Operator_out1046_out1            : std_logic;
  SIGNAL Logical_Operator_out1047_out1            : std_logic;
  SIGNAL Logical_Operator_out1048_out1            : std_logic;
  SIGNAL Logical_Operator_out1049_out1            : std_logic;
  SIGNAL Logical_Operator_out1050_out1            : std_logic;
  SIGNAL Logical_Operator_out1051_out1            : std_logic;
  SIGNAL Logical_Operator_out1052_out1            : std_logic;
  SIGNAL Logical_Operator_out1053_out1            : std_logic;
  SIGNAL Logical_Operator_out1054_out1            : std_logic;
  SIGNAL Logical_Operator_out1055_out1            : std_logic;
  SIGNAL Logical_Operator_out1056_out1            : std_logic;
  SIGNAL Logical_Operator_out1057_out1            : std_logic;
  SIGNAL Logical_Operator_out1058_out1            : std_logic;
  SIGNAL Logical_Operator_out1059_out1            : std_logic;
  SIGNAL Logical_Operator_out1060_out1            : std_logic;
  SIGNAL Logical_Operator_out1061_out1            : std_logic;
  SIGNAL Logical_Operator_out1062_out1            : std_logic;
  SIGNAL Logical_Operator_out1063_out1            : std_logic;
  SIGNAL Logical_Operator_out1064_out1            : std_logic;
  SIGNAL Logical_Operator_out1065_out1            : std_logic;
  SIGNAL Logical_Operator_out1066_out1            : std_logic;
  SIGNAL Logical_Operator_out1067_out1            : std_logic;
  SIGNAL Logical_Operator_out1068_out1            : std_logic;
  SIGNAL Logical_Operator_out1069_out1            : std_logic;
  SIGNAL Logical_Operator_out1070_out1            : std_logic;
  SIGNAL Logical_Operator_out1071_out1            : std_logic;
  SIGNAL Logical_Operator_out1072_out1            : std_logic;
  SIGNAL Logical_Operator_out1073_out1            : std_logic;
  SIGNAL Logical_Operator_out1074_out1            : std_logic;
  SIGNAL Logical_Operator_out1075_out1            : std_logic;
  SIGNAL Logical_Operator_out1076_out1            : std_logic;
  SIGNAL Logical_Operator_out1077_out1            : std_logic;
  SIGNAL Logical_Operator_out1078_out1            : std_logic;
  SIGNAL Logical_Operator_out1079_out1            : std_logic;
  SIGNAL Logical_Operator_out1080_out1            : std_logic;
  SIGNAL Logical_Operator_out1081_out1            : std_logic;
  SIGNAL Logical_Operator_out1082_out1            : std_logic;
  SIGNAL Logical_Operator_out1083_out1            : std_logic;
  SIGNAL Logical_Operator_out1084_out1            : std_logic;
  SIGNAL Logical_Operator_out1085_out1            : std_logic;
  SIGNAL Logical_Operator_out1086_out1            : std_logic;
  SIGNAL Logical_Operator_out1087_out1            : std_logic;
  SIGNAL Logical_Operator_out1088_out1            : std_logic;
  SIGNAL Logical_Operator_out1089_out1            : std_logic;
  SIGNAL Logical_Operator_out1090_out1            : std_logic;
  SIGNAL Logical_Operator_out1091_out1            : std_logic;
  SIGNAL Logical_Operator_out1092_out1            : std_logic;
  SIGNAL Logical_Operator_out1093_out1            : std_logic;
  SIGNAL Logical_Operator_out1094_out1            : std_logic;
  SIGNAL Logical_Operator_out1095_out1            : std_logic;
  SIGNAL Logical_Operator_out1096_out1            : std_logic;
  SIGNAL Logical_Operator_out1097_out1            : std_logic;
  SIGNAL Logical_Operator_out1098_out1            : std_logic;
  SIGNAL Logical_Operator_out1099_out1            : std_logic;
  SIGNAL Logical_Operator_out1100_out1            : std_logic;
  SIGNAL Logical_Operator_out1101_out1            : std_logic;
  SIGNAL Logical_Operator_out1102_out1            : std_logic;
  SIGNAL Logical_Operator_out1103_out1            : std_logic;
  SIGNAL Logical_Operator_out1104_out1            : std_logic;
  SIGNAL Logical_Operator_out1105_out1            : std_logic;
  SIGNAL Logical_Operator_out1106_out1            : std_logic;
  SIGNAL Logical_Operator_out1107_out1            : std_logic;
  SIGNAL Logical_Operator_out1108_out1            : std_logic;
  SIGNAL Logical_Operator_out1109_out1            : std_logic;
  SIGNAL Logical_Operator_out1110_out1            : std_logic;
  SIGNAL Logical_Operator_out1111_out1            : std_logic;
  SIGNAL Logical_Operator_out1112_out1            : std_logic;
  SIGNAL Logical_Operator_out1113_out1            : std_logic;
  SIGNAL Logical_Operator_out1114_out1            : std_logic;
  SIGNAL Logical_Operator_out1115_out1            : std_logic;
  SIGNAL Logical_Operator_out1116_out1            : std_logic;
  SIGNAL Logical_Operator_out1117_out1            : std_logic;
  SIGNAL Logical_Operator_out1118_out1            : std_logic;
  SIGNAL Logical_Operator_out1119_out1            : std_logic;
  SIGNAL Logical_Operator_out1120_out1            : std_logic;
  SIGNAL Logical_Operator_out1121_out1            : std_logic;
  SIGNAL Logical_Operator_out1122_out1            : std_logic;
  SIGNAL Logical_Operator_out1123_out1            : std_logic;
  SIGNAL Logical_Operator_out1124_out1            : std_logic;
  SIGNAL Logical_Operator_out1125_out1            : std_logic;
  SIGNAL Logical_Operator_out1126_out1            : std_logic;
  SIGNAL Logical_Operator_out1127_out1            : std_logic;
  SIGNAL Logical_Operator_out1128_out1            : std_logic;
  SIGNAL Logical_Operator_out1129_out1            : std_logic;
  SIGNAL Logical_Operator_out1130_out1            : std_logic;
  SIGNAL Logical_Operator_out1131_out1            : std_logic;
  SIGNAL Logical_Operator_out1132_out1            : std_logic;
  SIGNAL Logical_Operator_out1133_out1            : std_logic;
  SIGNAL Logical_Operator_out1134_out1            : std_logic;
  SIGNAL Logical_Operator_out1135_out1            : std_logic;
  SIGNAL Logical_Operator_out1136_out1            : std_logic;
  SIGNAL Logical_Operator_out1137_out1            : std_logic;
  SIGNAL Logical_Operator_out1138_out1            : std_logic;
  SIGNAL Logical_Operator_out1139_out1            : std_logic;
  SIGNAL Logical_Operator_out1140_out1            : std_logic;
  SIGNAL Logical_Operator_out1141_out1            : std_logic;
  SIGNAL Logical_Operator_out1142_out1            : std_logic;
  SIGNAL Logical_Operator_out1143_out1            : std_logic;
  SIGNAL Logical_Operator_out1144_out1            : std_logic;
  SIGNAL Logical_Operator_out1145_out1            : std_logic;
  SIGNAL Logical_Operator_out1146_out1            : std_logic;
  SIGNAL Logical_Operator_out1147_out1            : std_logic;
  SIGNAL Logical_Operator_out1148_out1            : std_logic;
  SIGNAL Logical_Operator_out1149_out1            : std_logic;
  SIGNAL Logical_Operator_out1150_out1            : std_logic;
  SIGNAL Logical_Operator_out1151_out1            : std_logic;
  SIGNAL Logical_Operator_out1152_out1            : std_logic;
  SIGNAL Logical_Operator_out1153_out1            : std_logic;
  SIGNAL Logical_Operator_out1154_out1            : std_logic;
  SIGNAL Logical_Operator_out1155_out1            : std_logic;
  SIGNAL Logical_Operator_out1156_out1            : std_logic;
  SIGNAL Logical_Operator_out1157_out1            : std_logic;
  SIGNAL Logical_Operator_out1158_out1            : std_logic;
  SIGNAL Logical_Operator_out1159_out1            : std_logic;
  SIGNAL Logical_Operator_out1160_out1            : std_logic;
  SIGNAL Logical_Operator_out1161_out1            : std_logic;
  SIGNAL Logical_Operator_out1162_out1            : std_logic;
  SIGNAL Logical_Operator_out1163_out1            : std_logic;
  SIGNAL Logical_Operator_out1164_out1            : std_logic;
  SIGNAL Logical_Operator_out1165_out1            : std_logic;
  SIGNAL Logical_Operator_out1166_out1            : std_logic;
  SIGNAL Logical_Operator_out1167_out1            : std_logic;
  SIGNAL Logical_Operator_out1168_out1            : std_logic;
  SIGNAL Logical_Operator_out1169_out1            : std_logic;
  SIGNAL Logical_Operator_out1170_out1            : std_logic;
  SIGNAL Logical_Operator_out1171_out1            : std_logic;
  SIGNAL Logical_Operator_out1172_out1            : std_logic;
  SIGNAL Logical_Operator_out1173_out1            : std_logic;
  SIGNAL Logical_Operator_out1174_out1            : std_logic;
  SIGNAL Logical_Operator_out1175_out1            : std_logic;
  SIGNAL Logical_Operator_out1176_out1            : std_logic;
  SIGNAL Logical_Operator_out1177_out1            : std_logic;
  SIGNAL Logical_Operator_out1178_out1            : std_logic;
  SIGNAL Logical_Operator_out1179_out1            : std_logic;
  SIGNAL Logical_Operator_out1180_out1            : std_logic;
  SIGNAL Logical_Operator_out1181_out1            : std_logic;
  SIGNAL Logical_Operator_out1182_out1            : std_logic;
  SIGNAL Logical_Operator_out1183_out1            : std_logic;
  SIGNAL Logical_Operator_out1184_out1            : std_logic;
  SIGNAL Logical_Operator_out1185_out1            : std_logic;
  SIGNAL Logical_Operator_out1186_out1            : std_logic;
  SIGNAL Logical_Operator_out1187_out1            : std_logic;
  SIGNAL Logical_Operator_out1188_out1            : std_logic;
  SIGNAL Logical_Operator_out1189_out1            : std_logic;
  SIGNAL Logical_Operator_out1190_out1            : std_logic;
  SIGNAL Logical_Operator_out1191_out1            : std_logic;
  SIGNAL Logical_Operator_out1192_out1            : std_logic;
  SIGNAL Logical_Operator_out1193_out1            : std_logic;
  SIGNAL Logical_Operator_out1194_out1            : std_logic;
  SIGNAL Logical_Operator_out1195_out1            : std_logic;
  SIGNAL Logical_Operator_out1196_out1            : std_logic;
  SIGNAL Logical_Operator_out1197_out1            : std_logic;
  SIGNAL Logical_Operator_out1198_out1            : std_logic;
  SIGNAL Logical_Operator_out1199_out1            : std_logic;
  SIGNAL Logical_Operator_out1200_out1            : std_logic;
  SIGNAL Logical_Operator_out1201_out1            : std_logic;
  SIGNAL Logical_Operator_out1202_out1            : std_logic;
  SIGNAL Logical_Operator_out1203_out1            : std_logic;
  SIGNAL Logical_Operator_out1204_out1            : std_logic;
  SIGNAL Logical_Operator_out1205_out1            : std_logic;
  SIGNAL Logical_Operator_out1206_out1            : std_logic;
  SIGNAL Logical_Operator_out1207_out1            : std_logic;
  SIGNAL Logical_Operator_out1208_out1            : std_logic;
  SIGNAL Logical_Operator_out1209_out1            : std_logic;
  SIGNAL Logical_Operator_out1210_out1            : std_logic;
  SIGNAL Logical_Operator_out1211_out1            : std_logic;
  SIGNAL Logical_Operator_out1212_out1            : std_logic;
  SIGNAL Logical_Operator_out1213_out1            : std_logic;
  SIGNAL Logical_Operator_out1214_out1            : std_logic;
  SIGNAL Logical_Operator_out1215_out1            : std_logic;
  SIGNAL Logical_Operator_out1216_out1            : std_logic;
  SIGNAL Logical_Operator_out1217_out1            : std_logic;
  SIGNAL Logical_Operator_out1218_out1            : std_logic;
  SIGNAL Logical_Operator_out1219_out1            : std_logic;
  SIGNAL Logical_Operator_out1220_out1            : std_logic;
  SIGNAL Logical_Operator_out1221_out1            : std_logic;
  SIGNAL Logical_Operator_out1222_out1            : std_logic;
  SIGNAL Logical_Operator_out1223_out1            : std_logic;
  SIGNAL Logical_Operator_out1224_out1            : std_logic;
  SIGNAL Logical_Operator_out1225_out1            : std_logic;
  SIGNAL Logical_Operator_out1226_out1            : std_logic;
  SIGNAL Logical_Operator_out1227_out1            : std_logic;
  SIGNAL Logical_Operator_out1228_out1            : std_logic;
  SIGNAL Logical_Operator_out1229_out1            : std_logic;
  SIGNAL Logical_Operator_out1230_out1            : std_logic;
  SIGNAL Logical_Operator_out1231_out1            : std_logic;
  SIGNAL Logical_Operator_out1232_out1            : std_logic;
  SIGNAL Logical_Operator_out1233_out1            : std_logic;
  SIGNAL Logical_Operator_out1234_out1            : std_logic;
  SIGNAL Logical_Operator_out1235_out1            : std_logic;
  SIGNAL Logical_Operator_out1236_out1            : std_logic;
  SIGNAL Logical_Operator_out1237_out1            : std_logic;
  SIGNAL Logical_Operator_out1238_out1            : std_logic;
  SIGNAL Logical_Operator_out1239_out1            : std_logic;
  SIGNAL Logical_Operator_out1240_out1            : std_logic;
  SIGNAL Logical_Operator_out1241_out1            : std_logic;
  SIGNAL Logical_Operator_out1242_out1            : std_logic;
  SIGNAL Logical_Operator_out1243_out1            : std_logic;
  SIGNAL Logical_Operator_out1244_out1            : std_logic;
  SIGNAL Logical_Operator_out1245_out1            : std_logic;
  SIGNAL Logical_Operator_out1246_out1            : std_logic;
  SIGNAL Logical_Operator_out1247_out1            : std_logic;
  SIGNAL Logical_Operator_out1248_out1            : std_logic;
  SIGNAL Logical_Operator_out1249_out1            : std_logic;
  SIGNAL Logical_Operator_out1250_out1            : std_logic;
  SIGNAL Logical_Operator_out1251_out1            : std_logic;
  SIGNAL Logical_Operator_out1252_out1            : std_logic;
  SIGNAL Logical_Operator_out1253_out1            : std_logic;
  SIGNAL Logical_Operator_out1254_out1            : std_logic;
  SIGNAL Logical_Operator_out1255_out1            : std_logic;
  SIGNAL Logical_Operator_out1256_out1            : std_logic;
  SIGNAL Logical_Operator_out1257_out1            : std_logic;
  SIGNAL Logical_Operator_out1258_out1            : std_logic;
  SIGNAL Logical_Operator_out1259_out1            : std_logic;
  SIGNAL Logical_Operator_out1260_out1            : std_logic;
  SIGNAL Logical_Operator_out1261_out1            : std_logic;
  SIGNAL Logical_Operator_out1262_out1            : std_logic;
  SIGNAL Logical_Operator_out1263_out1            : std_logic;
  SIGNAL Logical_Operator_out1264_out1            : std_logic;
  SIGNAL Logical_Operator_out1265_out1            : std_logic;
  SIGNAL Logical_Operator_out1266_out1            : std_logic;
  SIGNAL Logical_Operator_out1267_out1            : std_logic;
  SIGNAL Logical_Operator_out1268_out1            : std_logic;
  SIGNAL Logical_Operator_out1269_out1            : std_logic;
  SIGNAL Logical_Operator_out1270_out1            : std_logic;
  SIGNAL Logical_Operator_out1271_out1            : std_logic;
  SIGNAL Logical_Operator_out1272_out1            : std_logic;
  SIGNAL Logical_Operator_out1273_out1            : std_logic;
  SIGNAL Logical_Operator_out1274_out1            : std_logic;
  SIGNAL Logical_Operator_out1275_out1            : std_logic;
  SIGNAL Logical_Operator_out1276_out1            : std_logic;
  SIGNAL Logical_Operator_out1277_out1            : std_logic;
  SIGNAL Logical_Operator_out1278_out1            : std_logic;
  SIGNAL Logical_Operator_out1279_out1            : std_logic;
  SIGNAL Logical_Operator_out1280_out1            : std_logic;
  SIGNAL Logical_Operator_out1281_out1            : std_logic;
  SIGNAL Logical_Operator_out1282_out1            : std_logic;
  SIGNAL Logical_Operator_out1283_out1            : std_logic;
  SIGNAL Logical_Operator_out1284_out1            : std_logic;
  SIGNAL Logical_Operator_out1285_out1            : std_logic;
  SIGNAL Logical_Operator_out1286_out1            : std_logic;
  SIGNAL Logical_Operator_out1287_out1            : std_logic;
  SIGNAL Logical_Operator_out1288_out1            : std_logic;
  SIGNAL Logical_Operator_out1289_out1            : std_logic;
  SIGNAL Logical_Operator_out1290_out1            : std_logic;
  SIGNAL Logical_Operator_out1291_out1            : std_logic;
  SIGNAL Logical_Operator_out1292_out1            : std_logic;
  SIGNAL Logical_Operator_out1293_out1            : std_logic;
  SIGNAL Logical_Operator_out1294_out1            : std_logic;
  SIGNAL Logical_Operator_out1295_out1            : std_logic;
  SIGNAL Logical_Operator_out1296_out1            : std_logic;
  SIGNAL Logical_Operator_out1297_out1            : std_logic;
  SIGNAL Logical_Operator_out1298_out1            : std_logic;
  SIGNAL Logical_Operator_out1299_out1            : std_logic;
  SIGNAL Logical_Operator_out1300_out1            : std_logic;
  SIGNAL Logical_Operator_out1301_out1            : std_logic;
  SIGNAL Logical_Operator_out1302_out1            : std_logic;
  SIGNAL Logical_Operator_out1303_out1            : std_logic;
  SIGNAL Logical_Operator_out1304_out1            : std_logic;
  SIGNAL Logical_Operator_out1305_out1            : std_logic;
  SIGNAL Logical_Operator_out1306_out1            : std_logic;
  SIGNAL Logical_Operator_out1307_out1            : std_logic;
  SIGNAL Logical_Operator_out1308_out1            : std_logic;
  SIGNAL Logical_Operator_out1309_out1            : std_logic;
  SIGNAL Logical_Operator_out1310_out1            : std_logic;
  SIGNAL Logical_Operator_out1311_out1            : std_logic;
  SIGNAL Logical_Operator_out1312_out1            : std_logic;
  SIGNAL Logical_Operator_out1313_out1            : std_logic;
  SIGNAL Logical_Operator_out1314_out1            : std_logic;
  SIGNAL Logical_Operator_out1315_out1            : std_logic;
  SIGNAL Logical_Operator_out1316_out1            : std_logic;
  SIGNAL Logical_Operator_out1317_out1            : std_logic;
  SIGNAL Logical_Operator_out1318_out1            : std_logic;
  SIGNAL Logical_Operator_out1319_out1            : std_logic;
  SIGNAL Logical_Operator_out1320_out1            : std_logic;
  SIGNAL Logical_Operator_out1321_out1            : std_logic;
  SIGNAL Logical_Operator_out1322_out1            : std_logic;
  SIGNAL Logical_Operator_out1323_out1            : std_logic;
  SIGNAL Logical_Operator_out1324_out1            : std_logic;
  SIGNAL Logical_Operator_out1325_out1            : std_logic;
  SIGNAL Logical_Operator_out1326_out1            : std_logic;
  SIGNAL Logical_Operator_out1327_out1            : std_logic;
  SIGNAL Logical_Operator_out1328_out1            : std_logic;
  SIGNAL Logical_Operator_out1329_out1            : std_logic;
  SIGNAL Logical_Operator_out1330_out1            : std_logic;
  SIGNAL Logical_Operator_out1331_out1            : std_logic;
  SIGNAL Logical_Operator_out1332_out1            : std_logic;
  SIGNAL Logical_Operator_out1333_out1            : std_logic;
  SIGNAL Logical_Operator_out1334_out1            : std_logic;
  SIGNAL Logical_Operator_out1335_out1            : std_logic;
  SIGNAL Logical_Operator_out1336_out1            : std_logic;
  SIGNAL Logical_Operator_out1337_out1            : std_logic;
  SIGNAL Logical_Operator_out1338_out1            : std_logic;
  SIGNAL Logical_Operator_out1339_out1            : std_logic;
  SIGNAL Logical_Operator_out1340_out1            : std_logic;
  SIGNAL Logical_Operator_out1341_out1            : std_logic;
  SIGNAL Logical_Operator_out1342_out1            : std_logic;
  SIGNAL Logical_Operator_out1343_out1            : std_logic;
  SIGNAL Logical_Operator_out1344_out1            : std_logic;
  SIGNAL Logical_Operator_out1345_out1            : std_logic;
  SIGNAL Logical_Operator_out1346_out1            : std_logic;
  SIGNAL Logical_Operator_out1347_out1            : std_logic;
  SIGNAL Logical_Operator_out1348_out1            : std_logic;
  SIGNAL Logical_Operator_out1349_out1            : std_logic;
  SIGNAL Logical_Operator_out1350_out1            : std_logic;
  SIGNAL Logical_Operator_out1351_out1            : std_logic;
  SIGNAL Logical_Operator_out1352_out1            : std_logic;
  SIGNAL Logical_Operator_out1353_out1            : std_logic;
  SIGNAL Logical_Operator_out1354_out1            : std_logic;
  SIGNAL Logical_Operator_out1355_out1            : std_logic;
  SIGNAL Logical_Operator_out1356_out1            : std_logic;
  SIGNAL Logical_Operator_out1357_out1            : std_logic;
  SIGNAL Logical_Operator_out1358_out1            : std_logic;
  SIGNAL Logical_Operator_out1359_out1            : std_logic;
  SIGNAL Logical_Operator_out1360_out1            : std_logic;
  SIGNAL Logical_Operator_out1361_out1            : std_logic;
  SIGNAL Logical_Operator_out1362_out1            : std_logic;
  SIGNAL Logical_Operator_out1363_out1            : std_logic;
  SIGNAL Logical_Operator_out1364_out1            : std_logic;
  SIGNAL Logical_Operator_out1365_out1            : std_logic;
  SIGNAL Logical_Operator_out1366_out1            : std_logic;
  SIGNAL Logical_Operator_out1367_out1            : std_logic;
  SIGNAL Logical_Operator_out1368_out1            : std_logic;
  SIGNAL Logical_Operator_out1369_out1            : std_logic;
  SIGNAL Logical_Operator_out1370_out1            : std_logic;
  SIGNAL Logical_Operator_out1371_out1            : std_logic;
  SIGNAL Logical_Operator_out1372_out1            : std_logic;
  SIGNAL Logical_Operator_out1373_out1            : std_logic;
  SIGNAL Logical_Operator_out1374_out1            : std_logic;
  SIGNAL Logical_Operator_out1375_out1            : std_logic;
  SIGNAL Logical_Operator_out1376_out1            : std_logic;
  SIGNAL Logical_Operator_out1377_out1            : std_logic;
  SIGNAL Logical_Operator_out1378_out1            : std_logic;
  SIGNAL Logical_Operator_out1379_out1            : std_logic;
  SIGNAL Logical_Operator_out1380_out1            : std_logic;
  SIGNAL Logical_Operator_out1381_out1            : std_logic;
  SIGNAL Logical_Operator_out1382_out1            : std_logic;
  SIGNAL Logical_Operator_out1383_out1            : std_logic;
  SIGNAL Logical_Operator_out1384_out1            : std_logic;
  SIGNAL Logical_Operator_out1385_out1            : std_logic;
  SIGNAL Logical_Operator_out1386_out1            : std_logic;
  SIGNAL Logical_Operator_out1387_out1            : std_logic;
  SIGNAL Logical_Operator_out1388_out1            : std_logic;
  SIGNAL Logical_Operator_out1389_out1            : std_logic;
  SIGNAL Logical_Operator_out1390_out1            : std_logic;
  SIGNAL Logical_Operator_out1391_out1            : std_logic;
  SIGNAL Logical_Operator_out1392_out1            : std_logic;
  SIGNAL Logical_Operator_out1393_out1            : std_logic;
  SIGNAL Logical_Operator_out1394_out1            : std_logic;
  SIGNAL Logical_Operator_out1395_out1            : std_logic;
  SIGNAL Logical_Operator_out1396_out1            : std_logic;
  SIGNAL Logical_Operator_out1397_out1            : std_logic;
  SIGNAL Logical_Operator_out1398_out1            : std_logic;
  SIGNAL Logical_Operator_out1399_out1            : std_logic;
  SIGNAL Logical_Operator_out1400_out1            : std_logic;
  SIGNAL Logical_Operator_out1401_out1            : std_logic;
  SIGNAL Logical_Operator_out1402_out1            : std_logic;
  SIGNAL Logical_Operator_out1403_out1            : std_logic;
  SIGNAL Logical_Operator_out1404_out1            : std_logic;
  SIGNAL Logical_Operator_out1405_out1            : std_logic;
  SIGNAL Logical_Operator_out1406_out1            : std_logic;
  SIGNAL Logical_Operator_out1407_out1            : std_logic;
  SIGNAL Logical_Operator_out1408_out1            : std_logic;
  SIGNAL Logical_Operator_out1409_out1            : std_logic;
  SIGNAL Logical_Operator_out1410_out1            : std_logic;
  SIGNAL Logical_Operator_out1411_out1            : std_logic;
  SIGNAL Logical_Operator_out1412_out1            : std_logic;
  SIGNAL Logical_Operator_out1413_out1            : std_logic;
  SIGNAL Logical_Operator_out1414_out1            : std_logic;
  SIGNAL Logical_Operator_out1415_out1            : std_logic;
  SIGNAL Logical_Operator_out1416_out1            : std_logic;
  SIGNAL Logical_Operator_out1417_out1            : std_logic;
  SIGNAL Logical_Operator_out1418_out1            : std_logic;
  SIGNAL Logical_Operator_out1419_out1            : std_logic;
  SIGNAL Logical_Operator_out1420_out1            : std_logic;
  SIGNAL Logical_Operator_out1421_out1            : std_logic;
  SIGNAL Logical_Operator_out1422_out1            : std_logic;
  SIGNAL Logical_Operator_out1423_out1            : std_logic;
  SIGNAL Logical_Operator_out1424_out1            : std_logic;
  SIGNAL Logical_Operator_out1425_out1            : std_logic;
  SIGNAL Logical_Operator_out1426_out1            : std_logic;
  SIGNAL Logical_Operator_out1427_out1            : std_logic;
  SIGNAL Logical_Operator_out1428_out1            : std_logic;
  SIGNAL Logical_Operator_out1429_out1            : std_logic;
  SIGNAL Logical_Operator_out1430_out1            : std_logic;
  SIGNAL Logical_Operator_out1431_out1            : std_logic;
  SIGNAL Logical_Operator_out1432_out1            : std_logic;
  SIGNAL Logical_Operator_out1433_out1            : std_logic;
  SIGNAL Logical_Operator_out1434_out1            : std_logic;
  SIGNAL Logical_Operator_out1435_out1            : std_logic;
  SIGNAL Logical_Operator_out1436_out1            : std_logic;
  SIGNAL Logical_Operator_out1437_out1            : std_logic;
  SIGNAL Logical_Operator_out1438_out1            : std_logic;
  SIGNAL Logical_Operator_out1439_out1            : std_logic;
  SIGNAL Logical_Operator_out1440_out1            : std_logic;
  SIGNAL Logical_Operator_out1441_out1            : std_logic;
  SIGNAL Logical_Operator_out1442_out1            : std_logic;
  SIGNAL Logical_Operator_out1443_out1            : std_logic;
  SIGNAL Logical_Operator_out1444_out1            : std_logic;
  SIGNAL Logical_Operator_out1445_out1            : std_logic;
  SIGNAL Logical_Operator_out1446_out1            : std_logic;
  SIGNAL Logical_Operator_out1447_out1            : std_logic;
  SIGNAL Logical_Operator_out1448_out1            : std_logic;
  SIGNAL Logical_Operator_out1449_out1            : std_logic;
  SIGNAL Logical_Operator_out1450_out1            : std_logic;
  SIGNAL Logical_Operator_out1451_out1            : std_logic;
  SIGNAL Logical_Operator_out1452_out1            : std_logic;
  SIGNAL Logical_Operator_out1453_out1            : std_logic;
  SIGNAL Logical_Operator_out1454_out1            : std_logic;
  SIGNAL Logical_Operator_out1455_out1            : std_logic;
  SIGNAL Logical_Operator_out1456_out1            : std_logic;
  SIGNAL Logical_Operator_out1457_out1            : std_logic;
  SIGNAL Logical_Operator_out1458_out1            : std_logic;
  SIGNAL Logical_Operator_out1459_out1            : std_logic;
  SIGNAL Logical_Operator_out1460_out1            : std_logic;
  SIGNAL Logical_Operator_out1461_out1            : std_logic;
  SIGNAL Logical_Operator_out1462_out1            : std_logic;
  SIGNAL Logical_Operator_out1463_out1            : std_logic;
  SIGNAL Logical_Operator_out1464_out1            : std_logic;
  SIGNAL Logical_Operator_out1465_out1            : std_logic;
  SIGNAL Logical_Operator_out1466_out1            : std_logic;
  SIGNAL Logical_Operator_out1467_out1            : std_logic;
  SIGNAL Logical_Operator_out1468_out1            : std_logic;
  SIGNAL Logical_Operator_out1469_out1            : std_logic;
  SIGNAL Logical_Operator_out1470_out1            : std_logic;
  SIGNAL Logical_Operator_out1471_out1            : std_logic;
  SIGNAL Logical_Operator_out1472_out1            : std_logic;
  SIGNAL Logical_Operator_out1473_out1            : std_logic;
  SIGNAL Logical_Operator_out1474_out1            : std_logic;
  SIGNAL Logical_Operator_out1475_out1            : std_logic;
  SIGNAL Logical_Operator_out1476_out1            : std_logic;
  SIGNAL Logical_Operator_out1477_out1            : std_logic;
  SIGNAL Logical_Operator_out1478_out1            : std_logic;
  SIGNAL Logical_Operator_out1479_out1            : std_logic;
  SIGNAL Logical_Operator_out1480_out1            : std_logic;
  SIGNAL Logical_Operator_out1481_out1            : std_logic;
  SIGNAL Logical_Operator_out1482_out1            : std_logic;
  SIGNAL Logical_Operator_out1483_out1            : std_logic;
  SIGNAL Logical_Operator_out1484_out1            : std_logic;
  SIGNAL Logical_Operator_out1485_out1            : std_logic;
  SIGNAL Logical_Operator_out1486_out1            : std_logic;
  SIGNAL Logical_Operator_out1487_out1            : std_logic;
  SIGNAL Logical_Operator_out1488_out1            : std_logic;
  SIGNAL Logical_Operator_out1489_out1            : std_logic;
  SIGNAL Logical_Operator_out1490_out1            : std_logic;
  SIGNAL Logical_Operator_out1491_out1            : std_logic;
  SIGNAL Logical_Operator_out1492_out1            : std_logic;
  SIGNAL Logical_Operator_out1493_out1            : std_logic;
  SIGNAL Logical_Operator_out1494_out1            : std_logic;
  SIGNAL Logical_Operator_out1495_out1            : std_logic;
  SIGNAL Logical_Operator_out1496_out1            : std_logic;
  SIGNAL Logical_Operator_out1497_out1            : std_logic;
  SIGNAL Logical_Operator_out1498_out1            : std_logic;
  SIGNAL Logical_Operator_out1499_out1            : std_logic;
  SIGNAL Logical_Operator_out1500_out1            : std_logic;
  SIGNAL Logical_Operator_out1501_out1            : std_logic;
  SIGNAL Logical_Operator_out1502_out1            : std_logic;
  SIGNAL Logical_Operator_out1503_out1            : std_logic;
  SIGNAL Logical_Operator_out1504_out1            : std_logic;
  SIGNAL Logical_Operator_out1505_out1            : std_logic;
  SIGNAL Logical_Operator_out1506_out1            : std_logic;
  SIGNAL Logical_Operator_out1507_out1            : std_logic;
  SIGNAL Logical_Operator_out1508_out1            : std_logic;
  SIGNAL Logical_Operator_out1509_out1            : std_logic;
  SIGNAL Logical_Operator_out1510_out1            : std_logic;
  SIGNAL Logical_Operator_out1511_out1            : std_logic;
  SIGNAL Logical_Operator_out1512_out1            : std_logic;
  SIGNAL Logical_Operator_out1513_out1            : std_logic;
  SIGNAL Logical_Operator_out1514_out1            : std_logic;
  SIGNAL Logical_Operator_out1515_out1            : std_logic;
  SIGNAL Logical_Operator_out1516_out1            : std_logic;
  SIGNAL Logical_Operator_out1517_out1            : std_logic;
  SIGNAL Logical_Operator_out1518_out1            : std_logic;
  SIGNAL Logical_Operator_out1519_out1            : std_logic;
  SIGNAL Logical_Operator_out1520_out1            : std_logic;
  SIGNAL Logical_Operator_out1521_out1            : std_logic;
  SIGNAL Logical_Operator_out1522_out1            : std_logic;
  SIGNAL Logical_Operator_out1523_out1            : std_logic;
  SIGNAL Logical_Operator_out1524_out1            : std_logic;
  SIGNAL Logical_Operator_out1525_out1            : std_logic;
  SIGNAL Logical_Operator_out1526_out1            : std_logic;
  SIGNAL Logical_Operator_out1527_out1            : std_logic;
  SIGNAL Logical_Operator_out1528_out1            : std_logic;
  SIGNAL Logical_Operator_out1529_out1            : std_logic;
  SIGNAL Logical_Operator_out1530_out1            : std_logic;
  SIGNAL Logical_Operator_out1531_out1            : std_logic;
  SIGNAL Logical_Operator_out1532_out1            : std_logic;
  SIGNAL Logical_Operator_out1533_out1            : std_logic;
  SIGNAL Logical_Operator_out1534_out1            : std_logic;
  SIGNAL Logical_Operator_out1535_out1            : std_logic;
  SIGNAL Logical_Operator_out1536_out1            : std_logic;
  SIGNAL Logical_Operator_out1537_out1            : std_logic;
  SIGNAL Logical_Operator_out1538_out1            : std_logic;
  SIGNAL Logical_Operator_out1539_out1            : std_logic;
  SIGNAL Logical_Operator_out1540_out1            : std_logic;
  SIGNAL Logical_Operator_out1541_out1            : std_logic;
  SIGNAL Logical_Operator_out1542_out1            : std_logic;
  SIGNAL Logical_Operator_out1543_out1            : std_logic;
  SIGNAL Logical_Operator_out1544_out1            : std_logic;
  SIGNAL Logical_Operator_out1545_out1            : std_logic;
  SIGNAL Logical_Operator_out1546_out1            : std_logic;
  SIGNAL Logical_Operator_out1547_out1            : std_logic;
  SIGNAL Logical_Operator_out1548_out1            : std_logic;
  SIGNAL Logical_Operator_out1549_out1            : std_logic;
  SIGNAL Logical_Operator_out1550_out1            : std_logic;
  SIGNAL Logical_Operator_out1551_out1            : std_logic;
  SIGNAL Logical_Operator_out1552_out1            : std_logic;
  SIGNAL Logical_Operator_out1553_out1            : std_logic;
  SIGNAL Logical_Operator_out1554_out1            : std_logic;
  SIGNAL Logical_Operator_out1555_out1            : std_logic;
  SIGNAL Logical_Operator_out1556_out1            : std_logic;
  SIGNAL Logical_Operator_out1557_out1            : std_logic;
  SIGNAL Logical_Operator_out1558_out1            : std_logic;
  SIGNAL Logical_Operator_out1559_out1            : std_logic;
  SIGNAL Logical_Operator_out1560_out1            : std_logic;
  SIGNAL Logical_Operator_out1561_out1            : std_logic;
  SIGNAL Logical_Operator_out1562_out1            : std_logic;
  SIGNAL Logical_Operator_out1563_out1            : std_logic;
  SIGNAL Logical_Operator_out1564_out1            : std_logic;
  SIGNAL Logical_Operator_out1565_out1            : std_logic;
  SIGNAL Logical_Operator_out1566_out1            : std_logic;
  SIGNAL Logical_Operator_out1567_out1            : std_logic;
  SIGNAL Logical_Operator_out1568_out1            : std_logic;
  SIGNAL Logical_Operator_out1569_out1            : std_logic;
  SIGNAL Logical_Operator_out1570_out1            : std_logic;
  SIGNAL Logical_Operator_out1571_out1            : std_logic;
  SIGNAL Logical_Operator_out1572_out1            : std_logic;
  SIGNAL Logical_Operator_out1573_out1            : std_logic;
  SIGNAL Logical_Operator_out1574_out1            : std_logic;
  SIGNAL Logical_Operator_out1575_out1            : std_logic;
  SIGNAL Logical_Operator_out1576_out1            : std_logic;
  SIGNAL Logical_Operator_out1577_out1            : std_logic;
  SIGNAL Logical_Operator_out1578_out1            : std_logic;
  SIGNAL Logical_Operator_out1579_out1            : std_logic;
  SIGNAL Logical_Operator_out1580_out1            : std_logic;
  SIGNAL Logical_Operator_out1581_out1            : std_logic;
  SIGNAL Logical_Operator_out1582_out1            : std_logic;
  SIGNAL Logical_Operator_out1583_out1            : std_logic;
  SIGNAL Logical_Operator_out1584_out1            : std_logic;
  SIGNAL Logical_Operator_out1585_out1            : std_logic;
  SIGNAL Logical_Operator_out1586_out1            : std_logic;
  SIGNAL Logical_Operator_out1587_out1            : std_logic;
  SIGNAL Logical_Operator_out1588_out1            : std_logic;
  SIGNAL Logical_Operator_out1589_out1            : std_logic;
  SIGNAL Logical_Operator_out1590_out1            : std_logic;
  SIGNAL Logical_Operator_out1591_out1            : std_logic;
  SIGNAL Logical_Operator_out1592_out1            : std_logic;
  SIGNAL Logical_Operator_out1593_out1            : std_logic;
  SIGNAL Logical_Operator_out1594_out1            : std_logic;
  SIGNAL Logical_Operator_out1595_out1            : std_logic;
  SIGNAL Logical_Operator_out1596_out1            : std_logic;
  SIGNAL Logical_Operator_out1597_out1            : std_logic;
  SIGNAL Logical_Operator_out1598_out1            : std_logic;
  SIGNAL Logical_Operator_out1599_out1            : std_logic;
  SIGNAL Logical_Operator_out1600_out1            : std_logic;
  SIGNAL Logical_Operator_out1601_out1            : std_logic;
  SIGNAL Logical_Operator_out1602_out1            : std_logic;
  SIGNAL Logical_Operator_out1603_out1            : std_logic;
  SIGNAL Logical_Operator_out1604_out1            : std_logic;
  SIGNAL Logical_Operator_out1605_out1            : std_logic;
  SIGNAL Logical_Operator_out1606_out1            : std_logic;
  SIGNAL Logical_Operator_out1607_out1            : std_logic;
  SIGNAL Logical_Operator_out1608_out1            : std_logic;
  SIGNAL Logical_Operator_out1609_out1            : std_logic;
  SIGNAL Logical_Operator_out1610_out1            : std_logic;
  SIGNAL Logical_Operator_out1611_out1            : std_logic;
  SIGNAL Logical_Operator_out1612_out1            : std_logic;
  SIGNAL Logical_Operator_out1613_out1            : std_logic;
  SIGNAL Logical_Operator_out1614_out1            : std_logic;
  SIGNAL Logical_Operator_out1615_out1            : std_logic;
  SIGNAL Logical_Operator_out1616_out1            : std_logic;
  SIGNAL Logical_Operator_out1617_out1            : std_logic;
  SIGNAL Logical_Operator_out1618_out1            : std_logic;
  SIGNAL Logical_Operator_out1619_out1            : std_logic;
  SIGNAL Logical_Operator_out1620_out1            : std_logic;
  SIGNAL Logical_Operator_out1621_out1            : std_logic;
  SIGNAL Logical_Operator_out1622_out1            : std_logic;
  SIGNAL Logical_Operator_out1623_out1            : std_logic;
  SIGNAL Logical_Operator_out1624_out1            : std_logic;
  SIGNAL Logical_Operator_out1625_out1            : std_logic;
  SIGNAL Logical_Operator_out1626_out1            : std_logic;
  SIGNAL Logical_Operator_out1627_out1            : std_logic;
  SIGNAL Logical_Operator_out1628_out1            : std_logic;
  SIGNAL Logical_Operator_out1629_out1            : std_logic;
  SIGNAL Logical_Operator_out1630_out1            : std_logic;
  SIGNAL Logical_Operator_out1631_out1            : std_logic;
  SIGNAL Logical_Operator_out1632_out1            : std_logic;
  SIGNAL Logical_Operator_out1633_out1            : std_logic;
  SIGNAL Logical_Operator_out1634_out1            : std_logic;
  SIGNAL Logical_Operator_out1635_out1            : std_logic;
  SIGNAL Logical_Operator_out1636_out1            : std_logic;
  SIGNAL Logical_Operator_out1637_out1            : std_logic;
  SIGNAL Logical_Operator_out1638_out1            : std_logic;
  SIGNAL Logical_Operator_out1639_out1            : std_logic;
  SIGNAL Logical_Operator_out1640_out1            : std_logic;
  SIGNAL Logical_Operator_out1641_out1            : std_logic;
  SIGNAL Logical_Operator_out1642_out1            : std_logic;
  SIGNAL Logical_Operator_out1643_out1            : std_logic;
  SIGNAL Logical_Operator_out1644_out1            : std_logic;
  SIGNAL Logical_Operator_out1645_out1            : std_logic;
  SIGNAL Logical_Operator_out1646_out1            : std_logic;
  SIGNAL Logical_Operator_out1647_out1            : std_logic;
  SIGNAL Logical_Operator_out1648_out1            : std_logic;
  SIGNAL Logical_Operator_out1649_out1            : std_logic;
  SIGNAL Logical_Operator_out1650_out1            : std_logic;
  SIGNAL Logical_Operator_out1651_out1            : std_logic;
  SIGNAL Logical_Operator_out1652_out1            : std_logic;
  SIGNAL Logical_Operator_out1653_out1            : std_logic;
  SIGNAL Logical_Operator_out1654_out1            : std_logic;
  SIGNAL Logical_Operator_out1655_out1            : std_logic;
  SIGNAL Logical_Operator_out1656_out1            : std_logic;
  SIGNAL Logical_Operator_out1657_out1            : std_logic;
  SIGNAL Logical_Operator_out1658_out1            : std_logic;
  SIGNAL Logical_Operator_out1659_out1            : std_logic;
  SIGNAL Logical_Operator_out1660_out1            : std_logic;
  SIGNAL Logical_Operator_out1661_out1            : std_logic;
  SIGNAL Logical_Operator_out1662_out1            : std_logic;
  SIGNAL Logical_Operator_out1663_out1            : std_logic;
  SIGNAL Logical_Operator_out1664_out1            : std_logic;
  SIGNAL Logical_Operator_out1665_out1            : std_logic;
  SIGNAL Logical_Operator_out1666_out1            : std_logic;
  SIGNAL Logical_Operator_out1667_out1            : std_logic;
  SIGNAL Logical_Operator_out1668_out1            : std_logic;
  SIGNAL Logical_Operator_out1669_out1            : std_logic;
  SIGNAL Logical_Operator_out1670_out1            : std_logic;
  SIGNAL Logical_Operator_out1671_out1            : std_logic;
  SIGNAL Logical_Operator_out1672_out1            : std_logic;
  SIGNAL Logical_Operator_out1673_out1            : std_logic;
  SIGNAL Logical_Operator_out1674_out1            : std_logic;
  SIGNAL Logical_Operator_out1675_out1            : std_logic;
  SIGNAL Logical_Operator_out1676_out1            : std_logic;
  SIGNAL Logical_Operator_out1677_out1            : std_logic;
  SIGNAL Logical_Operator_out1678_out1            : std_logic;
  SIGNAL Logical_Operator_out1679_out1            : std_logic;
  SIGNAL Logical_Operator_out1680_out1            : std_logic;
  SIGNAL Logical_Operator_out1681_out1            : std_logic;
  SIGNAL Logical_Operator_out1682_out1            : std_logic;
  SIGNAL Logical_Operator_out1683_out1            : std_logic;
  SIGNAL Logical_Operator_out1684_out1            : std_logic;
  SIGNAL Logical_Operator_out1685_out1            : std_logic;
  SIGNAL Logical_Operator_out1686_out1            : std_logic;
  SIGNAL Logical_Operator_out1687_out1            : std_logic;
  SIGNAL Logical_Operator_out1688_out1            : std_logic;
  SIGNAL Logical_Operator_out1689_out1            : std_logic;
  SIGNAL Logical_Operator_out1690_out1            : std_logic;
  SIGNAL Logical_Operator_out1691_out1            : std_logic;
  SIGNAL Logical_Operator_out1692_out1            : std_logic;
  SIGNAL Logical_Operator_out1693_out1            : std_logic;
  SIGNAL Logical_Operator_out1694_out1            : std_logic;
  SIGNAL Logical_Operator_out1695_out1            : std_logic;
  SIGNAL Logical_Operator_out1696_out1            : std_logic;
  SIGNAL Logical_Operator_out1697_out1            : std_logic;
  SIGNAL Logical_Operator_out1698_out1            : std_logic;
  SIGNAL Logical_Operator_out1699_out1            : std_logic;
  SIGNAL Logical_Operator_out1700_out1            : std_logic;
  SIGNAL Logical_Operator_out1701_out1            : std_logic;
  SIGNAL Logical_Operator_out1702_out1            : std_logic;
  SIGNAL Logical_Operator_out1703_out1            : std_logic;
  SIGNAL Logical_Operator_out1704_out1            : std_logic;
  SIGNAL Logical_Operator_out1705_out1            : std_logic;
  SIGNAL Logical_Operator_out1706_out1            : std_logic;
  SIGNAL Logical_Operator_out1707_out1            : std_logic;
  SIGNAL Logical_Operator_out1708_out1            : std_logic;
  SIGNAL Logical_Operator_out1709_out1            : std_logic;
  SIGNAL Logical_Operator_out1710_out1            : std_logic;
  SIGNAL Logical_Operator_out1711_out1            : std_logic;
  SIGNAL Logical_Operator_out1712_out1            : std_logic;
  SIGNAL Logical_Operator_out1713_out1            : std_logic;
  SIGNAL Logical_Operator_out1714_out1            : std_logic;
  SIGNAL Logical_Operator_out1715_out1            : std_logic;
  SIGNAL Logical_Operator_out1716_out1            : std_logic;
  SIGNAL Logical_Operator_out1717_out1            : std_logic;
  SIGNAL Logical_Operator_out1718_out1            : std_logic;
  SIGNAL Logical_Operator_out1719_out1            : std_logic;
  SIGNAL Logical_Operator_out1720_out1            : std_logic;
  SIGNAL Logical_Operator_out1721_out1            : std_logic;
  SIGNAL Logical_Operator_out1722_out1            : std_logic;
  SIGNAL Logical_Operator_out1723_out1            : std_logic;
  SIGNAL Logical_Operator_out1724_out1            : std_logic;
  SIGNAL Logical_Operator_out1725_out1            : std_logic;
  SIGNAL Logical_Operator_out1726_out1            : std_logic;
  SIGNAL Logical_Operator_out1727_out1            : std_logic;
  SIGNAL Logical_Operator_out1728_out1            : std_logic;
  SIGNAL Logical_Operator_out1729_out1            : std_logic;
  SIGNAL Logical_Operator_out1730_out1            : std_logic;
  SIGNAL Logical_Operator_out1731_out1            : std_logic;
  SIGNAL Logical_Operator_out1732_out1            : std_logic;
  SIGNAL Logical_Operator_out1733_out1            : std_logic;
  SIGNAL Logical_Operator_out1734_out1            : std_logic;
  SIGNAL Logical_Operator_out1735_out1            : std_logic;
  SIGNAL Logical_Operator_out1736_out1            : std_logic;
  SIGNAL Logical_Operator_out1737_out1            : std_logic;
  SIGNAL Logical_Operator_out1738_out1            : std_logic;
  SIGNAL Logical_Operator_out1739_out1            : std_logic;
  SIGNAL Logical_Operator_out1740_out1            : std_logic;
  SIGNAL Logical_Operator_out1741_out1            : std_logic;
  SIGNAL Logical_Operator_out1742_out1            : std_logic;
  SIGNAL Logical_Operator_out1743_out1            : std_logic;
  SIGNAL Logical_Operator_out1744_out1            : std_logic;
  SIGNAL Logical_Operator_out1745_out1            : std_logic;
  SIGNAL Logical_Operator_out1746_out1            : std_logic;
  SIGNAL Logical_Operator_out1747_out1            : std_logic;
  SIGNAL Logical_Operator_out1748_out1            : std_logic;
  SIGNAL Logical_Operator_out1749_out1            : std_logic;
  SIGNAL Logical_Operator_out1750_out1            : std_logic;
  SIGNAL Logical_Operator_out1751_out1            : std_logic;
  SIGNAL Logical_Operator_out1752_out1            : std_logic;
  SIGNAL Logical_Operator_out1753_out1            : std_logic;
  SIGNAL Logical_Operator_out1754_out1            : std_logic;
  SIGNAL Logical_Operator_out1755_out1            : std_logic;
  SIGNAL Logical_Operator_out1756_out1            : std_logic;
  SIGNAL Logical_Operator_out1757_out1            : std_logic;
  SIGNAL Logical_Operator_out1758_out1            : std_logic;
  SIGNAL Logical_Operator_out1759_out1            : std_logic;
  SIGNAL Logical_Operator_out1760_out1            : std_logic;
  SIGNAL Logical_Operator_out1761_out1            : std_logic;
  SIGNAL Logical_Operator_out1762_out1            : std_logic;
  SIGNAL Logical_Operator_out1763_out1            : std_logic;
  SIGNAL Logical_Operator_out1764_out1            : std_logic;
  SIGNAL Logical_Operator_out1765_out1            : std_logic;
  SIGNAL Logical_Operator_out1766_out1            : std_logic;
  SIGNAL Logical_Operator_out1767_out1            : std_logic;
  SIGNAL Logical_Operator_out1768_out1            : std_logic;
  SIGNAL Logical_Operator_out1769_out1            : std_logic;
  SIGNAL Logical_Operator_out1770_out1            : std_logic;
  SIGNAL Logical_Operator_out1771_out1            : std_logic;
  SIGNAL Logical_Operator_out1772_out1            : std_logic;
  SIGNAL Logical_Operator_out1773_out1            : std_logic;
  SIGNAL Logical_Operator_out1774_out1            : std_logic;
  SIGNAL Logical_Operator_out1775_out1            : std_logic;
  SIGNAL Logical_Operator_out1776_out1            : std_logic;
  SIGNAL Logical_Operator_out1777_out1            : std_logic;
  SIGNAL Logical_Operator_out1778_out1            : std_logic;
  SIGNAL Logical_Operator_out1779_out1            : std_logic;
  SIGNAL Logical_Operator_out1780_out1            : std_logic;
  SIGNAL Logical_Operator_out1781_out1            : std_logic;
  SIGNAL Logical_Operator_out1782_out1            : std_logic;
  SIGNAL Logical_Operator_out1783_out1            : std_logic;
  SIGNAL Logical_Operator_out1784_out1            : std_logic;
  SIGNAL Logical_Operator_out1785_out1            : std_logic;
  SIGNAL Logical_Operator_out1786_out1            : std_logic;
  SIGNAL Logical_Operator_out1787_out1            : std_logic;
  SIGNAL Logical_Operator_out1788_out1            : std_logic;
  SIGNAL Logical_Operator_out1789_out1            : std_logic;
  SIGNAL Logical_Operator_out1790_out1            : std_logic;
  SIGNAL Logical_Operator_out1791_out1            : std_logic;
  SIGNAL Logical_Operator_out1792_out1            : std_logic;
  SIGNAL Logical_Operator_out1793_out1            : std_logic;
  SIGNAL Logical_Operator_out1794_out1            : std_logic;
  SIGNAL Logical_Operator_out1795_out1            : std_logic;
  SIGNAL Logical_Operator_out1796_out1            : std_logic;
  SIGNAL Logical_Operator_out1797_out1            : std_logic;
  SIGNAL Logical_Operator_out1798_out1            : std_logic;
  SIGNAL Logical_Operator_out1799_out1            : std_logic;
  SIGNAL Logical_Operator_out1800_out1            : std_logic;
  SIGNAL Logical_Operator_out1801_out1            : std_logic;
  SIGNAL Logical_Operator_out1802_out1            : std_logic;
  SIGNAL Logical_Operator_out1803_out1            : std_logic;
  SIGNAL Logical_Operator_out1804_out1            : std_logic;
  SIGNAL Logical_Operator_out1805_out1            : std_logic;
  SIGNAL Logical_Operator_out1806_out1            : std_logic;
  SIGNAL Logical_Operator_out1807_out1            : std_logic;
  SIGNAL Logical_Operator_out1808_out1            : std_logic;
  SIGNAL Logical_Operator_out1809_out1            : std_logic;
  SIGNAL Logical_Operator_out1810_out1            : std_logic;
  SIGNAL Logical_Operator_out1811_out1            : std_logic;
  SIGNAL Logical_Operator_out1812_out1            : std_logic;
  SIGNAL Logical_Operator_out1813_out1            : std_logic;
  SIGNAL Logical_Operator_out1814_out1            : std_logic;
  SIGNAL Logical_Operator_out1815_out1            : std_logic;
  SIGNAL Logical_Operator_out1816_out1            : std_logic;
  SIGNAL Logical_Operator_out1817_out1            : std_logic;
  SIGNAL Logical_Operator_out1818_out1            : std_logic;
  SIGNAL Logical_Operator_out1819_out1            : std_logic;
  SIGNAL Logical_Operator_out1820_out1            : std_logic;
  SIGNAL Logical_Operator_out1821_out1            : std_logic;
  SIGNAL Logical_Operator_out1822_out1            : std_logic;
  SIGNAL Logical_Operator_out1823_out1            : std_logic;
  SIGNAL Logical_Operator_out1824_out1            : std_logic;
  SIGNAL Logical_Operator_out1825_out1            : std_logic;
  SIGNAL Logical_Operator_out1826_out1            : std_logic;
  SIGNAL Logical_Operator_out1827_out1            : std_logic;
  SIGNAL Logical_Operator_out1828_out1            : std_logic;
  SIGNAL Logical_Operator_out1829_out1            : std_logic;
  SIGNAL Logical_Operator_out1830_out1            : std_logic;
  SIGNAL Logical_Operator_out1831_out1            : std_logic;
  SIGNAL Logical_Operator_out1832_out1            : std_logic;
  SIGNAL Logical_Operator_out1833_out1            : std_logic;
  SIGNAL Logical_Operator_out1834_out1            : std_logic;
  SIGNAL Logical_Operator_out1835_out1            : std_logic;
  SIGNAL Logical_Operator_out1836_out1            : std_logic;
  SIGNAL Logical_Operator_out1837_out1            : std_logic;
  SIGNAL Logical_Operator_out1838_out1            : std_logic;
  SIGNAL Logical_Operator_out1839_out1            : std_logic;
  SIGNAL Logical_Operator_out1840_out1            : std_logic;
  SIGNAL Logical_Operator_out1841_out1            : std_logic;
  SIGNAL Logical_Operator_out1842_out1            : std_logic;
  SIGNAL Logical_Operator_out1843_out1            : std_logic;
  SIGNAL Logical_Operator_out1844_out1            : std_logic;
  SIGNAL Logical_Operator_out1845_out1            : std_logic;
  SIGNAL Logical_Operator_out1846_out1            : std_logic;
  SIGNAL Logical_Operator_out1847_out1            : std_logic;
  SIGNAL Logical_Operator_out1848_out1            : std_logic;
  SIGNAL Logical_Operator_out1849_out1            : std_logic;
  SIGNAL Logical_Operator_out1850_out1            : std_logic;
  SIGNAL Logical_Operator_out1851_out1            : std_logic;
  SIGNAL Logical_Operator_out1852_out1            : std_logic;
  SIGNAL Logical_Operator_out1853_out1            : std_logic;
  SIGNAL Logical_Operator_out1854_out1            : std_logic;
  SIGNAL Logical_Operator_out1855_out1            : std_logic;
  SIGNAL Logical_Operator_out1856_out1            : std_logic;
  SIGNAL Logical_Operator_out1857_out1            : std_logic;
  SIGNAL Logical_Operator_out1858_out1            : std_logic;
  SIGNAL Logical_Operator_out1859_out1            : std_logic;
  SIGNAL Logical_Operator_out1860_out1            : std_logic;
  SIGNAL Logical_Operator_out1861_out1            : std_logic;
  SIGNAL Logical_Operator_out1862_out1            : std_logic;
  SIGNAL Logical_Operator_out1863_out1            : std_logic;
  SIGNAL Logical_Operator_out1864_out1            : std_logic;
  SIGNAL Logical_Operator_out1865_out1            : std_logic;
  SIGNAL Logical_Operator_out1866_out1            : std_logic;
  SIGNAL Logical_Operator_out1867_out1            : std_logic;
  SIGNAL Logical_Operator_out1868_out1            : std_logic;
  SIGNAL Logical_Operator_out1869_out1            : std_logic;
  SIGNAL Logical_Operator_out1870_out1            : std_logic;
  SIGNAL Logical_Operator_out1871_out1            : std_logic;
  SIGNAL Logical_Operator_out1872_out1            : std_logic;
  SIGNAL Logical_Operator_out1873_out1            : std_logic;
  SIGNAL Logical_Operator_out1874_out1            : std_logic;
  SIGNAL Logical_Operator_out1875_out1            : std_logic;
  SIGNAL Logical_Operator_out1876_out1            : std_logic;
  SIGNAL Logical_Operator_out1877_out1            : std_logic;
  SIGNAL Logical_Operator_out1878_out1            : std_logic;
  SIGNAL Logical_Operator_out1879_out1            : std_logic;
  SIGNAL Logical_Operator_out1880_out1            : std_logic;
  SIGNAL Logical_Operator_out1881_out1            : std_logic;
  SIGNAL Logical_Operator_out1882_out1            : std_logic;
  SIGNAL Logical_Operator_out1883_out1            : std_logic;
  SIGNAL Logical_Operator_out1884_out1            : std_logic;
  SIGNAL Logical_Operator_out1885_out1            : std_logic;
  SIGNAL Logical_Operator_out1886_out1            : std_logic;
  SIGNAL Logical_Operator_out1887_out1            : std_logic;
  SIGNAL Logical_Operator_out1888_out1            : std_logic;
  SIGNAL Logical_Operator_out1889_out1            : std_logic;
  SIGNAL Logical_Operator_out1890_out1            : std_logic;
  SIGNAL Logical_Operator_out1891_out1            : std_logic;
  SIGNAL Logical_Operator_out1892_out1            : std_logic;
  SIGNAL Logical_Operator_out1893_out1            : std_logic;
  SIGNAL Logical_Operator_out1894_out1            : std_logic;
  SIGNAL Logical_Operator_out1895_out1            : std_logic;
  SIGNAL Logical_Operator_out1896_out1            : std_logic;
  SIGNAL Logical_Operator_out1897_out1            : std_logic;
  SIGNAL Logical_Operator_out1898_out1            : std_logic;
  SIGNAL Logical_Operator_out1899_out1            : std_logic;
  SIGNAL Logical_Operator_out1900_out1            : std_logic;
  SIGNAL Logical_Operator_out1901_out1            : std_logic;
  SIGNAL Logical_Operator_out1902_out1            : std_logic;
  SIGNAL Logical_Operator_out1903_out1            : std_logic;
  SIGNAL Logical_Operator_out1904_out1            : std_logic;
  SIGNAL Logical_Operator_out1905_out1            : std_logic;
  SIGNAL Logical_Operator_out1906_out1            : std_logic;
  SIGNAL Logical_Operator_out1907_out1            : std_logic;
  SIGNAL Logical_Operator_out1908_out1            : std_logic;
  SIGNAL Logical_Operator_out1909_out1            : std_logic;
  SIGNAL Logical_Operator_out1910_out1            : std_logic;
  SIGNAL Logical_Operator_out1911_out1            : std_logic;
  SIGNAL Logical_Operator_out1912_out1            : std_logic;
  SIGNAL Logical_Operator_out1913_out1            : std_logic;
  SIGNAL Logical_Operator_out1914_out1            : std_logic;
  SIGNAL Logical_Operator_out1915_out1            : std_logic;
  SIGNAL Logical_Operator_out1916_out1            : std_logic;
  SIGNAL Logical_Operator_out1917_out1            : std_logic;
  SIGNAL Logical_Operator_out1918_out1            : std_logic;
  SIGNAL Logical_Operator_out1919_out1            : std_logic;
  SIGNAL Logical_Operator_out1920_out1            : std_logic;
  SIGNAL Logical_Operator_out1921_out1            : std_logic;
  SIGNAL Logical_Operator_out1922_out1            : std_logic;
  SIGNAL Logical_Operator_out1923_out1            : std_logic;
  SIGNAL Logical_Operator_out1924_out1            : std_logic;
  SIGNAL Logical_Operator_out1925_out1            : std_logic;
  SIGNAL Logical_Operator_out1926_out1            : std_logic;
  SIGNAL Logical_Operator_out1927_out1            : std_logic;
  SIGNAL Logical_Operator_out1928_out1            : std_logic;
  SIGNAL Logical_Operator_out1929_out1            : std_logic;
  SIGNAL Logical_Operator_out1930_out1            : std_logic;
  SIGNAL Logical_Operator_out1931_out1            : std_logic;
  SIGNAL Logical_Operator_out1932_out1            : std_logic;
  SIGNAL Logical_Operator_out1933_out1            : std_logic;
  SIGNAL Logical_Operator_out1934_out1            : std_logic;
  SIGNAL Logical_Operator_out1935_out1            : std_logic;
  SIGNAL Logical_Operator_out1936_out1            : std_logic;
  SIGNAL Logical_Operator_out1937_out1            : std_logic;
  SIGNAL Logical_Operator_out1938_out1            : std_logic;
  SIGNAL Logical_Operator_out1939_out1            : std_logic;
  SIGNAL Logical_Operator_out1940_out1            : std_logic;
  SIGNAL Logical_Operator_out1941_out1            : std_logic;
  SIGNAL Logical_Operator_out1942_out1            : std_logic;
  SIGNAL Logical_Operator_out1943_out1            : std_logic;
  SIGNAL Logical_Operator_out1944_out1            : std_logic;
  SIGNAL Logical_Operator_out1945_out1            : std_logic;
  SIGNAL Logical_Operator_out1946_out1            : std_logic;
  SIGNAL Logical_Operator_out1947_out1            : std_logic;
  SIGNAL Logical_Operator_out1948_out1            : std_logic;
  SIGNAL Logical_Operator_out1949_out1            : std_logic;
  SIGNAL Logical_Operator_out1950_out1            : std_logic;
  SIGNAL Logical_Operator_out1951_out1            : std_logic;
  SIGNAL Logical_Operator_out1952_out1            : std_logic;
  SIGNAL Logical_Operator_out1953_out1            : std_logic;
  SIGNAL Logical_Operator_out1954_out1            : std_logic;
  SIGNAL Logical_Operator_out1955_out1            : std_logic;
  SIGNAL Logical_Operator_out1956_out1            : std_logic;
  SIGNAL Logical_Operator_out1957_out1            : std_logic;
  SIGNAL Logical_Operator_out1958_out1            : std_logic;
  SIGNAL Logical_Operator_out1959_out1            : std_logic;
  SIGNAL Logical_Operator_out1960_out1            : std_logic;
  SIGNAL Logical_Operator_out1961_out1            : std_logic;
  SIGNAL Logical_Operator_out1962_out1            : std_logic;
  SIGNAL Logical_Operator_out1963_out1            : std_logic;
  SIGNAL Logical_Operator_out1964_out1            : std_logic;
  SIGNAL Logical_Operator_out1965_out1            : std_logic;
  SIGNAL Logical_Operator_out1966_out1            : std_logic;
  SIGNAL Logical_Operator_out1967_out1            : std_logic;
  SIGNAL Logical_Operator_out1968_out1            : std_logic;
  SIGNAL Logical_Operator_out1969_out1            : std_logic;
  SIGNAL Logical_Operator_out1970_out1            : std_logic;
  SIGNAL Logical_Operator_out1971_out1            : std_logic;
  SIGNAL Logical_Operator_out1972_out1            : std_logic;
  SIGNAL Logical_Operator_out1973_out1            : std_logic;
  SIGNAL Logical_Operator_out1974_out1            : std_logic;
  SIGNAL Logical_Operator_out1975_out1            : std_logic;
  SIGNAL Logical_Operator_out1976_out1            : std_logic;
  SIGNAL Logical_Operator_out1977_out1            : std_logic;
  SIGNAL Logical_Operator_out1978_out1            : std_logic;
  SIGNAL Logical_Operator_out1979_out1            : std_logic;
  SIGNAL Logical_Operator_out1980_out1            : std_logic;
  SIGNAL Logical_Operator_out1981_out1            : std_logic;
  SIGNAL Logical_Operator_out1982_out1            : std_logic;
  SIGNAL Logical_Operator_out1983_out1            : std_logic;
  SIGNAL Logical_Operator_out1984_out1            : std_logic;
  SIGNAL Logical_Operator_out1985_out1            : std_logic;
  SIGNAL Logical_Operator_out1986_out1            : std_logic;
  SIGNAL Logical_Operator_out1987_out1            : std_logic;
  SIGNAL Logical_Operator_out1988_out1            : std_logic;
  SIGNAL Logical_Operator_out1989_out1            : std_logic;
  SIGNAL Logical_Operator_out1990_out1            : std_logic;
  SIGNAL Logical_Operator_out1991_out1            : std_logic;
  SIGNAL Logical_Operator_out1992_out1            : std_logic;
  SIGNAL Logical_Operator_out1993_out1            : std_logic;
  SIGNAL Logical_Operator_out1994_out1            : std_logic;
  SIGNAL Logical_Operator_out1995_out1            : std_logic;
  SIGNAL Logical_Operator_out1996_out1            : std_logic;
  SIGNAL Logical_Operator_out1997_out1            : std_logic;
  SIGNAL Logical_Operator_out1998_out1            : std_logic;
  SIGNAL Logical_Operator_out1999_out1            : std_logic;
  SIGNAL Logical_Operator_out2000_out1            : std_logic;
  SIGNAL Logical_Operator_out2001_out1            : std_logic;
  SIGNAL Logical_Operator_out2002_out1            : std_logic;
  SIGNAL Logical_Operator_out2003_out1            : std_logic;
  SIGNAL Logical_Operator_out2004_out1            : std_logic;
  SIGNAL Logical_Operator_out2005_out1            : std_logic;
  SIGNAL Logical_Operator_out2006_out1            : std_logic;
  SIGNAL Logical_Operator_out2007_out1            : std_logic;
  SIGNAL Logical_Operator_out2008_out1            : std_logic;
  SIGNAL Logical_Operator_out2009_out1            : std_logic;
  SIGNAL Logical_Operator_out2010_out1            : std_logic;
  SIGNAL Logical_Operator_out2011_out1            : std_logic;
  SIGNAL Logical_Operator_out2012_out1            : std_logic;
  SIGNAL Logical_Operator_out2013_out1            : std_logic;
  SIGNAL Logical_Operator_out2014_out1            : std_logic;
  SIGNAL Logical_Operator_out2015_out1            : std_logic;
  SIGNAL Logical_Operator_out2016_out1            : std_logic;
  SIGNAL Logical_Operator_out2017_out1            : std_logic;
  SIGNAL Logical_Operator_out2018_out1            : std_logic;
  SIGNAL Logical_Operator_out2019_out1            : std_logic;
  SIGNAL Logical_Operator_out2020_out1            : std_logic;
  SIGNAL Logical_Operator_out2021_out1            : std_logic;
  SIGNAL Logical_Operator_out2022_out1            : std_logic;
  SIGNAL Logical_Operator_out2023_out1            : std_logic;
  SIGNAL Logical_Operator_out2024_out1            : std_logic;
  SIGNAL Logical_Operator_out2025_out1            : std_logic;
  SIGNAL Logical_Operator_out2026_out1            : std_logic;
  SIGNAL Logical_Operator_out2027_out1            : std_logic;
  SIGNAL Logical_Operator_out2028_out1            : std_logic;
  SIGNAL Logical_Operator_out2029_out1            : std_logic;
  SIGNAL Logical_Operator_out2030_out1            : std_logic;
  SIGNAL Logical_Operator_out2031_out1            : std_logic;
  SIGNAL Logical_Operator_out2032_out1            : std_logic;
  SIGNAL Logical_Operator_out2033_out1            : std_logic;
  SIGNAL Logical_Operator_out2034_out1            : std_logic;
  SIGNAL Logical_Operator_out2035_out1            : std_logic;
  SIGNAL Logical_Operator_out2036_out1            : std_logic;
  SIGNAL Logical_Operator_out2037_out1            : std_logic;
  SIGNAL Logical_Operator_out2038_out1            : std_logic;
  SIGNAL Logical_Operator_out2039_out1            : std_logic;
  SIGNAL Logical_Operator_out2040_out1            : std_logic;
  SIGNAL Logical_Operator_out2041_out1            : std_logic;
  SIGNAL Logical_Operator_out2042_out1            : std_logic;
  SIGNAL Logical_Operator_out2043_out1            : std_logic;
  SIGNAL Logical_Operator_out2044_out1            : std_logic;
  SIGNAL Logical_Operator_out2045_out1            : std_logic;
  SIGNAL Logical_Operator_out2046_out1            : std_logic;
  SIGNAL Logical_Operator_out2047_out1            : std_logic;
  SIGNAL Logical_Operator_out2048_out1            : std_logic;
  SIGNAL Logical_Operator_out2049_out1            : std_logic;
  SIGNAL Logical_Operator_out2050_out1            : std_logic;
  SIGNAL Logical_Operator_out2051_out1            : std_logic;
  SIGNAL Logical_Operator_out2052_out1            : std_logic;
  SIGNAL Logical_Operator_out2053_out1            : std_logic;
  SIGNAL Logical_Operator_out2054_out1            : std_logic;
  SIGNAL Logical_Operator_out2055_out1            : std_logic;
  SIGNAL Logical_Operator_out2056_out1            : std_logic;
  SIGNAL Logical_Operator_out2057_out1            : std_logic;
  SIGNAL Logical_Operator_out2058_out1            : std_logic;
  SIGNAL Logical_Operator_out2059_out1            : std_logic;
  SIGNAL Logical_Operator_out2060_out1            : std_logic;
  SIGNAL Logical_Operator_out2061_out1            : std_logic;
  SIGNAL Logical_Operator_out2062_out1            : std_logic;
  SIGNAL Logical_Operator_out2063_out1            : std_logic;
  SIGNAL Logical_Operator_out2064_out1            : std_logic;
  SIGNAL Logical_Operator_out2065_out1            : std_logic;
  SIGNAL Logical_Operator_out2066_out1            : std_logic;
  SIGNAL Logical_Operator_out2067_out1            : std_logic;
  SIGNAL Logical_Operator_out2068_out1            : std_logic;
  SIGNAL Logical_Operator_out2069_out1            : std_logic;
  SIGNAL Logical_Operator_out2070_out1            : std_logic;
  SIGNAL Logical_Operator_out2071_out1            : std_logic;
  SIGNAL Logical_Operator_out2072_out1            : std_logic;
  SIGNAL Logical_Operator_out2073_out1            : std_logic;
  SIGNAL Logical_Operator_out2074_out1            : std_logic;
  SIGNAL Logical_Operator_out2075_out1            : std_logic;
  SIGNAL Logical_Operator_out2076_out1            : std_logic;
  SIGNAL Logical_Operator_out2077_out1            : std_logic;
  SIGNAL Logical_Operator_out2078_out1            : std_logic;
  SIGNAL Logical_Operator_out2079_out1            : std_logic;
  SIGNAL Logical_Operator_out2080_out1            : std_logic;
  SIGNAL Logical_Operator_out2081_out1            : std_logic;
  SIGNAL Logical_Operator_out2082_out1            : std_logic;
  SIGNAL Logical_Operator_out2083_out1            : std_logic;
  SIGNAL Logical_Operator_out2084_out1            : std_logic;
  SIGNAL Logical_Operator_out2085_out1            : std_logic;
  SIGNAL Logical_Operator_out2086_out1            : std_logic;
  SIGNAL Logical_Operator_out2087_out1            : std_logic;
  SIGNAL Logical_Operator_out2088_out1            : std_logic;
  SIGNAL Logical_Operator_out2089_out1            : std_logic;
  SIGNAL Logical_Operator_out2090_out1            : std_logic;
  SIGNAL Logical_Operator_out2091_out1            : std_logic;
  SIGNAL Logical_Operator_out2092_out1            : std_logic;
  SIGNAL Logical_Operator_out2093_out1            : std_logic;
  SIGNAL Logical_Operator_out2094_out1            : std_logic;
  SIGNAL Logical_Operator_out2095_out1            : std_logic;
  SIGNAL Logical_Operator_out2096_out1            : std_logic;
  SIGNAL Logical_Operator_out2097_out1            : std_logic;
  SIGNAL Logical_Operator_out2098_out1            : std_logic;
  SIGNAL Logical_Operator_out2099_out1            : std_logic;
  SIGNAL Logical_Operator_out2100_out1            : std_logic;
  SIGNAL Logical_Operator_out2101_out1            : std_logic;
  SIGNAL Logical_Operator_out2102_out1            : std_logic;
  SIGNAL Logical_Operator_out2103_out1            : std_logic;
  SIGNAL Logical_Operator_out2104_out1            : std_logic;
  SIGNAL Logical_Operator_out2105_out1            : std_logic;
  SIGNAL Logical_Operator_out2106_out1            : std_logic;
  SIGNAL Logical_Operator_out2107_out1            : std_logic;
  SIGNAL Logical_Operator_out2108_out1            : std_logic;
  SIGNAL Logical_Operator_out2109_out1            : std_logic;
  SIGNAL Logical_Operator_out2110_out1            : std_logic;
  SIGNAL Logical_Operator_out2111_out1            : std_logic;
  SIGNAL Logical_Operator_out2112_out1            : std_logic;
  SIGNAL Logical_Operator_out2113_out1            : std_logic;
  SIGNAL Logical_Operator_out2114_out1            : std_logic;
  SIGNAL Logical_Operator_out2115_out1            : std_logic;
  SIGNAL Logical_Operator_out2116_out1            : std_logic;
  SIGNAL Logical_Operator_out2117_out1            : std_logic;
  SIGNAL Logical_Operator_out2118_out1            : std_logic;
  SIGNAL Logical_Operator_out2119_out1            : std_logic;
  SIGNAL Logical_Operator_out2120_out1            : std_logic;
  SIGNAL Logical_Operator_out2121_out1            : std_logic;
  SIGNAL Logical_Operator_out2122_out1            : std_logic;
  SIGNAL Logical_Operator_out2123_out1            : std_logic;
  SIGNAL Logical_Operator_out2124_out1            : std_logic;
  SIGNAL Logical_Operator_out2125_out1            : std_logic;
  SIGNAL Logical_Operator_out2126_out1            : std_logic;
  SIGNAL Logical_Operator_out2127_out1            : std_logic;
  SIGNAL Logical_Operator_out2128_out1            : std_logic;
  SIGNAL Logical_Operator_out2129_out1            : std_logic;
  SIGNAL Logical_Operator_out2130_out1            : std_logic;
  SIGNAL Logical_Operator_out2131_out1            : std_logic;
  SIGNAL Logical_Operator_out2132_out1            : std_logic;
  SIGNAL Logical_Operator_out2133_out1            : std_logic;
  SIGNAL Logical_Operator_out2134_out1            : std_logic;
  SIGNAL Logical_Operator_out2135_out1            : std_logic;
  SIGNAL Logical_Operator_out2136_out1            : std_logic;
  SIGNAL Logical_Operator_out2137_out1            : std_logic;
  SIGNAL Logical_Operator_out2138_out1            : std_logic;
  SIGNAL Logical_Operator_out2139_out1            : std_logic;
  SIGNAL Logical_Operator_out2140_out1            : std_logic;
  SIGNAL Logical_Operator_out2141_out1            : std_logic;
  SIGNAL Logical_Operator_out2142_out1            : std_logic;
  SIGNAL Logical_Operator_out2143_out1            : std_logic;
  SIGNAL Logical_Operator_out2144_out1            : std_logic;
  SIGNAL Logical_Operator_out2145_out1            : std_logic;
  SIGNAL Logical_Operator_out2146_out1            : std_logic;
  SIGNAL Logical_Operator_out2147_out1            : std_logic;
  SIGNAL Logical_Operator_out2148_out1            : std_logic;
  SIGNAL Logical_Operator_out2149_out1            : std_logic;
  SIGNAL Logical_Operator_out2150_out1            : std_logic;
  SIGNAL Logical_Operator_out2151_out1            : std_logic;
  SIGNAL Logical_Operator_out2152_out1            : std_logic;
  SIGNAL Logical_Operator_out2153_out1            : std_logic;
  SIGNAL Logical_Operator_out2154_out1            : std_logic;
  SIGNAL Logical_Operator_out2155_out1            : std_logic;
  SIGNAL Logical_Operator_out2156_out1            : std_logic;
  SIGNAL Logical_Operator_out2157_out1            : std_logic;
  SIGNAL Logical_Operator_out2158_out1            : std_logic;
  SIGNAL Logical_Operator_out2159_out1            : std_logic;
  SIGNAL Logical_Operator_out2160_out1            : std_logic;
  SIGNAL Logical_Operator_out2161_out1            : std_logic;
  SIGNAL Logical_Operator_out2162_out1            : std_logic;
  SIGNAL Logical_Operator_out2163_out1            : std_logic;
  SIGNAL Logical_Operator_out2164_out1            : std_logic;
  SIGNAL Logical_Operator_out2165_out1            : std_logic;
  SIGNAL Logical_Operator_out2166_out1            : std_logic;
  SIGNAL Logical_Operator_out2167_out1            : std_logic;
  SIGNAL Logical_Operator_out2168_out1            : std_logic;
  SIGNAL Logical_Operator_out2169_out1            : std_logic;
  SIGNAL Logical_Operator_out2170_out1            : std_logic;
  SIGNAL Logical_Operator_out2171_out1            : std_logic;
  SIGNAL Logical_Operator_out2172_out1            : std_logic;
  SIGNAL Logical_Operator_out2173_out1            : std_logic;
  SIGNAL Logical_Operator_out2174_out1            : std_logic;
  SIGNAL Logical_Operator_out2175_out1            : std_logic;
  SIGNAL Logical_Operator_out2176_out1            : std_logic;
  SIGNAL Logical_Operator_out2177_out1            : std_logic;
  SIGNAL Logical_Operator_out2178_out1            : std_logic;
  SIGNAL Logical_Operator_out2179_out1            : std_logic;
  SIGNAL Logical_Operator_out2180_out1            : std_logic;
  SIGNAL Logical_Operator_out2181_out1            : std_logic;
  SIGNAL Logical_Operator_out2182_out1            : std_logic;
  SIGNAL Logical_Operator_out2183_out1            : std_logic;
  SIGNAL Logical_Operator_out2184_out1            : std_logic;
  SIGNAL Logical_Operator_out2185_out1            : std_logic;
  SIGNAL Logical_Operator_out2186_out1            : std_logic;
  SIGNAL Logical_Operator_out2187_out1            : std_logic;
  SIGNAL Logical_Operator_out2188_out1            : std_logic;
  SIGNAL Logical_Operator_out2189_out1            : std_logic;
  SIGNAL Logical_Operator_out2190_out1            : std_logic;
  SIGNAL Logical_Operator_out2191_out1            : std_logic;
  SIGNAL Logical_Operator_out2192_out1            : std_logic;
  SIGNAL Logical_Operator_out2193_out1            : std_logic;
  SIGNAL Logical_Operator_out2194_out1            : std_logic;
  SIGNAL Logical_Operator_out2195_out1            : std_logic;
  SIGNAL Logical_Operator_out2196_out1            : std_logic;
  SIGNAL Logical_Operator_out2197_out1            : std_logic;
  SIGNAL Logical_Operator_out2198_out1            : std_logic;
  SIGNAL Logical_Operator_out2199_out1            : std_logic;
  SIGNAL Logical_Operator_out2200_out1            : std_logic;
  SIGNAL Logical_Operator_out2201_out1            : std_logic;
  SIGNAL Logical_Operator_out2202_out1            : std_logic;
  SIGNAL Logical_Operator_out2203_out1            : std_logic;
  SIGNAL Logical_Operator_out2204_out1            : std_logic;
  SIGNAL Logical_Operator_out2205_out1            : std_logic;
  SIGNAL Logical_Operator_out2206_out1            : std_logic;
  SIGNAL Logical_Operator_out2207_out1            : std_logic;
  SIGNAL Logical_Operator_out2208_out1            : std_logic;
  SIGNAL Logical_Operator_out2209_out1            : std_logic;
  SIGNAL Logical_Operator_out2210_out1            : std_logic;
  SIGNAL Logical_Operator_out2211_out1            : std_logic;
  SIGNAL Logical_Operator_out2212_out1            : std_logic;
  SIGNAL Logical_Operator_out2213_out1            : std_logic;
  SIGNAL Logical_Operator_out2214_out1            : std_logic;
  SIGNAL Logical_Operator_out2215_out1            : std_logic;
  SIGNAL Logical_Operator_out2216_out1            : std_logic;
  SIGNAL Logical_Operator_out2217_out1            : std_logic;
  SIGNAL Logical_Operator_out2218_out1            : std_logic;
  SIGNAL Logical_Operator_out2219_out1            : std_logic;
  SIGNAL Logical_Operator_out2220_out1            : std_logic;
  SIGNAL Logical_Operator_out2221_out1            : std_logic;
  SIGNAL Logical_Operator_out2222_out1            : std_logic;
  SIGNAL Logical_Operator_out2223_out1            : std_logic;
  SIGNAL Logical_Operator_out2224_out1            : std_logic;
  SIGNAL Logical_Operator_out2225_out1            : std_logic;
  SIGNAL Logical_Operator_out2226_out1            : std_logic;
  SIGNAL Logical_Operator_out2227_out1            : std_logic;
  SIGNAL Logical_Operator_out2228_out1            : std_logic;
  SIGNAL Logical_Operator_out2229_out1            : std_logic;
  SIGNAL Logical_Operator_out2230_out1            : std_logic;
  SIGNAL Logical_Operator_out2231_out1            : std_logic;
  SIGNAL Logical_Operator_out2232_out1            : std_logic;
  SIGNAL Logical_Operator_out2233_out1            : std_logic;
  SIGNAL Logical_Operator_out2234_out1            : std_logic;
  SIGNAL Logical_Operator_out2235_out1            : std_logic;
  SIGNAL Logical_Operator_out2236_out1            : std_logic;
  SIGNAL Logical_Operator_out2237_out1            : std_logic;
  SIGNAL Logical_Operator_out2238_out1            : std_logic;
  SIGNAL Logical_Operator_out2239_out1            : std_logic;
  SIGNAL Logical_Operator_out2240_out1            : std_logic;
  SIGNAL Logical_Operator_out2241_out1            : std_logic;
  SIGNAL Logical_Operator_out2242_out1            : std_logic;
  SIGNAL Logical_Operator_out2243_out1            : std_logic;
  SIGNAL Logical_Operator_out2244_out1            : std_logic;
  SIGNAL Logical_Operator_out2245_out1            : std_logic;
  SIGNAL Logical_Operator_out2246_out1            : std_logic;
  SIGNAL Logical_Operator_out2247_out1            : std_logic;
  SIGNAL Logical_Operator_out2248_out1            : std_logic;
  SIGNAL Logical_Operator_out2249_out1            : std_logic;
  SIGNAL Logical_Operator_out2250_out1            : std_logic;
  SIGNAL Logical_Operator_out2251_out1            : std_logic;
  SIGNAL Logical_Operator_out2252_out1            : std_logic;
  SIGNAL Logical_Operator_out2253_out1            : std_logic;
  SIGNAL Logical_Operator_out2254_out1            : std_logic;
  SIGNAL Logical_Operator_out2255_out1            : std_logic;
  SIGNAL Logical_Operator_out2256_out1            : std_logic;
  SIGNAL Logical_Operator_out2257_out1            : std_logic;
  SIGNAL Logical_Operator_out2258_out1            : std_logic;
  SIGNAL Logical_Operator_out2259_out1            : std_logic;
  SIGNAL Logical_Operator_out2260_out1            : std_logic;
  SIGNAL Logical_Operator_out2261_out1            : std_logic;
  SIGNAL Logical_Operator_out2262_out1            : std_logic;
  SIGNAL Logical_Operator_out2263_out1            : std_logic;
  SIGNAL Logical_Operator_out2264_out1            : std_logic;
  SIGNAL Logical_Operator_out2265_out1            : std_logic;
  SIGNAL Logical_Operator_out2266_out1            : std_logic;
  SIGNAL Logical_Operator_out2267_out1            : std_logic;
  SIGNAL Logical_Operator_out2268_out1            : std_logic;
  SIGNAL Logical_Operator_out2269_out1            : std_logic;
  SIGNAL Logical_Operator_out2270_out1            : std_logic;
  SIGNAL Logical_Operator_out2271_out1            : std_logic;
  SIGNAL Logical_Operator_out2272_out1            : std_logic;
  SIGNAL Logical_Operator_out2273_out1            : std_logic;
  SIGNAL Logical_Operator_out2274_out1            : std_logic;
  SIGNAL Logical_Operator_out2275_out1            : std_logic;
  SIGNAL Logical_Operator_out2276_out1            : std_logic;
  SIGNAL Logical_Operator_out2277_out1            : std_logic;
  SIGNAL Logical_Operator_out2278_out1            : std_logic;
  SIGNAL Logical_Operator_out2279_out1            : std_logic;
  SIGNAL Logical_Operator_out2280_out1            : std_logic;
  SIGNAL Logical_Operator_out2281_out1            : std_logic;
  SIGNAL Logical_Operator_out2282_out1            : std_logic;
  SIGNAL Logical_Operator_out2283_out1            : std_logic;
  SIGNAL Logical_Operator_out2284_out1            : std_logic;
  SIGNAL Logical_Operator_out2285_out1            : std_logic;
  SIGNAL Logical_Operator_out2286_out1            : std_logic;
  SIGNAL Logical_Operator_out2287_out1            : std_logic;
  SIGNAL Logical_Operator_out2288_out1            : std_logic;
  SIGNAL Logical_Operator_out2289_out1            : std_logic;
  SIGNAL Logical_Operator_out2290_out1            : std_logic;
  SIGNAL Logical_Operator_out2291_out1            : std_logic;
  SIGNAL Logical_Operator_out2292_out1            : std_logic;
  SIGNAL Logical_Operator_out2293_out1            : std_logic;
  SIGNAL Logical_Operator_out2294_out1            : std_logic;
  SIGNAL Logical_Operator_out2295_out1            : std_logic;
  SIGNAL Logical_Operator_out2296_out1            : std_logic;
  SIGNAL Logical_Operator_out2297_out1            : std_logic;
  SIGNAL Logical_Operator_out2298_out1            : std_logic;
  SIGNAL Logical_Operator_out2299_out1            : std_logic;
  SIGNAL Logical_Operator_out2300_out1            : std_logic;
  SIGNAL Logical_Operator_out2301_out1            : std_logic;
  SIGNAL Logical_Operator_out2302_out1            : std_logic;
  SIGNAL Logical_Operator_out2303_out1            : std_logic;
  SIGNAL Logical_Operator_out2304_out1            : std_logic;

BEGIN

  Logical_Operator_out1_out1 <= in1 XOR in2;

  Logical_Operator_out2_out1 <= in3 XOR in4;

  Logical_Operator_out3_out1 <= in5 XOR in6;

  Logical_Operator_out4_out1 <= in7 XOR in8;

  Logical_Operator_out5_out1 <= in9 XOR in10;

  Logical_Operator_out6_out1 <= in11 XOR in12;

  Logical_Operator_out7_out1 <= in13 XOR in14;

  Logical_Operator_out8_out1 <= in15 XOR in16;

  Logical_Operator_out9_out1 <= in17 XOR in18;

  Logical_Operator_out10_out1 <= in19 XOR in20;

  Logical_Operator_out11_out1 <= in21 XOR in22;

  Logical_Operator_out12_out1 <= in23 XOR in24;

  Logical_Operator_out13_out1 <= in25 XOR in26;

  Logical_Operator_out14_out1 <= in27 XOR in28;

  Logical_Operator_out15_out1 <= in29 XOR in30;

  Logical_Operator_out16_out1 <= in31 XOR in32;

  Logical_Operator_out17_out1 <= in33 XOR in34;

  Logical_Operator_out18_out1 <= in35 XOR in36;

  Logical_Operator_out19_out1 <= in37 XOR in38;

  Logical_Operator_out20_out1 <= in39 XOR in40;

  Logical_Operator_out21_out1 <= in41 XOR in42;

  Logical_Operator_out22_out1 <= in43 XOR in44;

  Logical_Operator_out23_out1 <= in45 XOR in46;

  Logical_Operator_out24_out1 <= in47 XOR in48;

  Logical_Operator_out25_out1 <= in49 XOR in50;

  Logical_Operator_out26_out1 <= in51 XOR in52;

  Logical_Operator_out27_out1 <= in53 XOR in54;

  Logical_Operator_out28_out1 <= in55 XOR in56;

  Logical_Operator_out29_out1 <= in57 XOR in58;

  Logical_Operator_out30_out1 <= in59 XOR in60;

  Logical_Operator_out31_out1 <= in61 XOR in62;

  Logical_Operator_out32_out1 <= in63 XOR in64;

  Logical_Operator_out33_out1 <= in65 XOR in66;

  Logical_Operator_out34_out1 <= in67 XOR in68;

  Logical_Operator_out35_out1 <= in69 XOR in70;

  Logical_Operator_out36_out1 <= in71 XOR in72;

  Logical_Operator_out37_out1 <= in73 XOR in74;

  Logical_Operator_out38_out1 <= in75 XOR in76;

  Logical_Operator_out39_out1 <= in77 XOR in78;

  Logical_Operator_out40_out1 <= in79 XOR in80;

  Logical_Operator_out41_out1 <= in81 XOR in82;

  Logical_Operator_out42_out1 <= in83 XOR in84;

  Logical_Operator_out43_out1 <= in85 XOR in86;

  Logical_Operator_out44_out1 <= in87 XOR in88;

  Logical_Operator_out45_out1 <= in89 XOR in90;

  Logical_Operator_out46_out1 <= in91 XOR in92;

  Logical_Operator_out47_out1 <= in93 XOR in94;

  Logical_Operator_out48_out1 <= in95 XOR in96;

  Logical_Operator_out49_out1 <= in97 XOR in98;

  Logical_Operator_out50_out1 <= in99 XOR in100;

  Logical_Operator_out51_out1 <= in101 XOR in102;

  Logical_Operator_out52_out1 <= in103 XOR in104;

  Logical_Operator_out53_out1 <= in105 XOR in106;

  Logical_Operator_out54_out1 <= in107 XOR in108;

  Logical_Operator_out55_out1 <= in109 XOR in110;

  Logical_Operator_out56_out1 <= in111 XOR in112;

  Logical_Operator_out57_out1 <= in113 XOR in114;

  Logical_Operator_out58_out1 <= in115 XOR in116;

  Logical_Operator_out59_out1 <= in117 XOR in118;

  Logical_Operator_out60_out1 <= in119 XOR in120;

  Logical_Operator_out61_out1 <= in121 XOR in122;

  Logical_Operator_out62_out1 <= in123 XOR in124;

  Logical_Operator_out63_out1 <= in125 XOR in126;

  Logical_Operator_out64_out1 <= in127 XOR in128;

  Logical_Operator_out65_out1 <= in129 XOR in130;

  Logical_Operator_out66_out1 <= in131 XOR in132;

  Logical_Operator_out67_out1 <= in133 XOR in134;

  Logical_Operator_out68_out1 <= in135 XOR in136;

  Logical_Operator_out69_out1 <= in137 XOR in138;

  Logical_Operator_out70_out1 <= in139 XOR in140;

  Logical_Operator_out71_out1 <= in141 XOR in142;

  Logical_Operator_out72_out1 <= in143 XOR in144;

  Logical_Operator_out73_out1 <= in145 XOR in146;

  Logical_Operator_out74_out1 <= in147 XOR in148;

  Logical_Operator_out75_out1 <= in149 XOR in150;

  Logical_Operator_out76_out1 <= in151 XOR in152;

  Logical_Operator_out77_out1 <= in153 XOR in154;

  Logical_Operator_out78_out1 <= in155 XOR in156;

  Logical_Operator_out79_out1 <= in157 XOR in158;

  Logical_Operator_out80_out1 <= in159 XOR in160;

  Logical_Operator_out81_out1 <= in161 XOR in162;

  Logical_Operator_out82_out1 <= in163 XOR in164;

  Logical_Operator_out83_out1 <= in165 XOR in166;

  Logical_Operator_out84_out1 <= in167 XOR in168;

  Logical_Operator_out85_out1 <= in169 XOR in170;

  Logical_Operator_out86_out1 <= in171 XOR in172;

  Logical_Operator_out87_out1 <= in173 XOR in174;

  Logical_Operator_out88_out1 <= in175 XOR in176;

  Logical_Operator_out89_out1 <= in177 XOR in178;

  Logical_Operator_out90_out1 <= in179 XOR in180;

  Logical_Operator_out91_out1 <= in181 XOR in182;

  Logical_Operator_out92_out1 <= in183 XOR in184;

  Logical_Operator_out93_out1 <= in185 XOR in186;

  Logical_Operator_out94_out1 <= in187 XOR in188;

  Logical_Operator_out95_out1 <= in189 XOR in190;

  Logical_Operator_out96_out1 <= in191 XOR in192;

  Logical_Operator_out97_out1 <= in193 XOR in194;

  Logical_Operator_out98_out1 <= in195 XOR in196;

  Logical_Operator_out99_out1 <= in197 XOR in198;

  Logical_Operator_out100_out1 <= in199 XOR in200;

  Logical_Operator_out101_out1 <= in201 XOR in202;

  Logical_Operator_out102_out1 <= in203 XOR in204;

  Logical_Operator_out103_out1 <= in205 XOR in206;

  Logical_Operator_out104_out1 <= in207 XOR in208;

  Logical_Operator_out105_out1 <= in209 XOR in210;

  Logical_Operator_out106_out1 <= in211 XOR in212;

  Logical_Operator_out107_out1 <= in213 XOR in214;

  Logical_Operator_out108_out1 <= in215 XOR in216;

  Logical_Operator_out109_out1 <= in217 XOR in218;

  Logical_Operator_out110_out1 <= in219 XOR in220;

  Logical_Operator_out111_out1 <= in221 XOR in222;

  Logical_Operator_out112_out1 <= in223 XOR in224;

  Logical_Operator_out113_out1 <= in225 XOR in226;

  Logical_Operator_out114_out1 <= in227 XOR in228;

  Logical_Operator_out115_out1 <= in229 XOR in230;

  Logical_Operator_out116_out1 <= in231 XOR in232;

  Logical_Operator_out117_out1 <= in233 XOR in234;

  Logical_Operator_out118_out1 <= in235 XOR in236;

  Logical_Operator_out119_out1 <= in237 XOR in238;

  Logical_Operator_out120_out1 <= in239 XOR in240;

  Logical_Operator_out121_out1 <= in241 XOR in242;

  Logical_Operator_out122_out1 <= in243 XOR in244;

  Logical_Operator_out123_out1 <= in245 XOR in246;

  Logical_Operator_out124_out1 <= in247 XOR in248;

  Logical_Operator_out125_out1 <= in249 XOR in250;

  Logical_Operator_out126_out1 <= in251 XOR in252;

  Logical_Operator_out127_out1 <= in253 XOR in254;

  Logical_Operator_out128_out1 <= in255 XOR in256;

  Logical_Operator_out129_out1 <= in257 XOR in258;

  Logical_Operator_out130_out1 <= in259 XOR in260;

  Logical_Operator_out131_out1 <= in261 XOR in262;

  Logical_Operator_out132_out1 <= in263 XOR in264;

  Logical_Operator_out133_out1 <= in265 XOR in266;

  Logical_Operator_out134_out1 <= in267 XOR in268;

  Logical_Operator_out135_out1 <= in269 XOR in270;

  Logical_Operator_out136_out1 <= in271 XOR in272;

  Logical_Operator_out137_out1 <= in273 XOR in274;

  Logical_Operator_out138_out1 <= in275 XOR in276;

  Logical_Operator_out139_out1 <= in277 XOR in278;

  Logical_Operator_out140_out1 <= in279 XOR in280;

  Logical_Operator_out141_out1 <= in281 XOR in282;

  Logical_Operator_out142_out1 <= in283 XOR in284;

  Logical_Operator_out143_out1 <= in285 XOR in286;

  Logical_Operator_out144_out1 <= in287 XOR in288;

  Logical_Operator_out145_out1 <= in289 XOR in290;

  Logical_Operator_out146_out1 <= in291 XOR in292;

  Logical_Operator_out147_out1 <= in293 XOR in294;

  Logical_Operator_out148_out1 <= in295 XOR in296;

  Logical_Operator_out149_out1 <= in297 XOR in298;

  Logical_Operator_out150_out1 <= in299 XOR in300;

  Logical_Operator_out151_out1 <= in301 XOR in302;

  Logical_Operator_out152_out1 <= in303 XOR in304;

  Logical_Operator_out153_out1 <= in305 XOR in306;

  Logical_Operator_out154_out1 <= in307 XOR in308;

  Logical_Operator_out155_out1 <= in309 XOR in310;

  Logical_Operator_out156_out1 <= in311 XOR in312;

  Logical_Operator_out157_out1 <= in313 XOR in314;

  Logical_Operator_out158_out1 <= in315 XOR in316;

  Logical_Operator_out159_out1 <= in317 XOR in318;

  Logical_Operator_out160_out1 <= in319 XOR in320;

  Logical_Operator_out161_out1 <= in321 XOR in322;

  Logical_Operator_out162_out1 <= in323 XOR in324;

  Logical_Operator_out163_out1 <= in325 XOR in326;

  Logical_Operator_out164_out1 <= in327 XOR in328;

  Logical_Operator_out165_out1 <= in329 XOR in330;

  Logical_Operator_out166_out1 <= in331 XOR in332;

  Logical_Operator_out167_out1 <= in333 XOR in334;

  Logical_Operator_out168_out1 <= in335 XOR in336;

  Logical_Operator_out169_out1 <= in337 XOR in338;

  Logical_Operator_out170_out1 <= in339 XOR in340;

  Logical_Operator_out171_out1 <= in341 XOR in342;

  Logical_Operator_out172_out1 <= in343 XOR in344;

  Logical_Operator_out173_out1 <= in345 XOR in346;

  Logical_Operator_out174_out1 <= in347 XOR in348;

  Logical_Operator_out175_out1 <= in349 XOR in350;

  Logical_Operator_out176_out1 <= in351 XOR in352;

  Logical_Operator_out177_out1 <= in353 XOR in354;

  Logical_Operator_out178_out1 <= in355 XOR in356;

  Logical_Operator_out179_out1 <= in357 XOR in358;

  Logical_Operator_out180_out1 <= in359 XOR in360;

  Logical_Operator_out181_out1 <= in361 XOR in362;

  Logical_Operator_out182_out1 <= in363 XOR in364;

  Logical_Operator_out183_out1 <= in365 XOR in366;

  Logical_Operator_out184_out1 <= in367 XOR in368;

  Logical_Operator_out185_out1 <= in369 XOR in370;

  Logical_Operator_out186_out1 <= in371 XOR in372;

  Logical_Operator_out187_out1 <= in373 XOR in374;

  Logical_Operator_out188_out1 <= in375 XOR in376;

  Logical_Operator_out189_out1 <= in377 XOR in378;

  Logical_Operator_out190_out1 <= in379 XOR in380;

  Logical_Operator_out191_out1 <= in381 XOR in382;

  Logical_Operator_out192_out1 <= in383 XOR in384;

  Logical_Operator_out193_out1 <= in385 XOR in386;

  Logical_Operator_out194_out1 <= in387 XOR in388;

  Logical_Operator_out195_out1 <= in389 XOR in390;

  Logical_Operator_out196_out1 <= in391 XOR in392;

  Logical_Operator_out197_out1 <= in393 XOR in394;

  Logical_Operator_out198_out1 <= in395 XOR in396;

  Logical_Operator_out199_out1 <= in397 XOR in398;

  Logical_Operator_out200_out1 <= in399 XOR in400;

  Logical_Operator_out201_out1 <= in401 XOR in402;

  Logical_Operator_out202_out1 <= in403 XOR in404;

  Logical_Operator_out203_out1 <= in405 XOR in406;

  Logical_Operator_out204_out1 <= in407 XOR in408;

  Logical_Operator_out205_out1 <= in409 XOR in410;

  Logical_Operator_out206_out1 <= in411 XOR in412;

  Logical_Operator_out207_out1 <= in413 XOR in414;

  Logical_Operator_out208_out1 <= in415 XOR in416;

  Logical_Operator_out209_out1 <= in417 XOR in418;

  Logical_Operator_out210_out1 <= in419 XOR in420;

  Logical_Operator_out211_out1 <= in421 XOR in422;

  Logical_Operator_out212_out1 <= in423 XOR in424;

  Logical_Operator_out213_out1 <= in425 XOR in426;

  Logical_Operator_out214_out1 <= in427 XOR in428;

  Logical_Operator_out215_out1 <= in429 XOR in430;

  Logical_Operator_out216_out1 <= in431 XOR in432;

  Logical_Operator_out217_out1 <= in433 XOR in434;

  Logical_Operator_out218_out1 <= in435 XOR in436;

  Logical_Operator_out219_out1 <= in437 XOR in438;

  Logical_Operator_out220_out1 <= in439 XOR in440;

  Logical_Operator_out221_out1 <= in441 XOR in442;

  Logical_Operator_out222_out1 <= in443 XOR in444;

  Logical_Operator_out223_out1 <= in445 XOR in446;

  Logical_Operator_out224_out1 <= in447 XOR in448;

  Logical_Operator_out225_out1 <= in449 XOR in450;

  Logical_Operator_out226_out1 <= in451 XOR in452;

  Logical_Operator_out227_out1 <= in453 XOR in454;

  Logical_Operator_out228_out1 <= in455 XOR in456;

  Logical_Operator_out229_out1 <= in457 XOR in458;

  Logical_Operator_out230_out1 <= in459 XOR in460;

  Logical_Operator_out231_out1 <= in461 XOR in462;

  Logical_Operator_out232_out1 <= in463 XOR in464;

  Logical_Operator_out233_out1 <= in465 XOR in466;

  Logical_Operator_out234_out1 <= in467 XOR in468;

  Logical_Operator_out235_out1 <= in469 XOR in470;

  Logical_Operator_out236_out1 <= in471 XOR in472;

  Logical_Operator_out237_out1 <= in473 XOR in474;

  Logical_Operator_out238_out1 <= in475 XOR in476;

  Logical_Operator_out239_out1 <= in477 XOR in478;

  Logical_Operator_out240_out1 <= in479 XOR in480;

  Logical_Operator_out241_out1 <= in481 XOR in482;

  Logical_Operator_out242_out1 <= in483 XOR in484;

  Logical_Operator_out243_out1 <= in485 XOR in486;

  Logical_Operator_out244_out1 <= in487 XOR in488;

  Logical_Operator_out245_out1 <= in489 XOR in490;

  Logical_Operator_out246_out1 <= in491 XOR in492;

  Logical_Operator_out247_out1 <= in493 XOR in494;

  Logical_Operator_out248_out1 <= in495 XOR in496;

  Logical_Operator_out249_out1 <= in497 XOR in498;

  Logical_Operator_out250_out1 <= in499 XOR in500;

  Logical_Operator_out251_out1 <= in501 XOR in502;

  Logical_Operator_out252_out1 <= in503 XOR in504;

  Logical_Operator_out253_out1 <= in505 XOR in506;

  Logical_Operator_out254_out1 <= in507 XOR in508;

  Logical_Operator_out255_out1 <= in509 XOR in510;

  Logical_Operator_out256_out1 <= in511 XOR in512;

  Logical_Operator_out257_out1 <= Logical_Operator_out1_out1 XOR Logical_Operator_out2_out1;

  Logical_Operator_out258_out1 <= in2 XOR in4;

  Logical_Operator_out259_out1 <= Logical_Operator_out3_out1 XOR Logical_Operator_out4_out1;

  Logical_Operator_out260_out1 <= in6 XOR in8;

  Logical_Operator_out261_out1 <= Logical_Operator_out5_out1 XOR Logical_Operator_out6_out1;

  Logical_Operator_out262_out1 <= in10 XOR in12;

  Logical_Operator_out263_out1 <= Logical_Operator_out7_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out264_out1 <= in14 XOR in16;

  Logical_Operator_out265_out1 <= Logical_Operator_out9_out1 XOR Logical_Operator_out10_out1;

  Logical_Operator_out266_out1 <= in18 XOR in20;

  Logical_Operator_out267_out1 <= Logical_Operator_out11_out1 XOR Logical_Operator_out12_out1;

  Logical_Operator_out268_out1 <= in22 XOR in24;

  Logical_Operator_out269_out1 <= Logical_Operator_out13_out1 XOR Logical_Operator_out14_out1;

  Logical_Operator_out270_out1 <= in26 XOR in28;

  Logical_Operator_out271_out1 <= Logical_Operator_out15_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out272_out1 <= in30 XOR in32;

  Logical_Operator_out273_out1 <= Logical_Operator_out17_out1 XOR Logical_Operator_out18_out1;

  Logical_Operator_out274_out1 <= in34 XOR in36;

  Logical_Operator_out275_out1 <= Logical_Operator_out19_out1 XOR Logical_Operator_out20_out1;

  Logical_Operator_out276_out1 <= in38 XOR in40;

  Logical_Operator_out277_out1 <= Logical_Operator_out21_out1 XOR Logical_Operator_out22_out1;

  Logical_Operator_out278_out1 <= in42 XOR in44;

  Logical_Operator_out279_out1 <= Logical_Operator_out23_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out280_out1 <= in46 XOR in48;

  Logical_Operator_out281_out1 <= Logical_Operator_out25_out1 XOR Logical_Operator_out26_out1;

  Logical_Operator_out282_out1 <= in50 XOR in52;

  Logical_Operator_out283_out1 <= Logical_Operator_out27_out1 XOR Logical_Operator_out28_out1;

  Logical_Operator_out284_out1 <= in54 XOR in56;

  Logical_Operator_out285_out1 <= Logical_Operator_out29_out1 XOR Logical_Operator_out30_out1;

  Logical_Operator_out286_out1 <= in58 XOR in60;

  Logical_Operator_out287_out1 <= Logical_Operator_out31_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out288_out1 <= in62 XOR in64;

  Logical_Operator_out289_out1 <= Logical_Operator_out33_out1 XOR Logical_Operator_out34_out1;

  Logical_Operator_out290_out1 <= in66 XOR in68;

  Logical_Operator_out291_out1 <= Logical_Operator_out35_out1 XOR Logical_Operator_out36_out1;

  Logical_Operator_out292_out1 <= in70 XOR in72;

  Logical_Operator_out293_out1 <= Logical_Operator_out37_out1 XOR Logical_Operator_out38_out1;

  Logical_Operator_out294_out1 <= in74 XOR in76;

  Logical_Operator_out295_out1 <= Logical_Operator_out39_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out296_out1 <= in78 XOR in80;

  Logical_Operator_out297_out1 <= Logical_Operator_out41_out1 XOR Logical_Operator_out42_out1;

  Logical_Operator_out298_out1 <= in82 XOR in84;

  Logical_Operator_out299_out1 <= Logical_Operator_out43_out1 XOR Logical_Operator_out44_out1;

  Logical_Operator_out300_out1 <= in86 XOR in88;

  Logical_Operator_out301_out1 <= Logical_Operator_out45_out1 XOR Logical_Operator_out46_out1;

  Logical_Operator_out302_out1 <= in90 XOR in92;

  Logical_Operator_out303_out1 <= Logical_Operator_out47_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out304_out1 <= in94 XOR in96;

  Logical_Operator_out305_out1 <= Logical_Operator_out49_out1 XOR Logical_Operator_out50_out1;

  Logical_Operator_out306_out1 <= in98 XOR in100;

  Logical_Operator_out307_out1 <= Logical_Operator_out51_out1 XOR Logical_Operator_out52_out1;

  Logical_Operator_out308_out1 <= in102 XOR in104;

  Logical_Operator_out309_out1 <= Logical_Operator_out53_out1 XOR Logical_Operator_out54_out1;

  Logical_Operator_out310_out1 <= in106 XOR in108;

  Logical_Operator_out311_out1 <= Logical_Operator_out55_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out312_out1 <= in110 XOR in112;

  Logical_Operator_out313_out1 <= Logical_Operator_out57_out1 XOR Logical_Operator_out58_out1;

  Logical_Operator_out314_out1 <= in114 XOR in116;

  Logical_Operator_out315_out1 <= Logical_Operator_out59_out1 XOR Logical_Operator_out60_out1;

  Logical_Operator_out316_out1 <= in118 XOR in120;

  Logical_Operator_out317_out1 <= Logical_Operator_out61_out1 XOR Logical_Operator_out62_out1;

  Logical_Operator_out318_out1 <= in122 XOR in124;

  Logical_Operator_out319_out1 <= Logical_Operator_out63_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out320_out1 <= in126 XOR in128;

  Logical_Operator_out321_out1 <= Logical_Operator_out65_out1 XOR Logical_Operator_out66_out1;

  Logical_Operator_out322_out1 <= in130 XOR in132;

  Logical_Operator_out323_out1 <= Logical_Operator_out67_out1 XOR Logical_Operator_out68_out1;

  Logical_Operator_out324_out1 <= in134 XOR in136;

  Logical_Operator_out325_out1 <= Logical_Operator_out69_out1 XOR Logical_Operator_out70_out1;

  Logical_Operator_out326_out1 <= in138 XOR in140;

  Logical_Operator_out327_out1 <= Logical_Operator_out71_out1 XOR Logical_Operator_out72_out1;

  Logical_Operator_out328_out1 <= in142 XOR in144;

  Logical_Operator_out329_out1 <= Logical_Operator_out73_out1 XOR Logical_Operator_out74_out1;

  Logical_Operator_out330_out1 <= in146 XOR in148;

  Logical_Operator_out331_out1 <= Logical_Operator_out75_out1 XOR Logical_Operator_out76_out1;

  Logical_Operator_out332_out1 <= in150 XOR in152;

  Logical_Operator_out333_out1 <= Logical_Operator_out77_out1 XOR Logical_Operator_out78_out1;

  Logical_Operator_out334_out1 <= in154 XOR in156;

  Logical_Operator_out335_out1 <= Logical_Operator_out79_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out336_out1 <= in158 XOR in160;

  Logical_Operator_out337_out1 <= Logical_Operator_out81_out1 XOR Logical_Operator_out82_out1;

  Logical_Operator_out338_out1 <= in162 XOR in164;

  Logical_Operator_out339_out1 <= Logical_Operator_out83_out1 XOR Logical_Operator_out84_out1;

  Logical_Operator_out340_out1 <= in166 XOR in168;

  Logical_Operator_out341_out1 <= Logical_Operator_out85_out1 XOR Logical_Operator_out86_out1;

  Logical_Operator_out342_out1 <= in170 XOR in172;

  Logical_Operator_out343_out1 <= Logical_Operator_out87_out1 XOR Logical_Operator_out88_out1;

  Logical_Operator_out344_out1 <= in174 XOR in176;

  Logical_Operator_out345_out1 <= Logical_Operator_out89_out1 XOR Logical_Operator_out90_out1;

  Logical_Operator_out346_out1 <= in178 XOR in180;

  Logical_Operator_out347_out1 <= Logical_Operator_out91_out1 XOR Logical_Operator_out92_out1;

  Logical_Operator_out348_out1 <= in182 XOR in184;

  Logical_Operator_out349_out1 <= Logical_Operator_out93_out1 XOR Logical_Operator_out94_out1;

  Logical_Operator_out350_out1 <= in186 XOR in188;

  Logical_Operator_out351_out1 <= Logical_Operator_out95_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out352_out1 <= in190 XOR in192;

  Logical_Operator_out353_out1 <= Logical_Operator_out97_out1 XOR Logical_Operator_out98_out1;

  Logical_Operator_out354_out1 <= in194 XOR in196;

  Logical_Operator_out355_out1 <= Logical_Operator_out99_out1 XOR Logical_Operator_out100_out1;

  Logical_Operator_out356_out1 <= in198 XOR in200;

  Logical_Operator_out357_out1 <= Logical_Operator_out101_out1 XOR Logical_Operator_out102_out1;

  Logical_Operator_out358_out1 <= in202 XOR in204;

  Logical_Operator_out359_out1 <= Logical_Operator_out103_out1 XOR Logical_Operator_out104_out1;

  Logical_Operator_out360_out1 <= in206 XOR in208;

  Logical_Operator_out361_out1 <= Logical_Operator_out105_out1 XOR Logical_Operator_out106_out1;

  Logical_Operator_out362_out1 <= in210 XOR in212;

  Logical_Operator_out363_out1 <= Logical_Operator_out107_out1 XOR Logical_Operator_out108_out1;

  Logical_Operator_out364_out1 <= in214 XOR in216;

  Logical_Operator_out365_out1 <= Logical_Operator_out109_out1 XOR Logical_Operator_out110_out1;

  Logical_Operator_out366_out1 <= in218 XOR in220;

  Logical_Operator_out367_out1 <= Logical_Operator_out111_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out368_out1 <= in222 XOR in224;

  Logical_Operator_out369_out1 <= Logical_Operator_out113_out1 XOR Logical_Operator_out114_out1;

  Logical_Operator_out370_out1 <= in226 XOR in228;

  Logical_Operator_out371_out1 <= Logical_Operator_out115_out1 XOR Logical_Operator_out116_out1;

  Logical_Operator_out372_out1 <= in230 XOR in232;

  Logical_Operator_out373_out1 <= Logical_Operator_out117_out1 XOR Logical_Operator_out118_out1;

  Logical_Operator_out374_out1 <= in234 XOR in236;

  Logical_Operator_out375_out1 <= Logical_Operator_out119_out1 XOR Logical_Operator_out120_out1;

  Logical_Operator_out376_out1 <= in238 XOR in240;

  Logical_Operator_out377_out1 <= Logical_Operator_out121_out1 XOR Logical_Operator_out122_out1;

  Logical_Operator_out378_out1 <= in242 XOR in244;

  Logical_Operator_out379_out1 <= Logical_Operator_out123_out1 XOR Logical_Operator_out124_out1;

  Logical_Operator_out380_out1 <= in246 XOR in248;

  Logical_Operator_out381_out1 <= Logical_Operator_out125_out1 XOR Logical_Operator_out126_out1;

  Logical_Operator_out382_out1 <= in250 XOR in252;

  Logical_Operator_out383_out1 <= Logical_Operator_out127_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out384_out1 <= in254 XOR in256;

  Logical_Operator_out385_out1 <= Logical_Operator_out129_out1 XOR Logical_Operator_out130_out1;

  Logical_Operator_out386_out1 <= in258 XOR in260;

  Logical_Operator_out387_out1 <= Logical_Operator_out131_out1 XOR Logical_Operator_out132_out1;

  Logical_Operator_out388_out1 <= in262 XOR in264;

  Logical_Operator_out389_out1 <= Logical_Operator_out133_out1 XOR Logical_Operator_out134_out1;

  Logical_Operator_out390_out1 <= in266 XOR in268;

  Logical_Operator_out391_out1 <= Logical_Operator_out135_out1 XOR Logical_Operator_out136_out1;

  Logical_Operator_out392_out1 <= in270 XOR in272;

  Logical_Operator_out393_out1 <= Logical_Operator_out137_out1 XOR Logical_Operator_out138_out1;

  Logical_Operator_out394_out1 <= in274 XOR in276;

  Logical_Operator_out395_out1 <= Logical_Operator_out139_out1 XOR Logical_Operator_out140_out1;

  Logical_Operator_out396_out1 <= in278 XOR in280;

  Logical_Operator_out397_out1 <= Logical_Operator_out141_out1 XOR Logical_Operator_out142_out1;

  Logical_Operator_out398_out1 <= in282 XOR in284;

  Logical_Operator_out399_out1 <= Logical_Operator_out143_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out400_out1 <= in286 XOR in288;

  Logical_Operator_out401_out1 <= Logical_Operator_out145_out1 XOR Logical_Operator_out146_out1;

  Logical_Operator_out402_out1 <= in290 XOR in292;

  Logical_Operator_out403_out1 <= Logical_Operator_out147_out1 XOR Logical_Operator_out148_out1;

  Logical_Operator_out404_out1 <= in294 XOR in296;

  Logical_Operator_out405_out1 <= Logical_Operator_out149_out1 XOR Logical_Operator_out150_out1;

  Logical_Operator_out406_out1 <= in298 XOR in300;

  Logical_Operator_out407_out1 <= Logical_Operator_out151_out1 XOR Logical_Operator_out152_out1;

  Logical_Operator_out408_out1 <= in302 XOR in304;

  Logical_Operator_out409_out1 <= Logical_Operator_out153_out1 XOR Logical_Operator_out154_out1;

  Logical_Operator_out410_out1 <= in306 XOR in308;

  Logical_Operator_out411_out1 <= Logical_Operator_out155_out1 XOR Logical_Operator_out156_out1;

  Logical_Operator_out412_out1 <= in310 XOR in312;

  Logical_Operator_out413_out1 <= Logical_Operator_out157_out1 XOR Logical_Operator_out158_out1;

  Logical_Operator_out414_out1 <= in314 XOR in316;

  Logical_Operator_out415_out1 <= Logical_Operator_out159_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out416_out1 <= in318 XOR in320;

  Logical_Operator_out417_out1 <= Logical_Operator_out161_out1 XOR Logical_Operator_out162_out1;

  Logical_Operator_out418_out1 <= in322 XOR in324;

  Logical_Operator_out419_out1 <= Logical_Operator_out163_out1 XOR Logical_Operator_out164_out1;

  Logical_Operator_out420_out1 <= in326 XOR in328;

  Logical_Operator_out421_out1 <= Logical_Operator_out165_out1 XOR Logical_Operator_out166_out1;

  Logical_Operator_out422_out1 <= in330 XOR in332;

  Logical_Operator_out423_out1 <= Logical_Operator_out167_out1 XOR Logical_Operator_out168_out1;

  Logical_Operator_out424_out1 <= in334 XOR in336;

  Logical_Operator_out425_out1 <= Logical_Operator_out169_out1 XOR Logical_Operator_out170_out1;

  Logical_Operator_out426_out1 <= in338 XOR in340;

  Logical_Operator_out427_out1 <= Logical_Operator_out171_out1 XOR Logical_Operator_out172_out1;

  Logical_Operator_out428_out1 <= in342 XOR in344;

  Logical_Operator_out429_out1 <= Logical_Operator_out173_out1 XOR Logical_Operator_out174_out1;

  Logical_Operator_out430_out1 <= in346 XOR in348;

  Logical_Operator_out431_out1 <= Logical_Operator_out175_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out432_out1 <= in350 XOR in352;

  Logical_Operator_out433_out1 <= Logical_Operator_out177_out1 XOR Logical_Operator_out178_out1;

  Logical_Operator_out434_out1 <= in354 XOR in356;

  Logical_Operator_out435_out1 <= Logical_Operator_out179_out1 XOR Logical_Operator_out180_out1;

  Logical_Operator_out436_out1 <= in358 XOR in360;

  Logical_Operator_out437_out1 <= Logical_Operator_out181_out1 XOR Logical_Operator_out182_out1;

  Logical_Operator_out438_out1 <= in362 XOR in364;

  Logical_Operator_out439_out1 <= Logical_Operator_out183_out1 XOR Logical_Operator_out184_out1;

  Logical_Operator_out440_out1 <= in366 XOR in368;

  Logical_Operator_out441_out1 <= Logical_Operator_out185_out1 XOR Logical_Operator_out186_out1;

  Logical_Operator_out442_out1 <= in370 XOR in372;

  Logical_Operator_out443_out1 <= Logical_Operator_out187_out1 XOR Logical_Operator_out188_out1;

  Logical_Operator_out444_out1 <= in374 XOR in376;

  Logical_Operator_out445_out1 <= Logical_Operator_out189_out1 XOR Logical_Operator_out190_out1;

  Logical_Operator_out446_out1 <= in378 XOR in380;

  Logical_Operator_out447_out1 <= Logical_Operator_out191_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out448_out1 <= in382 XOR in384;

  Logical_Operator_out449_out1 <= Logical_Operator_out193_out1 XOR Logical_Operator_out194_out1;

  Logical_Operator_out450_out1 <= in386 XOR in388;

  Logical_Operator_out451_out1 <= Logical_Operator_out195_out1 XOR Logical_Operator_out196_out1;

  Logical_Operator_out452_out1 <= in390 XOR in392;

  Logical_Operator_out453_out1 <= Logical_Operator_out197_out1 XOR Logical_Operator_out198_out1;

  Logical_Operator_out454_out1 <= in394 XOR in396;

  Logical_Operator_out455_out1 <= Logical_Operator_out199_out1 XOR Logical_Operator_out200_out1;

  Logical_Operator_out456_out1 <= in398 XOR in400;

  Logical_Operator_out457_out1 <= Logical_Operator_out201_out1 XOR Logical_Operator_out202_out1;

  Logical_Operator_out458_out1 <= in402 XOR in404;

  Logical_Operator_out459_out1 <= Logical_Operator_out203_out1 XOR Logical_Operator_out204_out1;

  Logical_Operator_out460_out1 <= in406 XOR in408;

  Logical_Operator_out461_out1 <= Logical_Operator_out205_out1 XOR Logical_Operator_out206_out1;

  Logical_Operator_out462_out1 <= in410 XOR in412;

  Logical_Operator_out463_out1 <= Logical_Operator_out207_out1 XOR Logical_Operator_out208_out1;

  Logical_Operator_out464_out1 <= in414 XOR in416;

  Logical_Operator_out465_out1 <= Logical_Operator_out209_out1 XOR Logical_Operator_out210_out1;

  Logical_Operator_out466_out1 <= in418 XOR in420;

  Logical_Operator_out467_out1 <= Logical_Operator_out211_out1 XOR Logical_Operator_out212_out1;

  Logical_Operator_out468_out1 <= in422 XOR in424;

  Logical_Operator_out469_out1 <= Logical_Operator_out213_out1 XOR Logical_Operator_out214_out1;

  Logical_Operator_out470_out1 <= in426 XOR in428;

  Logical_Operator_out471_out1 <= Logical_Operator_out215_out1 XOR Logical_Operator_out216_out1;

  Logical_Operator_out472_out1 <= in430 XOR in432;

  Logical_Operator_out473_out1 <= Logical_Operator_out217_out1 XOR Logical_Operator_out218_out1;

  Logical_Operator_out474_out1 <= in434 XOR in436;

  Logical_Operator_out475_out1 <= Logical_Operator_out219_out1 XOR Logical_Operator_out220_out1;

  Logical_Operator_out476_out1 <= in438 XOR in440;

  Logical_Operator_out477_out1 <= Logical_Operator_out221_out1 XOR Logical_Operator_out222_out1;

  Logical_Operator_out478_out1 <= in442 XOR in444;

  Logical_Operator_out479_out1 <= Logical_Operator_out223_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out480_out1 <= in446 XOR in448;

  Logical_Operator_out481_out1 <= Logical_Operator_out225_out1 XOR Logical_Operator_out226_out1;

  Logical_Operator_out482_out1 <= in450 XOR in452;

  Logical_Operator_out483_out1 <= Logical_Operator_out227_out1 XOR Logical_Operator_out228_out1;

  Logical_Operator_out484_out1 <= in454 XOR in456;

  Logical_Operator_out485_out1 <= Logical_Operator_out229_out1 XOR Logical_Operator_out230_out1;

  Logical_Operator_out486_out1 <= in458 XOR in460;

  Logical_Operator_out487_out1 <= Logical_Operator_out231_out1 XOR Logical_Operator_out232_out1;

  Logical_Operator_out488_out1 <= in462 XOR in464;

  Logical_Operator_out489_out1 <= Logical_Operator_out233_out1 XOR Logical_Operator_out234_out1;

  Logical_Operator_out490_out1 <= in466 XOR in468;

  Logical_Operator_out491_out1 <= Logical_Operator_out235_out1 XOR Logical_Operator_out236_out1;

  Logical_Operator_out492_out1 <= in470 XOR in472;

  Logical_Operator_out493_out1 <= Logical_Operator_out237_out1 XOR Logical_Operator_out238_out1;

  Logical_Operator_out494_out1 <= in474 XOR in476;

  Logical_Operator_out495_out1 <= Logical_Operator_out239_out1 XOR Logical_Operator_out240_out1;

  Logical_Operator_out496_out1 <= in478 XOR in480;

  Logical_Operator_out497_out1 <= Logical_Operator_out241_out1 XOR Logical_Operator_out242_out1;

  Logical_Operator_out498_out1 <= in482 XOR in484;

  Logical_Operator_out499_out1 <= Logical_Operator_out243_out1 XOR Logical_Operator_out244_out1;

  Logical_Operator_out500_out1 <= in486 XOR in488;

  Logical_Operator_out501_out1 <= Logical_Operator_out245_out1 XOR Logical_Operator_out246_out1;

  Logical_Operator_out502_out1 <= in490 XOR in492;

  Logical_Operator_out503_out1 <= Logical_Operator_out247_out1 XOR Logical_Operator_out248_out1;

  Logical_Operator_out504_out1 <= in494 XOR in496;

  Logical_Operator_out505_out1 <= Logical_Operator_out249_out1 XOR Logical_Operator_out250_out1;

  Logical_Operator_out506_out1 <= in498 XOR in500;

  Logical_Operator_out507_out1 <= Logical_Operator_out251_out1 XOR Logical_Operator_out252_out1;

  Logical_Operator_out508_out1 <= in502 XOR in504;

  Logical_Operator_out509_out1 <= Logical_Operator_out253_out1 XOR Logical_Operator_out254_out1;

  Logical_Operator_out510_out1 <= in506 XOR in508;

  Logical_Operator_out511_out1 <= Logical_Operator_out255_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out512_out1 <= in510 XOR in512;

  Logical_Operator_out513_out1 <= Logical_Operator_out257_out1 XOR Logical_Operator_out259_out1;

  Logical_Operator_out514_out1 <= Logical_Operator_out258_out1 XOR Logical_Operator_out260_out1;

  Logical_Operator_out515_out1 <= Logical_Operator_out2_out1 XOR Logical_Operator_out4_out1;

  Logical_Operator_out516_out1 <= in4 XOR in8;

  Logical_Operator_out517_out1 <= Logical_Operator_out261_out1 XOR Logical_Operator_out263_out1;

  Logical_Operator_out518_out1 <= Logical_Operator_out262_out1 XOR Logical_Operator_out264_out1;

  Logical_Operator_out519_out1 <= Logical_Operator_out6_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out520_out1 <= in12 XOR in16;

  Logical_Operator_out521_out1 <= Logical_Operator_out265_out1 XOR Logical_Operator_out267_out1;

  Logical_Operator_out522_out1 <= Logical_Operator_out266_out1 XOR Logical_Operator_out268_out1;

  Logical_Operator_out523_out1 <= Logical_Operator_out10_out1 XOR Logical_Operator_out12_out1;

  Logical_Operator_out524_out1 <= in20 XOR in24;

  Logical_Operator_out525_out1 <= Logical_Operator_out269_out1 XOR Logical_Operator_out271_out1;

  Logical_Operator_out526_out1 <= Logical_Operator_out270_out1 XOR Logical_Operator_out272_out1;

  Logical_Operator_out527_out1 <= Logical_Operator_out14_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out528_out1 <= in28 XOR in32;

  Logical_Operator_out529_out1 <= Logical_Operator_out273_out1 XOR Logical_Operator_out275_out1;

  Logical_Operator_out530_out1 <= Logical_Operator_out274_out1 XOR Logical_Operator_out276_out1;

  Logical_Operator_out531_out1 <= Logical_Operator_out18_out1 XOR Logical_Operator_out20_out1;

  Logical_Operator_out532_out1 <= in36 XOR in40;

  Logical_Operator_out533_out1 <= Logical_Operator_out277_out1 XOR Logical_Operator_out279_out1;

  Logical_Operator_out534_out1 <= Logical_Operator_out278_out1 XOR Logical_Operator_out280_out1;

  Logical_Operator_out535_out1 <= Logical_Operator_out22_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out536_out1 <= in44 XOR in48;

  Logical_Operator_out537_out1 <= Logical_Operator_out281_out1 XOR Logical_Operator_out283_out1;

  Logical_Operator_out538_out1 <= Logical_Operator_out282_out1 XOR Logical_Operator_out284_out1;

  Logical_Operator_out539_out1 <= Logical_Operator_out26_out1 XOR Logical_Operator_out28_out1;

  Logical_Operator_out540_out1 <= in52 XOR in56;

  Logical_Operator_out541_out1 <= Logical_Operator_out285_out1 XOR Logical_Operator_out287_out1;

  Logical_Operator_out542_out1 <= Logical_Operator_out286_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out543_out1 <= Logical_Operator_out30_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out544_out1 <= in60 XOR in64;

  Logical_Operator_out545_out1 <= Logical_Operator_out289_out1 XOR Logical_Operator_out291_out1;

  Logical_Operator_out546_out1 <= Logical_Operator_out290_out1 XOR Logical_Operator_out292_out1;

  Logical_Operator_out547_out1 <= Logical_Operator_out34_out1 XOR Logical_Operator_out36_out1;

  Logical_Operator_out548_out1 <= in68 XOR in72;

  Logical_Operator_out549_out1 <= Logical_Operator_out293_out1 XOR Logical_Operator_out295_out1;

  Logical_Operator_out550_out1 <= Logical_Operator_out294_out1 XOR Logical_Operator_out296_out1;

  Logical_Operator_out551_out1 <= Logical_Operator_out38_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out552_out1 <= in76 XOR in80;

  Logical_Operator_out553_out1 <= Logical_Operator_out297_out1 XOR Logical_Operator_out299_out1;

  Logical_Operator_out554_out1 <= Logical_Operator_out298_out1 XOR Logical_Operator_out300_out1;

  Logical_Operator_out555_out1 <= Logical_Operator_out42_out1 XOR Logical_Operator_out44_out1;

  Logical_Operator_out556_out1 <= in84 XOR in88;

  Logical_Operator_out557_out1 <= Logical_Operator_out301_out1 XOR Logical_Operator_out303_out1;

  Logical_Operator_out558_out1 <= Logical_Operator_out302_out1 XOR Logical_Operator_out304_out1;

  Logical_Operator_out559_out1 <= Logical_Operator_out46_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out560_out1 <= in92 XOR in96;

  Logical_Operator_out561_out1 <= Logical_Operator_out305_out1 XOR Logical_Operator_out307_out1;

  Logical_Operator_out562_out1 <= Logical_Operator_out306_out1 XOR Logical_Operator_out308_out1;

  Logical_Operator_out563_out1 <= Logical_Operator_out50_out1 XOR Logical_Operator_out52_out1;

  Logical_Operator_out564_out1 <= in100 XOR in104;

  Logical_Operator_out565_out1 <= Logical_Operator_out309_out1 XOR Logical_Operator_out311_out1;

  Logical_Operator_out566_out1 <= Logical_Operator_out310_out1 XOR Logical_Operator_out312_out1;

  Logical_Operator_out567_out1 <= Logical_Operator_out54_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out568_out1 <= in108 XOR in112;

  Logical_Operator_out569_out1 <= Logical_Operator_out313_out1 XOR Logical_Operator_out315_out1;

  Logical_Operator_out570_out1 <= Logical_Operator_out314_out1 XOR Logical_Operator_out316_out1;

  Logical_Operator_out571_out1 <= Logical_Operator_out58_out1 XOR Logical_Operator_out60_out1;

  Logical_Operator_out572_out1 <= in116 XOR in120;

  Logical_Operator_out573_out1 <= Logical_Operator_out317_out1 XOR Logical_Operator_out319_out1;

  Logical_Operator_out574_out1 <= Logical_Operator_out318_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out575_out1 <= Logical_Operator_out62_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out576_out1 <= in124 XOR in128;

  Logical_Operator_out577_out1 <= Logical_Operator_out321_out1 XOR Logical_Operator_out323_out1;

  Logical_Operator_out578_out1 <= Logical_Operator_out322_out1 XOR Logical_Operator_out324_out1;

  Logical_Operator_out579_out1 <= Logical_Operator_out66_out1 XOR Logical_Operator_out68_out1;

  Logical_Operator_out580_out1 <= in132 XOR in136;

  Logical_Operator_out581_out1 <= Logical_Operator_out325_out1 XOR Logical_Operator_out327_out1;

  Logical_Operator_out582_out1 <= Logical_Operator_out326_out1 XOR Logical_Operator_out328_out1;

  Logical_Operator_out583_out1 <= Logical_Operator_out70_out1 XOR Logical_Operator_out72_out1;

  Logical_Operator_out584_out1 <= in140 XOR in144;

  Logical_Operator_out585_out1 <= Logical_Operator_out329_out1 XOR Logical_Operator_out331_out1;

  Logical_Operator_out586_out1 <= Logical_Operator_out330_out1 XOR Logical_Operator_out332_out1;

  Logical_Operator_out587_out1 <= Logical_Operator_out74_out1 XOR Logical_Operator_out76_out1;

  Logical_Operator_out588_out1 <= in148 XOR in152;

  Logical_Operator_out589_out1 <= Logical_Operator_out333_out1 XOR Logical_Operator_out335_out1;

  Logical_Operator_out590_out1 <= Logical_Operator_out334_out1 XOR Logical_Operator_out336_out1;

  Logical_Operator_out591_out1 <= Logical_Operator_out78_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out592_out1 <= in156 XOR in160;

  Logical_Operator_out593_out1 <= Logical_Operator_out337_out1 XOR Logical_Operator_out339_out1;

  Logical_Operator_out594_out1 <= Logical_Operator_out338_out1 XOR Logical_Operator_out340_out1;

  Logical_Operator_out595_out1 <= Logical_Operator_out82_out1 XOR Logical_Operator_out84_out1;

  Logical_Operator_out596_out1 <= in164 XOR in168;

  Logical_Operator_out597_out1 <= Logical_Operator_out341_out1 XOR Logical_Operator_out343_out1;

  Logical_Operator_out598_out1 <= Logical_Operator_out342_out1 XOR Logical_Operator_out344_out1;

  Logical_Operator_out599_out1 <= Logical_Operator_out86_out1 XOR Logical_Operator_out88_out1;

  Logical_Operator_out600_out1 <= in172 XOR in176;

  Logical_Operator_out601_out1 <= Logical_Operator_out345_out1 XOR Logical_Operator_out347_out1;

  Logical_Operator_out602_out1 <= Logical_Operator_out346_out1 XOR Logical_Operator_out348_out1;

  Logical_Operator_out603_out1 <= Logical_Operator_out90_out1 XOR Logical_Operator_out92_out1;

  Logical_Operator_out604_out1 <= in180 XOR in184;

  Logical_Operator_out605_out1 <= Logical_Operator_out349_out1 XOR Logical_Operator_out351_out1;

  Logical_Operator_out606_out1 <= Logical_Operator_out350_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out607_out1 <= Logical_Operator_out94_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out608_out1 <= in188 XOR in192;

  Logical_Operator_out609_out1 <= Logical_Operator_out353_out1 XOR Logical_Operator_out355_out1;

  Logical_Operator_out610_out1 <= Logical_Operator_out354_out1 XOR Logical_Operator_out356_out1;

  Logical_Operator_out611_out1 <= Logical_Operator_out98_out1 XOR Logical_Operator_out100_out1;

  Logical_Operator_out612_out1 <= in196 XOR in200;

  Logical_Operator_out613_out1 <= Logical_Operator_out357_out1 XOR Logical_Operator_out359_out1;

  Logical_Operator_out614_out1 <= Logical_Operator_out358_out1 XOR Logical_Operator_out360_out1;

  Logical_Operator_out615_out1 <= Logical_Operator_out102_out1 XOR Logical_Operator_out104_out1;

  Logical_Operator_out616_out1 <= in204 XOR in208;

  Logical_Operator_out617_out1 <= Logical_Operator_out361_out1 XOR Logical_Operator_out363_out1;

  Logical_Operator_out618_out1 <= Logical_Operator_out362_out1 XOR Logical_Operator_out364_out1;

  Logical_Operator_out619_out1 <= Logical_Operator_out106_out1 XOR Logical_Operator_out108_out1;

  Logical_Operator_out620_out1 <= in212 XOR in216;

  Logical_Operator_out621_out1 <= Logical_Operator_out365_out1 XOR Logical_Operator_out367_out1;

  Logical_Operator_out622_out1 <= Logical_Operator_out366_out1 XOR Logical_Operator_out368_out1;

  Logical_Operator_out623_out1 <= Logical_Operator_out110_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out624_out1 <= in220 XOR in224;

  Logical_Operator_out625_out1 <= Logical_Operator_out369_out1 XOR Logical_Operator_out371_out1;

  Logical_Operator_out626_out1 <= Logical_Operator_out370_out1 XOR Logical_Operator_out372_out1;

  Logical_Operator_out627_out1 <= Logical_Operator_out114_out1 XOR Logical_Operator_out116_out1;

  Logical_Operator_out628_out1 <= in228 XOR in232;

  Logical_Operator_out629_out1 <= Logical_Operator_out373_out1 XOR Logical_Operator_out375_out1;

  Logical_Operator_out630_out1 <= Logical_Operator_out374_out1 XOR Logical_Operator_out376_out1;

  Logical_Operator_out631_out1 <= Logical_Operator_out118_out1 XOR Logical_Operator_out120_out1;

  Logical_Operator_out632_out1 <= in236 XOR in240;

  Logical_Operator_out633_out1 <= Logical_Operator_out377_out1 XOR Logical_Operator_out379_out1;

  Logical_Operator_out634_out1 <= Logical_Operator_out378_out1 XOR Logical_Operator_out380_out1;

  Logical_Operator_out635_out1 <= Logical_Operator_out122_out1 XOR Logical_Operator_out124_out1;

  Logical_Operator_out636_out1 <= in244 XOR in248;

  Logical_Operator_out637_out1 <= Logical_Operator_out381_out1 XOR Logical_Operator_out383_out1;

  Logical_Operator_out638_out1 <= Logical_Operator_out382_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out639_out1 <= Logical_Operator_out126_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out640_out1 <= in252 XOR in256;

  Logical_Operator_out641_out1 <= Logical_Operator_out385_out1 XOR Logical_Operator_out387_out1;

  Logical_Operator_out642_out1 <= Logical_Operator_out386_out1 XOR Logical_Operator_out388_out1;

  Logical_Operator_out643_out1 <= Logical_Operator_out130_out1 XOR Logical_Operator_out132_out1;

  Logical_Operator_out644_out1 <= in260 XOR in264;

  Logical_Operator_out645_out1 <= Logical_Operator_out389_out1 XOR Logical_Operator_out391_out1;

  Logical_Operator_out646_out1 <= Logical_Operator_out390_out1 XOR Logical_Operator_out392_out1;

  Logical_Operator_out647_out1 <= Logical_Operator_out134_out1 XOR Logical_Operator_out136_out1;

  Logical_Operator_out648_out1 <= in268 XOR in272;

  Logical_Operator_out649_out1 <= Logical_Operator_out393_out1 XOR Logical_Operator_out395_out1;

  Logical_Operator_out650_out1 <= Logical_Operator_out394_out1 XOR Logical_Operator_out396_out1;

  Logical_Operator_out651_out1 <= Logical_Operator_out138_out1 XOR Logical_Operator_out140_out1;

  Logical_Operator_out652_out1 <= in276 XOR in280;

  Logical_Operator_out653_out1 <= Logical_Operator_out397_out1 XOR Logical_Operator_out399_out1;

  Logical_Operator_out654_out1 <= Logical_Operator_out398_out1 XOR Logical_Operator_out400_out1;

  Logical_Operator_out655_out1 <= Logical_Operator_out142_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out656_out1 <= in284 XOR in288;

  Logical_Operator_out657_out1 <= Logical_Operator_out401_out1 XOR Logical_Operator_out403_out1;

  Logical_Operator_out658_out1 <= Logical_Operator_out402_out1 XOR Logical_Operator_out404_out1;

  Logical_Operator_out659_out1 <= Logical_Operator_out146_out1 XOR Logical_Operator_out148_out1;

  Logical_Operator_out660_out1 <= in292 XOR in296;

  Logical_Operator_out661_out1 <= Logical_Operator_out405_out1 XOR Logical_Operator_out407_out1;

  Logical_Operator_out662_out1 <= Logical_Operator_out406_out1 XOR Logical_Operator_out408_out1;

  Logical_Operator_out663_out1 <= Logical_Operator_out150_out1 XOR Logical_Operator_out152_out1;

  Logical_Operator_out664_out1 <= in300 XOR in304;

  Logical_Operator_out665_out1 <= Logical_Operator_out409_out1 XOR Logical_Operator_out411_out1;

  Logical_Operator_out666_out1 <= Logical_Operator_out410_out1 XOR Logical_Operator_out412_out1;

  Logical_Operator_out667_out1 <= Logical_Operator_out154_out1 XOR Logical_Operator_out156_out1;

  Logical_Operator_out668_out1 <= in308 XOR in312;

  Logical_Operator_out669_out1 <= Logical_Operator_out413_out1 XOR Logical_Operator_out415_out1;

  Logical_Operator_out670_out1 <= Logical_Operator_out414_out1 XOR Logical_Operator_out416_out1;

  Logical_Operator_out671_out1 <= Logical_Operator_out158_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out672_out1 <= in316 XOR in320;

  Logical_Operator_out673_out1 <= Logical_Operator_out417_out1 XOR Logical_Operator_out419_out1;

  Logical_Operator_out674_out1 <= Logical_Operator_out418_out1 XOR Logical_Operator_out420_out1;

  Logical_Operator_out675_out1 <= Logical_Operator_out162_out1 XOR Logical_Operator_out164_out1;

  Logical_Operator_out676_out1 <= in324 XOR in328;

  Logical_Operator_out677_out1 <= Logical_Operator_out421_out1 XOR Logical_Operator_out423_out1;

  Logical_Operator_out678_out1 <= Logical_Operator_out422_out1 XOR Logical_Operator_out424_out1;

  Logical_Operator_out679_out1 <= Logical_Operator_out166_out1 XOR Logical_Operator_out168_out1;

  Logical_Operator_out680_out1 <= in332 XOR in336;

  Logical_Operator_out681_out1 <= Logical_Operator_out425_out1 XOR Logical_Operator_out427_out1;

  Logical_Operator_out682_out1 <= Logical_Operator_out426_out1 XOR Logical_Operator_out428_out1;

  Logical_Operator_out683_out1 <= Logical_Operator_out170_out1 XOR Logical_Operator_out172_out1;

  Logical_Operator_out684_out1 <= in340 XOR in344;

  Logical_Operator_out685_out1 <= Logical_Operator_out429_out1 XOR Logical_Operator_out431_out1;

  Logical_Operator_out686_out1 <= Logical_Operator_out430_out1 XOR Logical_Operator_out432_out1;

  Logical_Operator_out687_out1 <= Logical_Operator_out174_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out688_out1 <= in348 XOR in352;

  Logical_Operator_out689_out1 <= Logical_Operator_out433_out1 XOR Logical_Operator_out435_out1;

  Logical_Operator_out690_out1 <= Logical_Operator_out434_out1 XOR Logical_Operator_out436_out1;

  Logical_Operator_out691_out1 <= Logical_Operator_out178_out1 XOR Logical_Operator_out180_out1;

  Logical_Operator_out692_out1 <= in356 XOR in360;

  Logical_Operator_out693_out1 <= Logical_Operator_out437_out1 XOR Logical_Operator_out439_out1;

  Logical_Operator_out694_out1 <= Logical_Operator_out438_out1 XOR Logical_Operator_out440_out1;

  Logical_Operator_out695_out1 <= Logical_Operator_out182_out1 XOR Logical_Operator_out184_out1;

  Logical_Operator_out696_out1 <= in364 XOR in368;

  Logical_Operator_out697_out1 <= Logical_Operator_out441_out1 XOR Logical_Operator_out443_out1;

  Logical_Operator_out698_out1 <= Logical_Operator_out442_out1 XOR Logical_Operator_out444_out1;

  Logical_Operator_out699_out1 <= Logical_Operator_out186_out1 XOR Logical_Operator_out188_out1;

  Logical_Operator_out700_out1 <= in372 XOR in376;

  Logical_Operator_out701_out1 <= Logical_Operator_out445_out1 XOR Logical_Operator_out447_out1;

  Logical_Operator_out702_out1 <= Logical_Operator_out446_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out703_out1 <= Logical_Operator_out190_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out704_out1 <= in380 XOR in384;

  Logical_Operator_out705_out1 <= Logical_Operator_out449_out1 XOR Logical_Operator_out451_out1;

  Logical_Operator_out706_out1 <= Logical_Operator_out450_out1 XOR Logical_Operator_out452_out1;

  Logical_Operator_out707_out1 <= Logical_Operator_out194_out1 XOR Logical_Operator_out196_out1;

  Logical_Operator_out708_out1 <= in388 XOR in392;

  Logical_Operator_out709_out1 <= Logical_Operator_out453_out1 XOR Logical_Operator_out455_out1;

  Logical_Operator_out710_out1 <= Logical_Operator_out454_out1 XOR Logical_Operator_out456_out1;

  Logical_Operator_out711_out1 <= Logical_Operator_out198_out1 XOR Logical_Operator_out200_out1;

  Logical_Operator_out712_out1 <= in396 XOR in400;

  Logical_Operator_out713_out1 <= Logical_Operator_out457_out1 XOR Logical_Operator_out459_out1;

  Logical_Operator_out714_out1 <= Logical_Operator_out458_out1 XOR Logical_Operator_out460_out1;

  Logical_Operator_out715_out1 <= Logical_Operator_out202_out1 XOR Logical_Operator_out204_out1;

  Logical_Operator_out716_out1 <= in404 XOR in408;

  Logical_Operator_out717_out1 <= Logical_Operator_out461_out1 XOR Logical_Operator_out463_out1;

  Logical_Operator_out718_out1 <= Logical_Operator_out462_out1 XOR Logical_Operator_out464_out1;

  Logical_Operator_out719_out1 <= Logical_Operator_out206_out1 XOR Logical_Operator_out208_out1;

  Logical_Operator_out720_out1 <= in412 XOR in416;

  Logical_Operator_out721_out1 <= Logical_Operator_out465_out1 XOR Logical_Operator_out467_out1;

  Logical_Operator_out722_out1 <= Logical_Operator_out466_out1 XOR Logical_Operator_out468_out1;

  Logical_Operator_out723_out1 <= Logical_Operator_out210_out1 XOR Logical_Operator_out212_out1;

  Logical_Operator_out724_out1 <= in420 XOR in424;

  Logical_Operator_out725_out1 <= Logical_Operator_out469_out1 XOR Logical_Operator_out471_out1;

  Logical_Operator_out726_out1 <= Logical_Operator_out470_out1 XOR Logical_Operator_out472_out1;

  Logical_Operator_out727_out1 <= Logical_Operator_out214_out1 XOR Logical_Operator_out216_out1;

  Logical_Operator_out728_out1 <= in428 XOR in432;

  Logical_Operator_out729_out1 <= Logical_Operator_out473_out1 XOR Logical_Operator_out475_out1;

  Logical_Operator_out730_out1 <= Logical_Operator_out474_out1 XOR Logical_Operator_out476_out1;

  Logical_Operator_out731_out1 <= Logical_Operator_out218_out1 XOR Logical_Operator_out220_out1;

  Logical_Operator_out732_out1 <= in436 XOR in440;

  Logical_Operator_out733_out1 <= Logical_Operator_out477_out1 XOR Logical_Operator_out479_out1;

  Logical_Operator_out734_out1 <= Logical_Operator_out478_out1 XOR Logical_Operator_out480_out1;

  Logical_Operator_out735_out1 <= Logical_Operator_out222_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out736_out1 <= in444 XOR in448;

  Logical_Operator_out737_out1 <= Logical_Operator_out481_out1 XOR Logical_Operator_out483_out1;

  Logical_Operator_out738_out1 <= Logical_Operator_out482_out1 XOR Logical_Operator_out484_out1;

  Logical_Operator_out739_out1 <= Logical_Operator_out226_out1 XOR Logical_Operator_out228_out1;

  Logical_Operator_out740_out1 <= in452 XOR in456;

  Logical_Operator_out741_out1 <= Logical_Operator_out485_out1 XOR Logical_Operator_out487_out1;

  Logical_Operator_out742_out1 <= Logical_Operator_out486_out1 XOR Logical_Operator_out488_out1;

  Logical_Operator_out743_out1 <= Logical_Operator_out230_out1 XOR Logical_Operator_out232_out1;

  Logical_Operator_out744_out1 <= in460 XOR in464;

  Logical_Operator_out745_out1 <= Logical_Operator_out489_out1 XOR Logical_Operator_out491_out1;

  Logical_Operator_out746_out1 <= Logical_Operator_out490_out1 XOR Logical_Operator_out492_out1;

  Logical_Operator_out747_out1 <= Logical_Operator_out234_out1 XOR Logical_Operator_out236_out1;

  Logical_Operator_out748_out1 <= in468 XOR in472;

  Logical_Operator_out749_out1 <= Logical_Operator_out493_out1 XOR Logical_Operator_out495_out1;

  Logical_Operator_out750_out1 <= Logical_Operator_out494_out1 XOR Logical_Operator_out496_out1;

  Logical_Operator_out751_out1 <= Logical_Operator_out238_out1 XOR Logical_Operator_out240_out1;

  Logical_Operator_out752_out1 <= in476 XOR in480;

  Logical_Operator_out753_out1 <= Logical_Operator_out497_out1 XOR Logical_Operator_out499_out1;

  Logical_Operator_out754_out1 <= Logical_Operator_out498_out1 XOR Logical_Operator_out500_out1;

  Logical_Operator_out755_out1 <= Logical_Operator_out242_out1 XOR Logical_Operator_out244_out1;

  Logical_Operator_out756_out1 <= in484 XOR in488;

  Logical_Operator_out757_out1 <= Logical_Operator_out501_out1 XOR Logical_Operator_out503_out1;

  Logical_Operator_out758_out1 <= Logical_Operator_out502_out1 XOR Logical_Operator_out504_out1;

  Logical_Operator_out759_out1 <= Logical_Operator_out246_out1 XOR Logical_Operator_out248_out1;

  Logical_Operator_out760_out1 <= in492 XOR in496;

  Logical_Operator_out761_out1 <= Logical_Operator_out505_out1 XOR Logical_Operator_out507_out1;

  Logical_Operator_out762_out1 <= Logical_Operator_out506_out1 XOR Logical_Operator_out508_out1;

  Logical_Operator_out763_out1 <= Logical_Operator_out250_out1 XOR Logical_Operator_out252_out1;

  Logical_Operator_out764_out1 <= in500 XOR in504;

  Logical_Operator_out765_out1 <= Logical_Operator_out509_out1 XOR Logical_Operator_out511_out1;

  Logical_Operator_out766_out1 <= Logical_Operator_out510_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out767_out1 <= Logical_Operator_out254_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out768_out1 <= in508 XOR in512;

  Logical_Operator_out769_out1 <= Logical_Operator_out513_out1 XOR Logical_Operator_out517_out1;

  Logical_Operator_out770_out1 <= Logical_Operator_out514_out1 XOR Logical_Operator_out518_out1;

  Logical_Operator_out771_out1 <= Logical_Operator_out515_out1 XOR Logical_Operator_out519_out1;

  Logical_Operator_out772_out1 <= Logical_Operator_out516_out1 XOR Logical_Operator_out520_out1;

  Logical_Operator_out773_out1 <= Logical_Operator_out259_out1 XOR Logical_Operator_out263_out1;

  Logical_Operator_out774_out1 <= Logical_Operator_out260_out1 XOR Logical_Operator_out264_out1;

  Logical_Operator_out775_out1 <= Logical_Operator_out4_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out776_out1 <= in8 XOR in16;

  Logical_Operator_out777_out1 <= Logical_Operator_out521_out1 XOR Logical_Operator_out525_out1;

  Logical_Operator_out778_out1 <= Logical_Operator_out522_out1 XOR Logical_Operator_out526_out1;

  Logical_Operator_out779_out1 <= Logical_Operator_out523_out1 XOR Logical_Operator_out527_out1;

  Logical_Operator_out780_out1 <= Logical_Operator_out524_out1 XOR Logical_Operator_out528_out1;

  Logical_Operator_out781_out1 <= Logical_Operator_out267_out1 XOR Logical_Operator_out271_out1;

  Logical_Operator_out782_out1 <= Logical_Operator_out268_out1 XOR Logical_Operator_out272_out1;

  Logical_Operator_out783_out1 <= Logical_Operator_out12_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out784_out1 <= in24 XOR in32;

  Logical_Operator_out785_out1 <= Logical_Operator_out529_out1 XOR Logical_Operator_out533_out1;

  Logical_Operator_out786_out1 <= Logical_Operator_out530_out1 XOR Logical_Operator_out534_out1;

  Logical_Operator_out787_out1 <= Logical_Operator_out531_out1 XOR Logical_Operator_out535_out1;

  Logical_Operator_out788_out1 <= Logical_Operator_out532_out1 XOR Logical_Operator_out536_out1;

  Logical_Operator_out789_out1 <= Logical_Operator_out275_out1 XOR Logical_Operator_out279_out1;

  Logical_Operator_out790_out1 <= Logical_Operator_out276_out1 XOR Logical_Operator_out280_out1;

  Logical_Operator_out791_out1 <= Logical_Operator_out20_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out792_out1 <= in40 XOR in48;

  Logical_Operator_out793_out1 <= Logical_Operator_out537_out1 XOR Logical_Operator_out541_out1;

  Logical_Operator_out794_out1 <= Logical_Operator_out538_out1 XOR Logical_Operator_out542_out1;

  Logical_Operator_out795_out1 <= Logical_Operator_out539_out1 XOR Logical_Operator_out543_out1;

  Logical_Operator_out796_out1 <= Logical_Operator_out540_out1 XOR Logical_Operator_out544_out1;

  Logical_Operator_out797_out1 <= Logical_Operator_out283_out1 XOR Logical_Operator_out287_out1;

  Logical_Operator_out798_out1 <= Logical_Operator_out284_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out799_out1 <= Logical_Operator_out28_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out800_out1 <= in56 XOR in64;

  Logical_Operator_out801_out1 <= Logical_Operator_out545_out1 XOR Logical_Operator_out549_out1;

  Logical_Operator_out802_out1 <= Logical_Operator_out546_out1 XOR Logical_Operator_out550_out1;

  Logical_Operator_out803_out1 <= Logical_Operator_out547_out1 XOR Logical_Operator_out551_out1;

  Logical_Operator_out804_out1 <= Logical_Operator_out548_out1 XOR Logical_Operator_out552_out1;

  Logical_Operator_out805_out1 <= Logical_Operator_out291_out1 XOR Logical_Operator_out295_out1;

  Logical_Operator_out806_out1 <= Logical_Operator_out292_out1 XOR Logical_Operator_out296_out1;

  Logical_Operator_out807_out1 <= Logical_Operator_out36_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out808_out1 <= in72 XOR in80;

  Logical_Operator_out809_out1 <= Logical_Operator_out553_out1 XOR Logical_Operator_out557_out1;

  Logical_Operator_out810_out1 <= Logical_Operator_out554_out1 XOR Logical_Operator_out558_out1;

  Logical_Operator_out811_out1 <= Logical_Operator_out555_out1 XOR Logical_Operator_out559_out1;

  Logical_Operator_out812_out1 <= Logical_Operator_out556_out1 XOR Logical_Operator_out560_out1;

  Logical_Operator_out813_out1 <= Logical_Operator_out299_out1 XOR Logical_Operator_out303_out1;

  Logical_Operator_out814_out1 <= Logical_Operator_out300_out1 XOR Logical_Operator_out304_out1;

  Logical_Operator_out815_out1 <= Logical_Operator_out44_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out816_out1 <= in88 XOR in96;

  Logical_Operator_out817_out1 <= Logical_Operator_out561_out1 XOR Logical_Operator_out565_out1;

  Logical_Operator_out818_out1 <= Logical_Operator_out562_out1 XOR Logical_Operator_out566_out1;

  Logical_Operator_out819_out1 <= Logical_Operator_out563_out1 XOR Logical_Operator_out567_out1;

  Logical_Operator_out820_out1 <= Logical_Operator_out564_out1 XOR Logical_Operator_out568_out1;

  Logical_Operator_out821_out1 <= Logical_Operator_out307_out1 XOR Logical_Operator_out311_out1;

  Logical_Operator_out822_out1 <= Logical_Operator_out308_out1 XOR Logical_Operator_out312_out1;

  Logical_Operator_out823_out1 <= Logical_Operator_out52_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out824_out1 <= in104 XOR in112;

  Logical_Operator_out825_out1 <= Logical_Operator_out569_out1 XOR Logical_Operator_out573_out1;

  Logical_Operator_out826_out1 <= Logical_Operator_out570_out1 XOR Logical_Operator_out574_out1;

  Logical_Operator_out827_out1 <= Logical_Operator_out571_out1 XOR Logical_Operator_out575_out1;

  Logical_Operator_out828_out1 <= Logical_Operator_out572_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out829_out1 <= Logical_Operator_out315_out1 XOR Logical_Operator_out319_out1;

  Logical_Operator_out830_out1 <= Logical_Operator_out316_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out831_out1 <= Logical_Operator_out60_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out832_out1 <= in120 XOR in128;

  Logical_Operator_out833_out1 <= Logical_Operator_out577_out1 XOR Logical_Operator_out581_out1;

  Logical_Operator_out834_out1 <= Logical_Operator_out578_out1 XOR Logical_Operator_out582_out1;

  Logical_Operator_out835_out1 <= Logical_Operator_out579_out1 XOR Logical_Operator_out583_out1;

  Logical_Operator_out836_out1 <= Logical_Operator_out580_out1 XOR Logical_Operator_out584_out1;

  Logical_Operator_out837_out1 <= Logical_Operator_out323_out1 XOR Logical_Operator_out327_out1;

  Logical_Operator_out838_out1 <= Logical_Operator_out324_out1 XOR Logical_Operator_out328_out1;

  Logical_Operator_out839_out1 <= Logical_Operator_out68_out1 XOR Logical_Operator_out72_out1;

  Logical_Operator_out840_out1 <= in136 XOR in144;

  Logical_Operator_out841_out1 <= Logical_Operator_out585_out1 XOR Logical_Operator_out589_out1;

  Logical_Operator_out842_out1 <= Logical_Operator_out586_out1 XOR Logical_Operator_out590_out1;

  Logical_Operator_out843_out1 <= Logical_Operator_out587_out1 XOR Logical_Operator_out591_out1;

  Logical_Operator_out844_out1 <= Logical_Operator_out588_out1 XOR Logical_Operator_out592_out1;

  Logical_Operator_out845_out1 <= Logical_Operator_out331_out1 XOR Logical_Operator_out335_out1;

  Logical_Operator_out846_out1 <= Logical_Operator_out332_out1 XOR Logical_Operator_out336_out1;

  Logical_Operator_out847_out1 <= Logical_Operator_out76_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out848_out1 <= in152 XOR in160;

  Logical_Operator_out849_out1 <= Logical_Operator_out593_out1 XOR Logical_Operator_out597_out1;

  Logical_Operator_out850_out1 <= Logical_Operator_out594_out1 XOR Logical_Operator_out598_out1;

  Logical_Operator_out851_out1 <= Logical_Operator_out595_out1 XOR Logical_Operator_out599_out1;

  Logical_Operator_out852_out1 <= Logical_Operator_out596_out1 XOR Logical_Operator_out600_out1;

  Logical_Operator_out853_out1 <= Logical_Operator_out339_out1 XOR Logical_Operator_out343_out1;

  Logical_Operator_out854_out1 <= Logical_Operator_out340_out1 XOR Logical_Operator_out344_out1;

  Logical_Operator_out855_out1 <= Logical_Operator_out84_out1 XOR Logical_Operator_out88_out1;

  Logical_Operator_out856_out1 <= in168 XOR in176;

  Logical_Operator_out857_out1 <= Logical_Operator_out601_out1 XOR Logical_Operator_out605_out1;

  Logical_Operator_out858_out1 <= Logical_Operator_out602_out1 XOR Logical_Operator_out606_out1;

  Logical_Operator_out859_out1 <= Logical_Operator_out603_out1 XOR Logical_Operator_out607_out1;

  Logical_Operator_out860_out1 <= Logical_Operator_out604_out1 XOR Logical_Operator_out608_out1;

  Logical_Operator_out861_out1 <= Logical_Operator_out347_out1 XOR Logical_Operator_out351_out1;

  Logical_Operator_out862_out1 <= Logical_Operator_out348_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out863_out1 <= Logical_Operator_out92_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out864_out1 <= in184 XOR in192;

  Logical_Operator_out865_out1 <= Logical_Operator_out609_out1 XOR Logical_Operator_out613_out1;

  Logical_Operator_out866_out1 <= Logical_Operator_out610_out1 XOR Logical_Operator_out614_out1;

  Logical_Operator_out867_out1 <= Logical_Operator_out611_out1 XOR Logical_Operator_out615_out1;

  Logical_Operator_out868_out1 <= Logical_Operator_out612_out1 XOR Logical_Operator_out616_out1;

  Logical_Operator_out869_out1 <= Logical_Operator_out355_out1 XOR Logical_Operator_out359_out1;

  Logical_Operator_out870_out1 <= Logical_Operator_out356_out1 XOR Logical_Operator_out360_out1;

  Logical_Operator_out871_out1 <= Logical_Operator_out100_out1 XOR Logical_Operator_out104_out1;

  Logical_Operator_out872_out1 <= in200 XOR in208;

  Logical_Operator_out873_out1 <= Logical_Operator_out617_out1 XOR Logical_Operator_out621_out1;

  Logical_Operator_out874_out1 <= Logical_Operator_out618_out1 XOR Logical_Operator_out622_out1;

  Logical_Operator_out875_out1 <= Logical_Operator_out619_out1 XOR Logical_Operator_out623_out1;

  Logical_Operator_out876_out1 <= Logical_Operator_out620_out1 XOR Logical_Operator_out624_out1;

  Logical_Operator_out877_out1 <= Logical_Operator_out363_out1 XOR Logical_Operator_out367_out1;

  Logical_Operator_out878_out1 <= Logical_Operator_out364_out1 XOR Logical_Operator_out368_out1;

  Logical_Operator_out879_out1 <= Logical_Operator_out108_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out880_out1 <= in216 XOR in224;

  Logical_Operator_out881_out1 <= Logical_Operator_out625_out1 XOR Logical_Operator_out629_out1;

  Logical_Operator_out882_out1 <= Logical_Operator_out626_out1 XOR Logical_Operator_out630_out1;

  Logical_Operator_out883_out1 <= Logical_Operator_out627_out1 XOR Logical_Operator_out631_out1;

  Logical_Operator_out884_out1 <= Logical_Operator_out628_out1 XOR Logical_Operator_out632_out1;

  Logical_Operator_out885_out1 <= Logical_Operator_out371_out1 XOR Logical_Operator_out375_out1;

  Logical_Operator_out886_out1 <= Logical_Operator_out372_out1 XOR Logical_Operator_out376_out1;

  Logical_Operator_out887_out1 <= Logical_Operator_out116_out1 XOR Logical_Operator_out120_out1;

  Logical_Operator_out888_out1 <= in232 XOR in240;

  Logical_Operator_out889_out1 <= Logical_Operator_out633_out1 XOR Logical_Operator_out637_out1;

  Logical_Operator_out890_out1 <= Logical_Operator_out634_out1 XOR Logical_Operator_out638_out1;

  Logical_Operator_out891_out1 <= Logical_Operator_out635_out1 XOR Logical_Operator_out639_out1;

  Logical_Operator_out892_out1 <= Logical_Operator_out636_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out893_out1 <= Logical_Operator_out379_out1 XOR Logical_Operator_out383_out1;

  Logical_Operator_out894_out1 <= Logical_Operator_out380_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out895_out1 <= Logical_Operator_out124_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out896_out1 <= in248 XOR in256;

  Logical_Operator_out897_out1 <= Logical_Operator_out641_out1 XOR Logical_Operator_out645_out1;

  Logical_Operator_out898_out1 <= Logical_Operator_out642_out1 XOR Logical_Operator_out646_out1;

  Logical_Operator_out899_out1 <= Logical_Operator_out643_out1 XOR Logical_Operator_out647_out1;

  Logical_Operator_out900_out1 <= Logical_Operator_out644_out1 XOR Logical_Operator_out648_out1;

  Logical_Operator_out901_out1 <= Logical_Operator_out387_out1 XOR Logical_Operator_out391_out1;

  Logical_Operator_out902_out1 <= Logical_Operator_out388_out1 XOR Logical_Operator_out392_out1;

  Logical_Operator_out903_out1 <= Logical_Operator_out132_out1 XOR Logical_Operator_out136_out1;

  Logical_Operator_out904_out1 <= in264 XOR in272;

  Logical_Operator_out905_out1 <= Logical_Operator_out649_out1 XOR Logical_Operator_out653_out1;

  Logical_Operator_out906_out1 <= Logical_Operator_out650_out1 XOR Logical_Operator_out654_out1;

  Logical_Operator_out907_out1 <= Logical_Operator_out651_out1 XOR Logical_Operator_out655_out1;

  Logical_Operator_out908_out1 <= Logical_Operator_out652_out1 XOR Logical_Operator_out656_out1;

  Logical_Operator_out909_out1 <= Logical_Operator_out395_out1 XOR Logical_Operator_out399_out1;

  Logical_Operator_out910_out1 <= Logical_Operator_out396_out1 XOR Logical_Operator_out400_out1;

  Logical_Operator_out911_out1 <= Logical_Operator_out140_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out912_out1 <= in280 XOR in288;

  Logical_Operator_out913_out1 <= Logical_Operator_out657_out1 XOR Logical_Operator_out661_out1;

  Logical_Operator_out914_out1 <= Logical_Operator_out658_out1 XOR Logical_Operator_out662_out1;

  Logical_Operator_out915_out1 <= Logical_Operator_out659_out1 XOR Logical_Operator_out663_out1;

  Logical_Operator_out916_out1 <= Logical_Operator_out660_out1 XOR Logical_Operator_out664_out1;

  Logical_Operator_out917_out1 <= Logical_Operator_out403_out1 XOR Logical_Operator_out407_out1;

  Logical_Operator_out918_out1 <= Logical_Operator_out404_out1 XOR Logical_Operator_out408_out1;

  Logical_Operator_out919_out1 <= Logical_Operator_out148_out1 XOR Logical_Operator_out152_out1;

  Logical_Operator_out920_out1 <= in296 XOR in304;

  Logical_Operator_out921_out1 <= Logical_Operator_out665_out1 XOR Logical_Operator_out669_out1;

  Logical_Operator_out922_out1 <= Logical_Operator_out666_out1 XOR Logical_Operator_out670_out1;

  Logical_Operator_out923_out1 <= Logical_Operator_out667_out1 XOR Logical_Operator_out671_out1;

  Logical_Operator_out924_out1 <= Logical_Operator_out668_out1 XOR Logical_Operator_out672_out1;

  Logical_Operator_out925_out1 <= Logical_Operator_out411_out1 XOR Logical_Operator_out415_out1;

  Logical_Operator_out926_out1 <= Logical_Operator_out412_out1 XOR Logical_Operator_out416_out1;

  Logical_Operator_out927_out1 <= Logical_Operator_out156_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out928_out1 <= in312 XOR in320;

  Logical_Operator_out929_out1 <= Logical_Operator_out673_out1 XOR Logical_Operator_out677_out1;

  Logical_Operator_out930_out1 <= Logical_Operator_out674_out1 XOR Logical_Operator_out678_out1;

  Logical_Operator_out931_out1 <= Logical_Operator_out675_out1 XOR Logical_Operator_out679_out1;

  Logical_Operator_out932_out1 <= Logical_Operator_out676_out1 XOR Logical_Operator_out680_out1;

  Logical_Operator_out933_out1 <= Logical_Operator_out419_out1 XOR Logical_Operator_out423_out1;

  Logical_Operator_out934_out1 <= Logical_Operator_out420_out1 XOR Logical_Operator_out424_out1;

  Logical_Operator_out935_out1 <= Logical_Operator_out164_out1 XOR Logical_Operator_out168_out1;

  Logical_Operator_out936_out1 <= in328 XOR in336;

  Logical_Operator_out937_out1 <= Logical_Operator_out681_out1 XOR Logical_Operator_out685_out1;

  Logical_Operator_out938_out1 <= Logical_Operator_out682_out1 XOR Logical_Operator_out686_out1;

  Logical_Operator_out939_out1 <= Logical_Operator_out683_out1 XOR Logical_Operator_out687_out1;

  Logical_Operator_out940_out1 <= Logical_Operator_out684_out1 XOR Logical_Operator_out688_out1;

  Logical_Operator_out941_out1 <= Logical_Operator_out427_out1 XOR Logical_Operator_out431_out1;

  Logical_Operator_out942_out1 <= Logical_Operator_out428_out1 XOR Logical_Operator_out432_out1;

  Logical_Operator_out943_out1 <= Logical_Operator_out172_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out944_out1 <= in344 XOR in352;

  Logical_Operator_out945_out1 <= Logical_Operator_out689_out1 XOR Logical_Operator_out693_out1;

  Logical_Operator_out946_out1 <= Logical_Operator_out690_out1 XOR Logical_Operator_out694_out1;

  Logical_Operator_out947_out1 <= Logical_Operator_out691_out1 XOR Logical_Operator_out695_out1;

  Logical_Operator_out948_out1 <= Logical_Operator_out692_out1 XOR Logical_Operator_out696_out1;

  Logical_Operator_out949_out1 <= Logical_Operator_out435_out1 XOR Logical_Operator_out439_out1;

  Logical_Operator_out950_out1 <= Logical_Operator_out436_out1 XOR Logical_Operator_out440_out1;

  Logical_Operator_out951_out1 <= Logical_Operator_out180_out1 XOR Logical_Operator_out184_out1;

  Logical_Operator_out952_out1 <= in360 XOR in368;

  Logical_Operator_out953_out1 <= Logical_Operator_out697_out1 XOR Logical_Operator_out701_out1;

  Logical_Operator_out954_out1 <= Logical_Operator_out698_out1 XOR Logical_Operator_out702_out1;

  Logical_Operator_out955_out1 <= Logical_Operator_out699_out1 XOR Logical_Operator_out703_out1;

  Logical_Operator_out956_out1 <= Logical_Operator_out700_out1 XOR Logical_Operator_out704_out1;

  Logical_Operator_out957_out1 <= Logical_Operator_out443_out1 XOR Logical_Operator_out447_out1;

  Logical_Operator_out958_out1 <= Logical_Operator_out444_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out959_out1 <= Logical_Operator_out188_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out960_out1 <= in376 XOR in384;

  Logical_Operator_out961_out1 <= Logical_Operator_out705_out1 XOR Logical_Operator_out709_out1;

  Logical_Operator_out962_out1 <= Logical_Operator_out706_out1 XOR Logical_Operator_out710_out1;

  Logical_Operator_out963_out1 <= Logical_Operator_out707_out1 XOR Logical_Operator_out711_out1;

  Logical_Operator_out964_out1 <= Logical_Operator_out708_out1 XOR Logical_Operator_out712_out1;

  Logical_Operator_out965_out1 <= Logical_Operator_out451_out1 XOR Logical_Operator_out455_out1;

  Logical_Operator_out966_out1 <= Logical_Operator_out452_out1 XOR Logical_Operator_out456_out1;

  Logical_Operator_out967_out1 <= Logical_Operator_out196_out1 XOR Logical_Operator_out200_out1;

  Logical_Operator_out968_out1 <= in392 XOR in400;

  Logical_Operator_out969_out1 <= Logical_Operator_out713_out1 XOR Logical_Operator_out717_out1;

  Logical_Operator_out970_out1 <= Logical_Operator_out714_out1 XOR Logical_Operator_out718_out1;

  Logical_Operator_out971_out1 <= Logical_Operator_out715_out1 XOR Logical_Operator_out719_out1;

  Logical_Operator_out972_out1 <= Logical_Operator_out716_out1 XOR Logical_Operator_out720_out1;

  Logical_Operator_out973_out1 <= Logical_Operator_out459_out1 XOR Logical_Operator_out463_out1;

  Logical_Operator_out974_out1 <= Logical_Operator_out460_out1 XOR Logical_Operator_out464_out1;

  Logical_Operator_out975_out1 <= Logical_Operator_out204_out1 XOR Logical_Operator_out208_out1;

  Logical_Operator_out976_out1 <= in408 XOR in416;

  Logical_Operator_out977_out1 <= Logical_Operator_out721_out1 XOR Logical_Operator_out725_out1;

  Logical_Operator_out978_out1 <= Logical_Operator_out722_out1 XOR Logical_Operator_out726_out1;

  Logical_Operator_out979_out1 <= Logical_Operator_out723_out1 XOR Logical_Operator_out727_out1;

  Logical_Operator_out980_out1 <= Logical_Operator_out724_out1 XOR Logical_Operator_out728_out1;

  Logical_Operator_out981_out1 <= Logical_Operator_out467_out1 XOR Logical_Operator_out471_out1;

  Logical_Operator_out982_out1 <= Logical_Operator_out468_out1 XOR Logical_Operator_out472_out1;

  Logical_Operator_out983_out1 <= Logical_Operator_out212_out1 XOR Logical_Operator_out216_out1;

  Logical_Operator_out984_out1 <= in424 XOR in432;

  Logical_Operator_out985_out1 <= Logical_Operator_out729_out1 XOR Logical_Operator_out733_out1;

  Logical_Operator_out986_out1 <= Logical_Operator_out730_out1 XOR Logical_Operator_out734_out1;

  Logical_Operator_out987_out1 <= Logical_Operator_out731_out1 XOR Logical_Operator_out735_out1;

  Logical_Operator_out988_out1 <= Logical_Operator_out732_out1 XOR Logical_Operator_out736_out1;

  Logical_Operator_out989_out1 <= Logical_Operator_out475_out1 XOR Logical_Operator_out479_out1;

  Logical_Operator_out990_out1 <= Logical_Operator_out476_out1 XOR Logical_Operator_out480_out1;

  Logical_Operator_out991_out1 <= Logical_Operator_out220_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out992_out1 <= in440 XOR in448;

  Logical_Operator_out993_out1 <= Logical_Operator_out737_out1 XOR Logical_Operator_out741_out1;

  Logical_Operator_out994_out1 <= Logical_Operator_out738_out1 XOR Logical_Operator_out742_out1;

  Logical_Operator_out995_out1 <= Logical_Operator_out739_out1 XOR Logical_Operator_out743_out1;

  Logical_Operator_out996_out1 <= Logical_Operator_out740_out1 XOR Logical_Operator_out744_out1;

  Logical_Operator_out997_out1 <= Logical_Operator_out483_out1 XOR Logical_Operator_out487_out1;

  Logical_Operator_out998_out1 <= Logical_Operator_out484_out1 XOR Logical_Operator_out488_out1;

  Logical_Operator_out999_out1 <= Logical_Operator_out228_out1 XOR Logical_Operator_out232_out1;

  Logical_Operator_out1000_out1 <= in456 XOR in464;

  Logical_Operator_out1001_out1 <= Logical_Operator_out745_out1 XOR Logical_Operator_out749_out1;

  Logical_Operator_out1002_out1 <= Logical_Operator_out746_out1 XOR Logical_Operator_out750_out1;

  Logical_Operator_out1003_out1 <= Logical_Operator_out747_out1 XOR Logical_Operator_out751_out1;

  Logical_Operator_out1004_out1 <= Logical_Operator_out748_out1 XOR Logical_Operator_out752_out1;

  Logical_Operator_out1005_out1 <= Logical_Operator_out491_out1 XOR Logical_Operator_out495_out1;

  Logical_Operator_out1006_out1 <= Logical_Operator_out492_out1 XOR Logical_Operator_out496_out1;

  Logical_Operator_out1007_out1 <= Logical_Operator_out236_out1 XOR Logical_Operator_out240_out1;

  Logical_Operator_out1008_out1 <= in472 XOR in480;

  Logical_Operator_out1009_out1 <= Logical_Operator_out753_out1 XOR Logical_Operator_out757_out1;

  Logical_Operator_out1010_out1 <= Logical_Operator_out754_out1 XOR Logical_Operator_out758_out1;

  Logical_Operator_out1011_out1 <= Logical_Operator_out755_out1 XOR Logical_Operator_out759_out1;

  Logical_Operator_out1012_out1 <= Logical_Operator_out756_out1 XOR Logical_Operator_out760_out1;

  Logical_Operator_out1013_out1 <= Logical_Operator_out499_out1 XOR Logical_Operator_out503_out1;

  Logical_Operator_out1014_out1 <= Logical_Operator_out500_out1 XOR Logical_Operator_out504_out1;

  Logical_Operator_out1015_out1 <= Logical_Operator_out244_out1 XOR Logical_Operator_out248_out1;

  Logical_Operator_out1016_out1 <= in488 XOR in496;

  Logical_Operator_out1017_out1 <= Logical_Operator_out761_out1 XOR Logical_Operator_out765_out1;

  Logical_Operator_out1018_out1 <= Logical_Operator_out762_out1 XOR Logical_Operator_out766_out1;

  Logical_Operator_out1019_out1 <= Logical_Operator_out763_out1 XOR Logical_Operator_out767_out1;

  Logical_Operator_out1020_out1 <= Logical_Operator_out764_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out1021_out1 <= Logical_Operator_out507_out1 XOR Logical_Operator_out511_out1;

  Logical_Operator_out1022_out1 <= Logical_Operator_out508_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out1023_out1 <= Logical_Operator_out252_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out1024_out1 <= in504 XOR in512;

  Logical_Operator_out1025_out1 <= Logical_Operator_out769_out1 XOR Logical_Operator_out777_out1;

  Logical_Operator_out1026_out1 <= Logical_Operator_out770_out1 XOR Logical_Operator_out778_out1;

  Logical_Operator_out1027_out1 <= Logical_Operator_out771_out1 XOR Logical_Operator_out779_out1;

  Logical_Operator_out1028_out1 <= Logical_Operator_out772_out1 XOR Logical_Operator_out780_out1;

  Logical_Operator_out1029_out1 <= Logical_Operator_out773_out1 XOR Logical_Operator_out781_out1;

  Logical_Operator_out1030_out1 <= Logical_Operator_out774_out1 XOR Logical_Operator_out782_out1;

  Logical_Operator_out1031_out1 <= Logical_Operator_out775_out1 XOR Logical_Operator_out783_out1;

  Logical_Operator_out1032_out1 <= Logical_Operator_out776_out1 XOR Logical_Operator_out784_out1;

  Logical_Operator_out1033_out1 <= Logical_Operator_out517_out1 XOR Logical_Operator_out525_out1;

  Logical_Operator_out1034_out1 <= Logical_Operator_out518_out1 XOR Logical_Operator_out526_out1;

  Logical_Operator_out1035_out1 <= Logical_Operator_out519_out1 XOR Logical_Operator_out527_out1;

  Logical_Operator_out1036_out1 <= Logical_Operator_out520_out1 XOR Logical_Operator_out528_out1;

  Logical_Operator_out1037_out1 <= Logical_Operator_out263_out1 XOR Logical_Operator_out271_out1;

  Logical_Operator_out1038_out1 <= Logical_Operator_out264_out1 XOR Logical_Operator_out272_out1;

  Logical_Operator_out1039_out1 <= Logical_Operator_out8_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out1040_out1 <= in16 XOR in32;

  Logical_Operator_out1041_out1 <= Logical_Operator_out785_out1 XOR Logical_Operator_out793_out1;

  Logical_Operator_out1042_out1 <= Logical_Operator_out786_out1 XOR Logical_Operator_out794_out1;

  Logical_Operator_out1043_out1 <= Logical_Operator_out787_out1 XOR Logical_Operator_out795_out1;

  Logical_Operator_out1044_out1 <= Logical_Operator_out788_out1 XOR Logical_Operator_out796_out1;

  Logical_Operator_out1045_out1 <= Logical_Operator_out789_out1 XOR Logical_Operator_out797_out1;

  Logical_Operator_out1046_out1 <= Logical_Operator_out790_out1 XOR Logical_Operator_out798_out1;

  Logical_Operator_out1047_out1 <= Logical_Operator_out791_out1 XOR Logical_Operator_out799_out1;

  Logical_Operator_out1048_out1 <= Logical_Operator_out792_out1 XOR Logical_Operator_out800_out1;

  Logical_Operator_out1049_out1 <= Logical_Operator_out533_out1 XOR Logical_Operator_out541_out1;

  Logical_Operator_out1050_out1 <= Logical_Operator_out534_out1 XOR Logical_Operator_out542_out1;

  Logical_Operator_out1051_out1 <= Logical_Operator_out535_out1 XOR Logical_Operator_out543_out1;

  Logical_Operator_out1052_out1 <= Logical_Operator_out536_out1 XOR Logical_Operator_out544_out1;

  Logical_Operator_out1053_out1 <= Logical_Operator_out279_out1 XOR Logical_Operator_out287_out1;

  Logical_Operator_out1054_out1 <= Logical_Operator_out280_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out1055_out1 <= Logical_Operator_out24_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out1056_out1 <= in48 XOR in64;

  Logical_Operator_out1057_out1 <= Logical_Operator_out801_out1 XOR Logical_Operator_out809_out1;

  Logical_Operator_out1058_out1 <= Logical_Operator_out802_out1 XOR Logical_Operator_out810_out1;

  Logical_Operator_out1059_out1 <= Logical_Operator_out803_out1 XOR Logical_Operator_out811_out1;

  Logical_Operator_out1060_out1 <= Logical_Operator_out804_out1 XOR Logical_Operator_out812_out1;

  Logical_Operator_out1061_out1 <= Logical_Operator_out805_out1 XOR Logical_Operator_out813_out1;

  Logical_Operator_out1062_out1 <= Logical_Operator_out806_out1 XOR Logical_Operator_out814_out1;

  Logical_Operator_out1063_out1 <= Logical_Operator_out807_out1 XOR Logical_Operator_out815_out1;

  Logical_Operator_out1064_out1 <= Logical_Operator_out808_out1 XOR Logical_Operator_out816_out1;

  Logical_Operator_out1065_out1 <= Logical_Operator_out549_out1 XOR Logical_Operator_out557_out1;

  Logical_Operator_out1066_out1 <= Logical_Operator_out550_out1 XOR Logical_Operator_out558_out1;

  Logical_Operator_out1067_out1 <= Logical_Operator_out551_out1 XOR Logical_Operator_out559_out1;

  Logical_Operator_out1068_out1 <= Logical_Operator_out552_out1 XOR Logical_Operator_out560_out1;

  Logical_Operator_out1069_out1 <= Logical_Operator_out295_out1 XOR Logical_Operator_out303_out1;

  Logical_Operator_out1070_out1 <= Logical_Operator_out296_out1 XOR Logical_Operator_out304_out1;

  Logical_Operator_out1071_out1 <= Logical_Operator_out40_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out1072_out1 <= in80 XOR in96;

  Logical_Operator_out1073_out1 <= Logical_Operator_out817_out1 XOR Logical_Operator_out825_out1;

  Logical_Operator_out1074_out1 <= Logical_Operator_out818_out1 XOR Logical_Operator_out826_out1;

  Logical_Operator_out1075_out1 <= Logical_Operator_out819_out1 XOR Logical_Operator_out827_out1;

  Logical_Operator_out1076_out1 <= Logical_Operator_out820_out1 XOR Logical_Operator_out828_out1;

  Logical_Operator_out1077_out1 <= Logical_Operator_out821_out1 XOR Logical_Operator_out829_out1;

  Logical_Operator_out1078_out1 <= Logical_Operator_out822_out1 XOR Logical_Operator_out830_out1;

  Logical_Operator_out1079_out1 <= Logical_Operator_out823_out1 XOR Logical_Operator_out831_out1;

  Logical_Operator_out1080_out1 <= Logical_Operator_out824_out1 XOR Logical_Operator_out832_out1;

  Logical_Operator_out1081_out1 <= Logical_Operator_out565_out1 XOR Logical_Operator_out573_out1;

  Logical_Operator_out1082_out1 <= Logical_Operator_out566_out1 XOR Logical_Operator_out574_out1;

  Logical_Operator_out1083_out1 <= Logical_Operator_out567_out1 XOR Logical_Operator_out575_out1;

  Logical_Operator_out1084_out1 <= Logical_Operator_out568_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out1085_out1 <= Logical_Operator_out311_out1 XOR Logical_Operator_out319_out1;

  Logical_Operator_out1086_out1 <= Logical_Operator_out312_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out1087_out1 <= Logical_Operator_out56_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out1088_out1 <= in112 XOR in128;

  Logical_Operator_out1089_out1 <= Logical_Operator_out833_out1 XOR Logical_Operator_out841_out1;

  Logical_Operator_out1090_out1 <= Logical_Operator_out834_out1 XOR Logical_Operator_out842_out1;

  Logical_Operator_out1091_out1 <= Logical_Operator_out835_out1 XOR Logical_Operator_out843_out1;

  Logical_Operator_out1092_out1 <= Logical_Operator_out836_out1 XOR Logical_Operator_out844_out1;

  Logical_Operator_out1093_out1 <= Logical_Operator_out837_out1 XOR Logical_Operator_out845_out1;

  Logical_Operator_out1094_out1 <= Logical_Operator_out838_out1 XOR Logical_Operator_out846_out1;

  Logical_Operator_out1095_out1 <= Logical_Operator_out839_out1 XOR Logical_Operator_out847_out1;

  Logical_Operator_out1096_out1 <= Logical_Operator_out840_out1 XOR Logical_Operator_out848_out1;

  Logical_Operator_out1097_out1 <= Logical_Operator_out581_out1 XOR Logical_Operator_out589_out1;

  Logical_Operator_out1098_out1 <= Logical_Operator_out582_out1 XOR Logical_Operator_out590_out1;

  Logical_Operator_out1099_out1 <= Logical_Operator_out583_out1 XOR Logical_Operator_out591_out1;

  Logical_Operator_out1100_out1 <= Logical_Operator_out584_out1 XOR Logical_Operator_out592_out1;

  Logical_Operator_out1101_out1 <= Logical_Operator_out327_out1 XOR Logical_Operator_out335_out1;

  Logical_Operator_out1102_out1 <= Logical_Operator_out328_out1 XOR Logical_Operator_out336_out1;

  Logical_Operator_out1103_out1 <= Logical_Operator_out72_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out1104_out1 <= in144 XOR in160;

  Logical_Operator_out1105_out1 <= Logical_Operator_out849_out1 XOR Logical_Operator_out857_out1;

  Logical_Operator_out1106_out1 <= Logical_Operator_out850_out1 XOR Logical_Operator_out858_out1;

  Logical_Operator_out1107_out1 <= Logical_Operator_out851_out1 XOR Logical_Operator_out859_out1;

  Logical_Operator_out1108_out1 <= Logical_Operator_out852_out1 XOR Logical_Operator_out860_out1;

  Logical_Operator_out1109_out1 <= Logical_Operator_out853_out1 XOR Logical_Operator_out861_out1;

  Logical_Operator_out1110_out1 <= Logical_Operator_out854_out1 XOR Logical_Operator_out862_out1;

  Logical_Operator_out1111_out1 <= Logical_Operator_out855_out1 XOR Logical_Operator_out863_out1;

  Logical_Operator_out1112_out1 <= Logical_Operator_out856_out1 XOR Logical_Operator_out864_out1;

  Logical_Operator_out1113_out1 <= Logical_Operator_out597_out1 XOR Logical_Operator_out605_out1;

  Logical_Operator_out1114_out1 <= Logical_Operator_out598_out1 XOR Logical_Operator_out606_out1;

  Logical_Operator_out1115_out1 <= Logical_Operator_out599_out1 XOR Logical_Operator_out607_out1;

  Logical_Operator_out1116_out1 <= Logical_Operator_out600_out1 XOR Logical_Operator_out608_out1;

  Logical_Operator_out1117_out1 <= Logical_Operator_out343_out1 XOR Logical_Operator_out351_out1;

  Logical_Operator_out1118_out1 <= Logical_Operator_out344_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out1119_out1 <= Logical_Operator_out88_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out1120_out1 <= in176 XOR in192;

  Logical_Operator_out1121_out1 <= Logical_Operator_out865_out1 XOR Logical_Operator_out873_out1;

  Logical_Operator_out1122_out1 <= Logical_Operator_out866_out1 XOR Logical_Operator_out874_out1;

  Logical_Operator_out1123_out1 <= Logical_Operator_out867_out1 XOR Logical_Operator_out875_out1;

  Logical_Operator_out1124_out1 <= Logical_Operator_out868_out1 XOR Logical_Operator_out876_out1;

  Logical_Operator_out1125_out1 <= Logical_Operator_out869_out1 XOR Logical_Operator_out877_out1;

  Logical_Operator_out1126_out1 <= Logical_Operator_out870_out1 XOR Logical_Operator_out878_out1;

  Logical_Operator_out1127_out1 <= Logical_Operator_out871_out1 XOR Logical_Operator_out879_out1;

  Logical_Operator_out1128_out1 <= Logical_Operator_out872_out1 XOR Logical_Operator_out880_out1;

  Logical_Operator_out1129_out1 <= Logical_Operator_out613_out1 XOR Logical_Operator_out621_out1;

  Logical_Operator_out1130_out1 <= Logical_Operator_out614_out1 XOR Logical_Operator_out622_out1;

  Logical_Operator_out1131_out1 <= Logical_Operator_out615_out1 XOR Logical_Operator_out623_out1;

  Logical_Operator_out1132_out1 <= Logical_Operator_out616_out1 XOR Logical_Operator_out624_out1;

  Logical_Operator_out1133_out1 <= Logical_Operator_out359_out1 XOR Logical_Operator_out367_out1;

  Logical_Operator_out1134_out1 <= Logical_Operator_out360_out1 XOR Logical_Operator_out368_out1;

  Logical_Operator_out1135_out1 <= Logical_Operator_out104_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out1136_out1 <= in208 XOR in224;

  Logical_Operator_out1137_out1 <= Logical_Operator_out881_out1 XOR Logical_Operator_out889_out1;

  Logical_Operator_out1138_out1 <= Logical_Operator_out882_out1 XOR Logical_Operator_out890_out1;

  Logical_Operator_out1139_out1 <= Logical_Operator_out883_out1 XOR Logical_Operator_out891_out1;

  Logical_Operator_out1140_out1 <= Logical_Operator_out884_out1 XOR Logical_Operator_out892_out1;

  Logical_Operator_out1141_out1 <= Logical_Operator_out885_out1 XOR Logical_Operator_out893_out1;

  Logical_Operator_out1142_out1 <= Logical_Operator_out886_out1 XOR Logical_Operator_out894_out1;

  Logical_Operator_out1143_out1 <= Logical_Operator_out887_out1 XOR Logical_Operator_out895_out1;

  Logical_Operator_out1144_out1 <= Logical_Operator_out888_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out1145_out1 <= Logical_Operator_out629_out1 XOR Logical_Operator_out637_out1;

  Logical_Operator_out1146_out1 <= Logical_Operator_out630_out1 XOR Logical_Operator_out638_out1;

  Logical_Operator_out1147_out1 <= Logical_Operator_out631_out1 XOR Logical_Operator_out639_out1;

  Logical_Operator_out1148_out1 <= Logical_Operator_out632_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out1149_out1 <= Logical_Operator_out375_out1 XOR Logical_Operator_out383_out1;

  Logical_Operator_out1150_out1 <= Logical_Operator_out376_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out1151_out1 <= Logical_Operator_out120_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out1152_out1 <= in240 XOR in256;

  Logical_Operator_out1153_out1 <= Logical_Operator_out897_out1 XOR Logical_Operator_out905_out1;

  Logical_Operator_out1154_out1 <= Logical_Operator_out898_out1 XOR Logical_Operator_out906_out1;

  Logical_Operator_out1155_out1 <= Logical_Operator_out899_out1 XOR Logical_Operator_out907_out1;

  Logical_Operator_out1156_out1 <= Logical_Operator_out900_out1 XOR Logical_Operator_out908_out1;

  Logical_Operator_out1157_out1 <= Logical_Operator_out901_out1 XOR Logical_Operator_out909_out1;

  Logical_Operator_out1158_out1 <= Logical_Operator_out902_out1 XOR Logical_Operator_out910_out1;

  Logical_Operator_out1159_out1 <= Logical_Operator_out903_out1 XOR Logical_Operator_out911_out1;

  Logical_Operator_out1160_out1 <= Logical_Operator_out904_out1 XOR Logical_Operator_out912_out1;

  Logical_Operator_out1161_out1 <= Logical_Operator_out645_out1 XOR Logical_Operator_out653_out1;

  Logical_Operator_out1162_out1 <= Logical_Operator_out646_out1 XOR Logical_Operator_out654_out1;

  Logical_Operator_out1163_out1 <= Logical_Operator_out647_out1 XOR Logical_Operator_out655_out1;

  Logical_Operator_out1164_out1 <= Logical_Operator_out648_out1 XOR Logical_Operator_out656_out1;

  Logical_Operator_out1165_out1 <= Logical_Operator_out391_out1 XOR Logical_Operator_out399_out1;

  Logical_Operator_out1166_out1 <= Logical_Operator_out392_out1 XOR Logical_Operator_out400_out1;

  Logical_Operator_out1167_out1 <= Logical_Operator_out136_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out1168_out1 <= in272 XOR in288;

  Logical_Operator_out1169_out1 <= Logical_Operator_out913_out1 XOR Logical_Operator_out921_out1;

  Logical_Operator_out1170_out1 <= Logical_Operator_out914_out1 XOR Logical_Operator_out922_out1;

  Logical_Operator_out1171_out1 <= Logical_Operator_out915_out1 XOR Logical_Operator_out923_out1;

  Logical_Operator_out1172_out1 <= Logical_Operator_out916_out1 XOR Logical_Operator_out924_out1;

  Logical_Operator_out1173_out1 <= Logical_Operator_out917_out1 XOR Logical_Operator_out925_out1;

  Logical_Operator_out1174_out1 <= Logical_Operator_out918_out1 XOR Logical_Operator_out926_out1;

  Logical_Operator_out1175_out1 <= Logical_Operator_out919_out1 XOR Logical_Operator_out927_out1;

  Logical_Operator_out1176_out1 <= Logical_Operator_out920_out1 XOR Logical_Operator_out928_out1;

  Logical_Operator_out1177_out1 <= Logical_Operator_out661_out1 XOR Logical_Operator_out669_out1;

  Logical_Operator_out1178_out1 <= Logical_Operator_out662_out1 XOR Logical_Operator_out670_out1;

  Logical_Operator_out1179_out1 <= Logical_Operator_out663_out1 XOR Logical_Operator_out671_out1;

  Logical_Operator_out1180_out1 <= Logical_Operator_out664_out1 XOR Logical_Operator_out672_out1;

  Logical_Operator_out1181_out1 <= Logical_Operator_out407_out1 XOR Logical_Operator_out415_out1;

  Logical_Operator_out1182_out1 <= Logical_Operator_out408_out1 XOR Logical_Operator_out416_out1;

  Logical_Operator_out1183_out1 <= Logical_Operator_out152_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out1184_out1 <= in304 XOR in320;

  Logical_Operator_out1185_out1 <= Logical_Operator_out929_out1 XOR Logical_Operator_out937_out1;

  Logical_Operator_out1186_out1 <= Logical_Operator_out930_out1 XOR Logical_Operator_out938_out1;

  Logical_Operator_out1187_out1 <= Logical_Operator_out931_out1 XOR Logical_Operator_out939_out1;

  Logical_Operator_out1188_out1 <= Logical_Operator_out932_out1 XOR Logical_Operator_out940_out1;

  Logical_Operator_out1189_out1 <= Logical_Operator_out933_out1 XOR Logical_Operator_out941_out1;

  Logical_Operator_out1190_out1 <= Logical_Operator_out934_out1 XOR Logical_Operator_out942_out1;

  Logical_Operator_out1191_out1 <= Logical_Operator_out935_out1 XOR Logical_Operator_out943_out1;

  Logical_Operator_out1192_out1 <= Logical_Operator_out936_out1 XOR Logical_Operator_out944_out1;

  Logical_Operator_out1193_out1 <= Logical_Operator_out677_out1 XOR Logical_Operator_out685_out1;

  Logical_Operator_out1194_out1 <= Logical_Operator_out678_out1 XOR Logical_Operator_out686_out1;

  Logical_Operator_out1195_out1 <= Logical_Operator_out679_out1 XOR Logical_Operator_out687_out1;

  Logical_Operator_out1196_out1 <= Logical_Operator_out680_out1 XOR Logical_Operator_out688_out1;

  Logical_Operator_out1197_out1 <= Logical_Operator_out423_out1 XOR Logical_Operator_out431_out1;

  Logical_Operator_out1198_out1 <= Logical_Operator_out424_out1 XOR Logical_Operator_out432_out1;

  Logical_Operator_out1199_out1 <= Logical_Operator_out168_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out1200_out1 <= in336 XOR in352;

  Logical_Operator_out1201_out1 <= Logical_Operator_out945_out1 XOR Logical_Operator_out953_out1;

  Logical_Operator_out1202_out1 <= Logical_Operator_out946_out1 XOR Logical_Operator_out954_out1;

  Logical_Operator_out1203_out1 <= Logical_Operator_out947_out1 XOR Logical_Operator_out955_out1;

  Logical_Operator_out1204_out1 <= Logical_Operator_out948_out1 XOR Logical_Operator_out956_out1;

  Logical_Operator_out1205_out1 <= Logical_Operator_out949_out1 XOR Logical_Operator_out957_out1;

  Logical_Operator_out1206_out1 <= Logical_Operator_out950_out1 XOR Logical_Operator_out958_out1;

  Logical_Operator_out1207_out1 <= Logical_Operator_out951_out1 XOR Logical_Operator_out959_out1;

  Logical_Operator_out1208_out1 <= Logical_Operator_out952_out1 XOR Logical_Operator_out960_out1;

  Logical_Operator_out1209_out1 <= Logical_Operator_out693_out1 XOR Logical_Operator_out701_out1;

  Logical_Operator_out1210_out1 <= Logical_Operator_out694_out1 XOR Logical_Operator_out702_out1;

  Logical_Operator_out1211_out1 <= Logical_Operator_out695_out1 XOR Logical_Operator_out703_out1;

  Logical_Operator_out1212_out1 <= Logical_Operator_out696_out1 XOR Logical_Operator_out704_out1;

  Logical_Operator_out1213_out1 <= Logical_Operator_out439_out1 XOR Logical_Operator_out447_out1;

  Logical_Operator_out1214_out1 <= Logical_Operator_out440_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out1215_out1 <= Logical_Operator_out184_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out1216_out1 <= in368 XOR in384;

  Logical_Operator_out1217_out1 <= Logical_Operator_out961_out1 XOR Logical_Operator_out969_out1;

  Logical_Operator_out1218_out1 <= Logical_Operator_out962_out1 XOR Logical_Operator_out970_out1;

  Logical_Operator_out1219_out1 <= Logical_Operator_out963_out1 XOR Logical_Operator_out971_out1;

  Logical_Operator_out1220_out1 <= Logical_Operator_out964_out1 XOR Logical_Operator_out972_out1;

  Logical_Operator_out1221_out1 <= Logical_Operator_out965_out1 XOR Logical_Operator_out973_out1;

  Logical_Operator_out1222_out1 <= Logical_Operator_out966_out1 XOR Logical_Operator_out974_out1;

  Logical_Operator_out1223_out1 <= Logical_Operator_out967_out1 XOR Logical_Operator_out975_out1;

  Logical_Operator_out1224_out1 <= Logical_Operator_out968_out1 XOR Logical_Operator_out976_out1;

  Logical_Operator_out1225_out1 <= Logical_Operator_out709_out1 XOR Logical_Operator_out717_out1;

  Logical_Operator_out1226_out1 <= Logical_Operator_out710_out1 XOR Logical_Operator_out718_out1;

  Logical_Operator_out1227_out1 <= Logical_Operator_out711_out1 XOR Logical_Operator_out719_out1;

  Logical_Operator_out1228_out1 <= Logical_Operator_out712_out1 XOR Logical_Operator_out720_out1;

  Logical_Operator_out1229_out1 <= Logical_Operator_out455_out1 XOR Logical_Operator_out463_out1;

  Logical_Operator_out1230_out1 <= Logical_Operator_out456_out1 XOR Logical_Operator_out464_out1;

  Logical_Operator_out1231_out1 <= Logical_Operator_out200_out1 XOR Logical_Operator_out208_out1;

  Logical_Operator_out1232_out1 <= in400 XOR in416;

  Logical_Operator_out1233_out1 <= Logical_Operator_out977_out1 XOR Logical_Operator_out985_out1;

  Logical_Operator_out1234_out1 <= Logical_Operator_out978_out1 XOR Logical_Operator_out986_out1;

  Logical_Operator_out1235_out1 <= Logical_Operator_out979_out1 XOR Logical_Operator_out987_out1;

  Logical_Operator_out1236_out1 <= Logical_Operator_out980_out1 XOR Logical_Operator_out988_out1;

  Logical_Operator_out1237_out1 <= Logical_Operator_out981_out1 XOR Logical_Operator_out989_out1;

  Logical_Operator_out1238_out1 <= Logical_Operator_out982_out1 XOR Logical_Operator_out990_out1;

  Logical_Operator_out1239_out1 <= Logical_Operator_out983_out1 XOR Logical_Operator_out991_out1;

  Logical_Operator_out1240_out1 <= Logical_Operator_out984_out1 XOR Logical_Operator_out992_out1;

  Logical_Operator_out1241_out1 <= Logical_Operator_out725_out1 XOR Logical_Operator_out733_out1;

  Logical_Operator_out1242_out1 <= Logical_Operator_out726_out1 XOR Logical_Operator_out734_out1;

  Logical_Operator_out1243_out1 <= Logical_Operator_out727_out1 XOR Logical_Operator_out735_out1;

  Logical_Operator_out1244_out1 <= Logical_Operator_out728_out1 XOR Logical_Operator_out736_out1;

  Logical_Operator_out1245_out1 <= Logical_Operator_out471_out1 XOR Logical_Operator_out479_out1;

  Logical_Operator_out1246_out1 <= Logical_Operator_out472_out1 XOR Logical_Operator_out480_out1;

  Logical_Operator_out1247_out1 <= Logical_Operator_out216_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out1248_out1 <= in432 XOR in448;

  Logical_Operator_out1249_out1 <= Logical_Operator_out993_out1 XOR Logical_Operator_out1001_out1;

  Logical_Operator_out1250_out1 <= Logical_Operator_out994_out1 XOR Logical_Operator_out1002_out1;

  Logical_Operator_out1251_out1 <= Logical_Operator_out995_out1 XOR Logical_Operator_out1003_out1;

  Logical_Operator_out1252_out1 <= Logical_Operator_out996_out1 XOR Logical_Operator_out1004_out1;

  Logical_Operator_out1253_out1 <= Logical_Operator_out997_out1 XOR Logical_Operator_out1005_out1;

  Logical_Operator_out1254_out1 <= Logical_Operator_out998_out1 XOR Logical_Operator_out1006_out1;

  Logical_Operator_out1255_out1 <= Logical_Operator_out999_out1 XOR Logical_Operator_out1007_out1;

  Logical_Operator_out1256_out1 <= Logical_Operator_out1000_out1 XOR Logical_Operator_out1008_out1;

  Logical_Operator_out1257_out1 <= Logical_Operator_out741_out1 XOR Logical_Operator_out749_out1;

  Logical_Operator_out1258_out1 <= Logical_Operator_out742_out1 XOR Logical_Operator_out750_out1;

  Logical_Operator_out1259_out1 <= Logical_Operator_out743_out1 XOR Logical_Operator_out751_out1;

  Logical_Operator_out1260_out1 <= Logical_Operator_out744_out1 XOR Logical_Operator_out752_out1;

  Logical_Operator_out1261_out1 <= Logical_Operator_out487_out1 XOR Logical_Operator_out495_out1;

  Logical_Operator_out1262_out1 <= Logical_Operator_out488_out1 XOR Logical_Operator_out496_out1;

  Logical_Operator_out1263_out1 <= Logical_Operator_out232_out1 XOR Logical_Operator_out240_out1;

  Logical_Operator_out1264_out1 <= in464 XOR in480;

  Logical_Operator_out1265_out1 <= Logical_Operator_out1009_out1 XOR Logical_Operator_out1017_out1;

  Logical_Operator_out1266_out1 <= Logical_Operator_out1010_out1 XOR Logical_Operator_out1018_out1;

  Logical_Operator_out1267_out1 <= Logical_Operator_out1011_out1 XOR Logical_Operator_out1019_out1;

  Logical_Operator_out1268_out1 <= Logical_Operator_out1012_out1 XOR Logical_Operator_out1020_out1;

  Logical_Operator_out1269_out1 <= Logical_Operator_out1013_out1 XOR Logical_Operator_out1021_out1;

  Logical_Operator_out1270_out1 <= Logical_Operator_out1014_out1 XOR Logical_Operator_out1022_out1;

  Logical_Operator_out1271_out1 <= Logical_Operator_out1015_out1 XOR Logical_Operator_out1023_out1;

  Logical_Operator_out1272_out1 <= Logical_Operator_out1016_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out1273_out1 <= Logical_Operator_out757_out1 XOR Logical_Operator_out765_out1;

  Logical_Operator_out1274_out1 <= Logical_Operator_out758_out1 XOR Logical_Operator_out766_out1;

  Logical_Operator_out1275_out1 <= Logical_Operator_out759_out1 XOR Logical_Operator_out767_out1;

  Logical_Operator_out1276_out1 <= Logical_Operator_out760_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out1277_out1 <= Logical_Operator_out503_out1 XOR Logical_Operator_out511_out1;

  Logical_Operator_out1278_out1 <= Logical_Operator_out504_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out1279_out1 <= Logical_Operator_out248_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out1280_out1 <= in496 XOR in512;

  Logical_Operator_out1281_out1 <= Logical_Operator_out1025_out1 XOR Logical_Operator_out1041_out1;

  Logical_Operator_out1282_out1 <= Logical_Operator_out1026_out1 XOR Logical_Operator_out1042_out1;

  Logical_Operator_out1283_out1 <= Logical_Operator_out1027_out1 XOR Logical_Operator_out1043_out1;

  Logical_Operator_out1284_out1 <= Logical_Operator_out1028_out1 XOR Logical_Operator_out1044_out1;

  Logical_Operator_out1285_out1 <= Logical_Operator_out1029_out1 XOR Logical_Operator_out1045_out1;

  Logical_Operator_out1286_out1 <= Logical_Operator_out1030_out1 XOR Logical_Operator_out1046_out1;

  Logical_Operator_out1287_out1 <= Logical_Operator_out1031_out1 XOR Logical_Operator_out1047_out1;

  Logical_Operator_out1288_out1 <= Logical_Operator_out1032_out1 XOR Logical_Operator_out1048_out1;

  Logical_Operator_out1289_out1 <= Logical_Operator_out1033_out1 XOR Logical_Operator_out1049_out1;

  Logical_Operator_out1290_out1 <= Logical_Operator_out1034_out1 XOR Logical_Operator_out1050_out1;

  Logical_Operator_out1291_out1 <= Logical_Operator_out1035_out1 XOR Logical_Operator_out1051_out1;

  Logical_Operator_out1292_out1 <= Logical_Operator_out1036_out1 XOR Logical_Operator_out1052_out1;

  Logical_Operator_out1293_out1 <= Logical_Operator_out1037_out1 XOR Logical_Operator_out1053_out1;

  Logical_Operator_out1294_out1 <= Logical_Operator_out1038_out1 XOR Logical_Operator_out1054_out1;

  Logical_Operator_out1295_out1 <= Logical_Operator_out1039_out1 XOR Logical_Operator_out1055_out1;

  Logical_Operator_out1296_out1 <= Logical_Operator_out1040_out1 XOR Logical_Operator_out1056_out1;

  Logical_Operator_out1297_out1 <= Logical_Operator_out777_out1 XOR Logical_Operator_out793_out1;

  Logical_Operator_out1298_out1 <= Logical_Operator_out778_out1 XOR Logical_Operator_out794_out1;

  Logical_Operator_out1299_out1 <= Logical_Operator_out779_out1 XOR Logical_Operator_out795_out1;

  Logical_Operator_out1300_out1 <= Logical_Operator_out780_out1 XOR Logical_Operator_out796_out1;

  Logical_Operator_out1301_out1 <= Logical_Operator_out781_out1 XOR Logical_Operator_out797_out1;

  Logical_Operator_out1302_out1 <= Logical_Operator_out782_out1 XOR Logical_Operator_out798_out1;

  Logical_Operator_out1303_out1 <= Logical_Operator_out783_out1 XOR Logical_Operator_out799_out1;

  Logical_Operator_out1304_out1 <= Logical_Operator_out784_out1 XOR Logical_Operator_out800_out1;

  Logical_Operator_out1305_out1 <= Logical_Operator_out525_out1 XOR Logical_Operator_out541_out1;

  Logical_Operator_out1306_out1 <= Logical_Operator_out526_out1 XOR Logical_Operator_out542_out1;

  Logical_Operator_out1307_out1 <= Logical_Operator_out527_out1 XOR Logical_Operator_out543_out1;

  Logical_Operator_out1308_out1 <= Logical_Operator_out528_out1 XOR Logical_Operator_out544_out1;

  Logical_Operator_out1309_out1 <= Logical_Operator_out271_out1 XOR Logical_Operator_out287_out1;

  Logical_Operator_out1310_out1 <= Logical_Operator_out272_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out1311_out1 <= Logical_Operator_out16_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out1312_out1 <= in32 XOR in64;

  Logical_Operator_out1313_out1 <= Logical_Operator_out1057_out1 XOR Logical_Operator_out1073_out1;

  Logical_Operator_out1314_out1 <= Logical_Operator_out1058_out1 XOR Logical_Operator_out1074_out1;

  Logical_Operator_out1315_out1 <= Logical_Operator_out1059_out1 XOR Logical_Operator_out1075_out1;

  Logical_Operator_out1316_out1 <= Logical_Operator_out1060_out1 XOR Logical_Operator_out1076_out1;

  Logical_Operator_out1317_out1 <= Logical_Operator_out1061_out1 XOR Logical_Operator_out1077_out1;

  Logical_Operator_out1318_out1 <= Logical_Operator_out1062_out1 XOR Logical_Operator_out1078_out1;

  Logical_Operator_out1319_out1 <= Logical_Operator_out1063_out1 XOR Logical_Operator_out1079_out1;

  Logical_Operator_out1320_out1 <= Logical_Operator_out1064_out1 XOR Logical_Operator_out1080_out1;

  Logical_Operator_out1321_out1 <= Logical_Operator_out1065_out1 XOR Logical_Operator_out1081_out1;

  Logical_Operator_out1322_out1 <= Logical_Operator_out1066_out1 XOR Logical_Operator_out1082_out1;

  Logical_Operator_out1323_out1 <= Logical_Operator_out1067_out1 XOR Logical_Operator_out1083_out1;

  Logical_Operator_out1324_out1 <= Logical_Operator_out1068_out1 XOR Logical_Operator_out1084_out1;

  Logical_Operator_out1325_out1 <= Logical_Operator_out1069_out1 XOR Logical_Operator_out1085_out1;

  Logical_Operator_out1326_out1 <= Logical_Operator_out1070_out1 XOR Logical_Operator_out1086_out1;

  Logical_Operator_out1327_out1 <= Logical_Operator_out1071_out1 XOR Logical_Operator_out1087_out1;

  Logical_Operator_out1328_out1 <= Logical_Operator_out1072_out1 XOR Logical_Operator_out1088_out1;

  Logical_Operator_out1329_out1 <= Logical_Operator_out809_out1 XOR Logical_Operator_out825_out1;

  Logical_Operator_out1330_out1 <= Logical_Operator_out810_out1 XOR Logical_Operator_out826_out1;

  Logical_Operator_out1331_out1 <= Logical_Operator_out811_out1 XOR Logical_Operator_out827_out1;

  Logical_Operator_out1332_out1 <= Logical_Operator_out812_out1 XOR Logical_Operator_out828_out1;

  Logical_Operator_out1333_out1 <= Logical_Operator_out813_out1 XOR Logical_Operator_out829_out1;

  Logical_Operator_out1334_out1 <= Logical_Operator_out814_out1 XOR Logical_Operator_out830_out1;

  Logical_Operator_out1335_out1 <= Logical_Operator_out815_out1 XOR Logical_Operator_out831_out1;

  Logical_Operator_out1336_out1 <= Logical_Operator_out816_out1 XOR Logical_Operator_out832_out1;

  Logical_Operator_out1337_out1 <= Logical_Operator_out557_out1 XOR Logical_Operator_out573_out1;

  Logical_Operator_out1338_out1 <= Logical_Operator_out558_out1 XOR Logical_Operator_out574_out1;

  Logical_Operator_out1339_out1 <= Logical_Operator_out559_out1 XOR Logical_Operator_out575_out1;

  Logical_Operator_out1340_out1 <= Logical_Operator_out560_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out1341_out1 <= Logical_Operator_out303_out1 XOR Logical_Operator_out319_out1;

  Logical_Operator_out1342_out1 <= Logical_Operator_out304_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out1343_out1 <= Logical_Operator_out48_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out1344_out1 <= in96 XOR in128;

  Logical_Operator_out1345_out1 <= Logical_Operator_out1089_out1 XOR Logical_Operator_out1105_out1;

  Logical_Operator_out1346_out1 <= Logical_Operator_out1090_out1 XOR Logical_Operator_out1106_out1;

  Logical_Operator_out1347_out1 <= Logical_Operator_out1091_out1 XOR Logical_Operator_out1107_out1;

  Logical_Operator_out1348_out1 <= Logical_Operator_out1092_out1 XOR Logical_Operator_out1108_out1;

  Logical_Operator_out1349_out1 <= Logical_Operator_out1093_out1 XOR Logical_Operator_out1109_out1;

  Logical_Operator_out1350_out1 <= Logical_Operator_out1094_out1 XOR Logical_Operator_out1110_out1;

  Logical_Operator_out1351_out1 <= Logical_Operator_out1095_out1 XOR Logical_Operator_out1111_out1;

  Logical_Operator_out1352_out1 <= Logical_Operator_out1096_out1 XOR Logical_Operator_out1112_out1;

  Logical_Operator_out1353_out1 <= Logical_Operator_out1097_out1 XOR Logical_Operator_out1113_out1;

  Logical_Operator_out1354_out1 <= Logical_Operator_out1098_out1 XOR Logical_Operator_out1114_out1;

  Logical_Operator_out1355_out1 <= Logical_Operator_out1099_out1 XOR Logical_Operator_out1115_out1;

  Logical_Operator_out1356_out1 <= Logical_Operator_out1100_out1 XOR Logical_Operator_out1116_out1;

  Logical_Operator_out1357_out1 <= Logical_Operator_out1101_out1 XOR Logical_Operator_out1117_out1;

  Logical_Operator_out1358_out1 <= Logical_Operator_out1102_out1 XOR Logical_Operator_out1118_out1;

  Logical_Operator_out1359_out1 <= Logical_Operator_out1103_out1 XOR Logical_Operator_out1119_out1;

  Logical_Operator_out1360_out1 <= Logical_Operator_out1104_out1 XOR Logical_Operator_out1120_out1;

  Logical_Operator_out1361_out1 <= Logical_Operator_out841_out1 XOR Logical_Operator_out857_out1;

  Logical_Operator_out1362_out1 <= Logical_Operator_out842_out1 XOR Logical_Operator_out858_out1;

  Logical_Operator_out1363_out1 <= Logical_Operator_out843_out1 XOR Logical_Operator_out859_out1;

  Logical_Operator_out1364_out1 <= Logical_Operator_out844_out1 XOR Logical_Operator_out860_out1;

  Logical_Operator_out1365_out1 <= Logical_Operator_out845_out1 XOR Logical_Operator_out861_out1;

  Logical_Operator_out1366_out1 <= Logical_Operator_out846_out1 XOR Logical_Operator_out862_out1;

  Logical_Operator_out1367_out1 <= Logical_Operator_out847_out1 XOR Logical_Operator_out863_out1;

  Logical_Operator_out1368_out1 <= Logical_Operator_out848_out1 XOR Logical_Operator_out864_out1;

  Logical_Operator_out1369_out1 <= Logical_Operator_out589_out1 XOR Logical_Operator_out605_out1;

  Logical_Operator_out1370_out1 <= Logical_Operator_out590_out1 XOR Logical_Operator_out606_out1;

  Logical_Operator_out1371_out1 <= Logical_Operator_out591_out1 XOR Logical_Operator_out607_out1;

  Logical_Operator_out1372_out1 <= Logical_Operator_out592_out1 XOR Logical_Operator_out608_out1;

  Logical_Operator_out1373_out1 <= Logical_Operator_out335_out1 XOR Logical_Operator_out351_out1;

  Logical_Operator_out1374_out1 <= Logical_Operator_out336_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out1375_out1 <= Logical_Operator_out80_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out1376_out1 <= in160 XOR in192;

  Logical_Operator_out1377_out1 <= Logical_Operator_out1121_out1 XOR Logical_Operator_out1137_out1;

  Logical_Operator_out1378_out1 <= Logical_Operator_out1122_out1 XOR Logical_Operator_out1138_out1;

  Logical_Operator_out1379_out1 <= Logical_Operator_out1123_out1 XOR Logical_Operator_out1139_out1;

  Logical_Operator_out1380_out1 <= Logical_Operator_out1124_out1 XOR Logical_Operator_out1140_out1;

  Logical_Operator_out1381_out1 <= Logical_Operator_out1125_out1 XOR Logical_Operator_out1141_out1;

  Logical_Operator_out1382_out1 <= Logical_Operator_out1126_out1 XOR Logical_Operator_out1142_out1;

  Logical_Operator_out1383_out1 <= Logical_Operator_out1127_out1 XOR Logical_Operator_out1143_out1;

  Logical_Operator_out1384_out1 <= Logical_Operator_out1128_out1 XOR Logical_Operator_out1144_out1;

  Logical_Operator_out1385_out1 <= Logical_Operator_out1129_out1 XOR Logical_Operator_out1145_out1;

  Logical_Operator_out1386_out1 <= Logical_Operator_out1130_out1 XOR Logical_Operator_out1146_out1;

  Logical_Operator_out1387_out1 <= Logical_Operator_out1131_out1 XOR Logical_Operator_out1147_out1;

  Logical_Operator_out1388_out1 <= Logical_Operator_out1132_out1 XOR Logical_Operator_out1148_out1;

  Logical_Operator_out1389_out1 <= Logical_Operator_out1133_out1 XOR Logical_Operator_out1149_out1;

  Logical_Operator_out1390_out1 <= Logical_Operator_out1134_out1 XOR Logical_Operator_out1150_out1;

  Logical_Operator_out1391_out1 <= Logical_Operator_out1135_out1 XOR Logical_Operator_out1151_out1;

  Logical_Operator_out1392_out1 <= Logical_Operator_out1136_out1 XOR Logical_Operator_out1152_out1;

  Logical_Operator_out1393_out1 <= Logical_Operator_out873_out1 XOR Logical_Operator_out889_out1;

  Logical_Operator_out1394_out1 <= Logical_Operator_out874_out1 XOR Logical_Operator_out890_out1;

  Logical_Operator_out1395_out1 <= Logical_Operator_out875_out1 XOR Logical_Operator_out891_out1;

  Logical_Operator_out1396_out1 <= Logical_Operator_out876_out1 XOR Logical_Operator_out892_out1;

  Logical_Operator_out1397_out1 <= Logical_Operator_out877_out1 XOR Logical_Operator_out893_out1;

  Logical_Operator_out1398_out1 <= Logical_Operator_out878_out1 XOR Logical_Operator_out894_out1;

  Logical_Operator_out1399_out1 <= Logical_Operator_out879_out1 XOR Logical_Operator_out895_out1;

  Logical_Operator_out1400_out1 <= Logical_Operator_out880_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out1401_out1 <= Logical_Operator_out621_out1 XOR Logical_Operator_out637_out1;

  Logical_Operator_out1402_out1 <= Logical_Operator_out622_out1 XOR Logical_Operator_out638_out1;

  Logical_Operator_out1403_out1 <= Logical_Operator_out623_out1 XOR Logical_Operator_out639_out1;

  Logical_Operator_out1404_out1 <= Logical_Operator_out624_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out1405_out1 <= Logical_Operator_out367_out1 XOR Logical_Operator_out383_out1;

  Logical_Operator_out1406_out1 <= Logical_Operator_out368_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out1407_out1 <= Logical_Operator_out112_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out1408_out1 <= in224 XOR in256;

  Logical_Operator_out1409_out1 <= Logical_Operator_out1153_out1 XOR Logical_Operator_out1169_out1;

  Logical_Operator_out1410_out1 <= Logical_Operator_out1154_out1 XOR Logical_Operator_out1170_out1;

  Logical_Operator_out1411_out1 <= Logical_Operator_out1155_out1 XOR Logical_Operator_out1171_out1;

  Logical_Operator_out1412_out1 <= Logical_Operator_out1156_out1 XOR Logical_Operator_out1172_out1;

  Logical_Operator_out1413_out1 <= Logical_Operator_out1157_out1 XOR Logical_Operator_out1173_out1;

  Logical_Operator_out1414_out1 <= Logical_Operator_out1158_out1 XOR Logical_Operator_out1174_out1;

  Logical_Operator_out1415_out1 <= Logical_Operator_out1159_out1 XOR Logical_Operator_out1175_out1;

  Logical_Operator_out1416_out1 <= Logical_Operator_out1160_out1 XOR Logical_Operator_out1176_out1;

  Logical_Operator_out1417_out1 <= Logical_Operator_out1161_out1 XOR Logical_Operator_out1177_out1;

  Logical_Operator_out1418_out1 <= Logical_Operator_out1162_out1 XOR Logical_Operator_out1178_out1;

  Logical_Operator_out1419_out1 <= Logical_Operator_out1163_out1 XOR Logical_Operator_out1179_out1;

  Logical_Operator_out1420_out1 <= Logical_Operator_out1164_out1 XOR Logical_Operator_out1180_out1;

  Logical_Operator_out1421_out1 <= Logical_Operator_out1165_out1 XOR Logical_Operator_out1181_out1;

  Logical_Operator_out1422_out1 <= Logical_Operator_out1166_out1 XOR Logical_Operator_out1182_out1;

  Logical_Operator_out1423_out1 <= Logical_Operator_out1167_out1 XOR Logical_Operator_out1183_out1;

  Logical_Operator_out1424_out1 <= Logical_Operator_out1168_out1 XOR Logical_Operator_out1184_out1;

  Logical_Operator_out1425_out1 <= Logical_Operator_out905_out1 XOR Logical_Operator_out921_out1;

  Logical_Operator_out1426_out1 <= Logical_Operator_out906_out1 XOR Logical_Operator_out922_out1;

  Logical_Operator_out1427_out1 <= Logical_Operator_out907_out1 XOR Logical_Operator_out923_out1;

  Logical_Operator_out1428_out1 <= Logical_Operator_out908_out1 XOR Logical_Operator_out924_out1;

  Logical_Operator_out1429_out1 <= Logical_Operator_out909_out1 XOR Logical_Operator_out925_out1;

  Logical_Operator_out1430_out1 <= Logical_Operator_out910_out1 XOR Logical_Operator_out926_out1;

  Logical_Operator_out1431_out1 <= Logical_Operator_out911_out1 XOR Logical_Operator_out927_out1;

  Logical_Operator_out1432_out1 <= Logical_Operator_out912_out1 XOR Logical_Operator_out928_out1;

  Logical_Operator_out1433_out1 <= Logical_Operator_out653_out1 XOR Logical_Operator_out669_out1;

  Logical_Operator_out1434_out1 <= Logical_Operator_out654_out1 XOR Logical_Operator_out670_out1;

  Logical_Operator_out1435_out1 <= Logical_Operator_out655_out1 XOR Logical_Operator_out671_out1;

  Logical_Operator_out1436_out1 <= Logical_Operator_out656_out1 XOR Logical_Operator_out672_out1;

  Logical_Operator_out1437_out1 <= Logical_Operator_out399_out1 XOR Logical_Operator_out415_out1;

  Logical_Operator_out1438_out1 <= Logical_Operator_out400_out1 XOR Logical_Operator_out416_out1;

  Logical_Operator_out1439_out1 <= Logical_Operator_out144_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out1440_out1 <= in288 XOR in320;

  Logical_Operator_out1441_out1 <= Logical_Operator_out1185_out1 XOR Logical_Operator_out1201_out1;

  Logical_Operator_out1442_out1 <= Logical_Operator_out1186_out1 XOR Logical_Operator_out1202_out1;

  Logical_Operator_out1443_out1 <= Logical_Operator_out1187_out1 XOR Logical_Operator_out1203_out1;

  Logical_Operator_out1444_out1 <= Logical_Operator_out1188_out1 XOR Logical_Operator_out1204_out1;

  Logical_Operator_out1445_out1 <= Logical_Operator_out1189_out1 XOR Logical_Operator_out1205_out1;

  Logical_Operator_out1446_out1 <= Logical_Operator_out1190_out1 XOR Logical_Operator_out1206_out1;

  Logical_Operator_out1447_out1 <= Logical_Operator_out1191_out1 XOR Logical_Operator_out1207_out1;

  Logical_Operator_out1448_out1 <= Logical_Operator_out1192_out1 XOR Logical_Operator_out1208_out1;

  Logical_Operator_out1449_out1 <= Logical_Operator_out1193_out1 XOR Logical_Operator_out1209_out1;

  Logical_Operator_out1450_out1 <= Logical_Operator_out1194_out1 XOR Logical_Operator_out1210_out1;

  Logical_Operator_out1451_out1 <= Logical_Operator_out1195_out1 XOR Logical_Operator_out1211_out1;

  Logical_Operator_out1452_out1 <= Logical_Operator_out1196_out1 XOR Logical_Operator_out1212_out1;

  Logical_Operator_out1453_out1 <= Logical_Operator_out1197_out1 XOR Logical_Operator_out1213_out1;

  Logical_Operator_out1454_out1 <= Logical_Operator_out1198_out1 XOR Logical_Operator_out1214_out1;

  Logical_Operator_out1455_out1 <= Logical_Operator_out1199_out1 XOR Logical_Operator_out1215_out1;

  Logical_Operator_out1456_out1 <= Logical_Operator_out1200_out1 XOR Logical_Operator_out1216_out1;

  Logical_Operator_out1457_out1 <= Logical_Operator_out937_out1 XOR Logical_Operator_out953_out1;

  Logical_Operator_out1458_out1 <= Logical_Operator_out938_out1 XOR Logical_Operator_out954_out1;

  Logical_Operator_out1459_out1 <= Logical_Operator_out939_out1 XOR Logical_Operator_out955_out1;

  Logical_Operator_out1460_out1 <= Logical_Operator_out940_out1 XOR Logical_Operator_out956_out1;

  Logical_Operator_out1461_out1 <= Logical_Operator_out941_out1 XOR Logical_Operator_out957_out1;

  Logical_Operator_out1462_out1 <= Logical_Operator_out942_out1 XOR Logical_Operator_out958_out1;

  Logical_Operator_out1463_out1 <= Logical_Operator_out943_out1 XOR Logical_Operator_out959_out1;

  Logical_Operator_out1464_out1 <= Logical_Operator_out944_out1 XOR Logical_Operator_out960_out1;

  Logical_Operator_out1465_out1 <= Logical_Operator_out685_out1 XOR Logical_Operator_out701_out1;

  Logical_Operator_out1466_out1 <= Logical_Operator_out686_out1 XOR Logical_Operator_out702_out1;

  Logical_Operator_out1467_out1 <= Logical_Operator_out687_out1 XOR Logical_Operator_out703_out1;

  Logical_Operator_out1468_out1 <= Logical_Operator_out688_out1 XOR Logical_Operator_out704_out1;

  Logical_Operator_out1469_out1 <= Logical_Operator_out431_out1 XOR Logical_Operator_out447_out1;

  Logical_Operator_out1470_out1 <= Logical_Operator_out432_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out1471_out1 <= Logical_Operator_out176_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out1472_out1 <= in352 XOR in384;

  Logical_Operator_out1473_out1 <= Logical_Operator_out1217_out1 XOR Logical_Operator_out1233_out1;

  Logical_Operator_out1474_out1 <= Logical_Operator_out1218_out1 XOR Logical_Operator_out1234_out1;

  Logical_Operator_out1475_out1 <= Logical_Operator_out1219_out1 XOR Logical_Operator_out1235_out1;

  Logical_Operator_out1476_out1 <= Logical_Operator_out1220_out1 XOR Logical_Operator_out1236_out1;

  Logical_Operator_out1477_out1 <= Logical_Operator_out1221_out1 XOR Logical_Operator_out1237_out1;

  Logical_Operator_out1478_out1 <= Logical_Operator_out1222_out1 XOR Logical_Operator_out1238_out1;

  Logical_Operator_out1479_out1 <= Logical_Operator_out1223_out1 XOR Logical_Operator_out1239_out1;

  Logical_Operator_out1480_out1 <= Logical_Operator_out1224_out1 XOR Logical_Operator_out1240_out1;

  Logical_Operator_out1481_out1 <= Logical_Operator_out1225_out1 XOR Logical_Operator_out1241_out1;

  Logical_Operator_out1482_out1 <= Logical_Operator_out1226_out1 XOR Logical_Operator_out1242_out1;

  Logical_Operator_out1483_out1 <= Logical_Operator_out1227_out1 XOR Logical_Operator_out1243_out1;

  Logical_Operator_out1484_out1 <= Logical_Operator_out1228_out1 XOR Logical_Operator_out1244_out1;

  Logical_Operator_out1485_out1 <= Logical_Operator_out1229_out1 XOR Logical_Operator_out1245_out1;

  Logical_Operator_out1486_out1 <= Logical_Operator_out1230_out1 XOR Logical_Operator_out1246_out1;

  Logical_Operator_out1487_out1 <= Logical_Operator_out1231_out1 XOR Logical_Operator_out1247_out1;

  Logical_Operator_out1488_out1 <= Logical_Operator_out1232_out1 XOR Logical_Operator_out1248_out1;

  Logical_Operator_out1489_out1 <= Logical_Operator_out969_out1 XOR Logical_Operator_out985_out1;

  Logical_Operator_out1490_out1 <= Logical_Operator_out970_out1 XOR Logical_Operator_out986_out1;

  Logical_Operator_out1491_out1 <= Logical_Operator_out971_out1 XOR Logical_Operator_out987_out1;

  Logical_Operator_out1492_out1 <= Logical_Operator_out972_out1 XOR Logical_Operator_out988_out1;

  Logical_Operator_out1493_out1 <= Logical_Operator_out973_out1 XOR Logical_Operator_out989_out1;

  Logical_Operator_out1494_out1 <= Logical_Operator_out974_out1 XOR Logical_Operator_out990_out1;

  Logical_Operator_out1495_out1 <= Logical_Operator_out975_out1 XOR Logical_Operator_out991_out1;

  Logical_Operator_out1496_out1 <= Logical_Operator_out976_out1 XOR Logical_Operator_out992_out1;

  Logical_Operator_out1497_out1 <= Logical_Operator_out717_out1 XOR Logical_Operator_out733_out1;

  Logical_Operator_out1498_out1 <= Logical_Operator_out718_out1 XOR Logical_Operator_out734_out1;

  Logical_Operator_out1499_out1 <= Logical_Operator_out719_out1 XOR Logical_Operator_out735_out1;

  Logical_Operator_out1500_out1 <= Logical_Operator_out720_out1 XOR Logical_Operator_out736_out1;

  Logical_Operator_out1501_out1 <= Logical_Operator_out463_out1 XOR Logical_Operator_out479_out1;

  Logical_Operator_out1502_out1 <= Logical_Operator_out464_out1 XOR Logical_Operator_out480_out1;

  Logical_Operator_out1503_out1 <= Logical_Operator_out208_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out1504_out1 <= in416 XOR in448;

  Logical_Operator_out1505_out1 <= Logical_Operator_out1249_out1 XOR Logical_Operator_out1265_out1;

  Logical_Operator_out1506_out1 <= Logical_Operator_out1250_out1 XOR Logical_Operator_out1266_out1;

  Logical_Operator_out1507_out1 <= Logical_Operator_out1251_out1 XOR Logical_Operator_out1267_out1;

  Logical_Operator_out1508_out1 <= Logical_Operator_out1252_out1 XOR Logical_Operator_out1268_out1;

  Logical_Operator_out1509_out1 <= Logical_Operator_out1253_out1 XOR Logical_Operator_out1269_out1;

  Logical_Operator_out1510_out1 <= Logical_Operator_out1254_out1 XOR Logical_Operator_out1270_out1;

  Logical_Operator_out1511_out1 <= Logical_Operator_out1255_out1 XOR Logical_Operator_out1271_out1;

  Logical_Operator_out1512_out1 <= Logical_Operator_out1256_out1 XOR Logical_Operator_out1272_out1;

  Logical_Operator_out1513_out1 <= Logical_Operator_out1257_out1 XOR Logical_Operator_out1273_out1;

  Logical_Operator_out1514_out1 <= Logical_Operator_out1258_out1 XOR Logical_Operator_out1274_out1;

  Logical_Operator_out1515_out1 <= Logical_Operator_out1259_out1 XOR Logical_Operator_out1275_out1;

  Logical_Operator_out1516_out1 <= Logical_Operator_out1260_out1 XOR Logical_Operator_out1276_out1;

  Logical_Operator_out1517_out1 <= Logical_Operator_out1261_out1 XOR Logical_Operator_out1277_out1;

  Logical_Operator_out1518_out1 <= Logical_Operator_out1262_out1 XOR Logical_Operator_out1278_out1;

  Logical_Operator_out1519_out1 <= Logical_Operator_out1263_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out1520_out1 <= Logical_Operator_out1264_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out1521_out1 <= Logical_Operator_out1001_out1 XOR Logical_Operator_out1017_out1;

  Logical_Operator_out1522_out1 <= Logical_Operator_out1002_out1 XOR Logical_Operator_out1018_out1;

  Logical_Operator_out1523_out1 <= Logical_Operator_out1003_out1 XOR Logical_Operator_out1019_out1;

  Logical_Operator_out1524_out1 <= Logical_Operator_out1004_out1 XOR Logical_Operator_out1020_out1;

  Logical_Operator_out1525_out1 <= Logical_Operator_out1005_out1 XOR Logical_Operator_out1021_out1;

  Logical_Operator_out1526_out1 <= Logical_Operator_out1006_out1 XOR Logical_Operator_out1022_out1;

  Logical_Operator_out1527_out1 <= Logical_Operator_out1007_out1 XOR Logical_Operator_out1023_out1;

  Logical_Operator_out1528_out1 <= Logical_Operator_out1008_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out1529_out1 <= Logical_Operator_out749_out1 XOR Logical_Operator_out765_out1;

  Logical_Operator_out1530_out1 <= Logical_Operator_out750_out1 XOR Logical_Operator_out766_out1;

  Logical_Operator_out1531_out1 <= Logical_Operator_out751_out1 XOR Logical_Operator_out767_out1;

  Logical_Operator_out1532_out1 <= Logical_Operator_out752_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out1533_out1 <= Logical_Operator_out495_out1 XOR Logical_Operator_out511_out1;

  Logical_Operator_out1534_out1 <= Logical_Operator_out496_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out1535_out1 <= Logical_Operator_out240_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out1536_out1 <= in480 XOR in512;

  Logical_Operator_out1537_out1 <= Logical_Operator_out1281_out1 XOR Logical_Operator_out1313_out1;

  Logical_Operator_out1538_out1 <= Logical_Operator_out1282_out1 XOR Logical_Operator_out1314_out1;

  Logical_Operator_out1539_out1 <= Logical_Operator_out1283_out1 XOR Logical_Operator_out1315_out1;

  Logical_Operator_out1540_out1 <= Logical_Operator_out1284_out1 XOR Logical_Operator_out1316_out1;

  Logical_Operator_out1541_out1 <= Logical_Operator_out1285_out1 XOR Logical_Operator_out1317_out1;

  Logical_Operator_out1542_out1 <= Logical_Operator_out1286_out1 XOR Logical_Operator_out1318_out1;

  Logical_Operator_out1543_out1 <= Logical_Operator_out1287_out1 XOR Logical_Operator_out1319_out1;

  Logical_Operator_out1544_out1 <= Logical_Operator_out1288_out1 XOR Logical_Operator_out1320_out1;

  Logical_Operator_out1545_out1 <= Logical_Operator_out1289_out1 XOR Logical_Operator_out1321_out1;

  Logical_Operator_out1546_out1 <= Logical_Operator_out1290_out1 XOR Logical_Operator_out1322_out1;

  Logical_Operator_out1547_out1 <= Logical_Operator_out1291_out1 XOR Logical_Operator_out1323_out1;

  Logical_Operator_out1548_out1 <= Logical_Operator_out1292_out1 XOR Logical_Operator_out1324_out1;

  Logical_Operator_out1549_out1 <= Logical_Operator_out1293_out1 XOR Logical_Operator_out1325_out1;

  Logical_Operator_out1550_out1 <= Logical_Operator_out1294_out1 XOR Logical_Operator_out1326_out1;

  Logical_Operator_out1551_out1 <= Logical_Operator_out1295_out1 XOR Logical_Operator_out1327_out1;

  Logical_Operator_out1552_out1 <= Logical_Operator_out1296_out1 XOR Logical_Operator_out1328_out1;

  Logical_Operator_out1553_out1 <= Logical_Operator_out1297_out1 XOR Logical_Operator_out1329_out1;

  Logical_Operator_out1554_out1 <= Logical_Operator_out1298_out1 XOR Logical_Operator_out1330_out1;

  Logical_Operator_out1555_out1 <= Logical_Operator_out1299_out1 XOR Logical_Operator_out1331_out1;

  Logical_Operator_out1556_out1 <= Logical_Operator_out1300_out1 XOR Logical_Operator_out1332_out1;

  Logical_Operator_out1557_out1 <= Logical_Operator_out1301_out1 XOR Logical_Operator_out1333_out1;

  Logical_Operator_out1558_out1 <= Logical_Operator_out1302_out1 XOR Logical_Operator_out1334_out1;

  Logical_Operator_out1559_out1 <= Logical_Operator_out1303_out1 XOR Logical_Operator_out1335_out1;

  Logical_Operator_out1560_out1 <= Logical_Operator_out1304_out1 XOR Logical_Operator_out1336_out1;

  Logical_Operator_out1561_out1 <= Logical_Operator_out1305_out1 XOR Logical_Operator_out1337_out1;

  Logical_Operator_out1562_out1 <= Logical_Operator_out1306_out1 XOR Logical_Operator_out1338_out1;

  Logical_Operator_out1563_out1 <= Logical_Operator_out1307_out1 XOR Logical_Operator_out1339_out1;

  Logical_Operator_out1564_out1 <= Logical_Operator_out1308_out1 XOR Logical_Operator_out1340_out1;

  Logical_Operator_out1565_out1 <= Logical_Operator_out1309_out1 XOR Logical_Operator_out1341_out1;

  Logical_Operator_out1566_out1 <= Logical_Operator_out1310_out1 XOR Logical_Operator_out1342_out1;

  Logical_Operator_out1567_out1 <= Logical_Operator_out1311_out1 XOR Logical_Operator_out1343_out1;

  Logical_Operator_out1568_out1 <= Logical_Operator_out1312_out1 XOR Logical_Operator_out1344_out1;

  Logical_Operator_out1569_out1 <= Logical_Operator_out1041_out1 XOR Logical_Operator_out1073_out1;

  Logical_Operator_out1570_out1 <= Logical_Operator_out1042_out1 XOR Logical_Operator_out1074_out1;

  Logical_Operator_out1571_out1 <= Logical_Operator_out1043_out1 XOR Logical_Operator_out1075_out1;

  Logical_Operator_out1572_out1 <= Logical_Operator_out1044_out1 XOR Logical_Operator_out1076_out1;

  Logical_Operator_out1573_out1 <= Logical_Operator_out1045_out1 XOR Logical_Operator_out1077_out1;

  Logical_Operator_out1574_out1 <= Logical_Operator_out1046_out1 XOR Logical_Operator_out1078_out1;

  Logical_Operator_out1575_out1 <= Logical_Operator_out1047_out1 XOR Logical_Operator_out1079_out1;

  Logical_Operator_out1576_out1 <= Logical_Operator_out1048_out1 XOR Logical_Operator_out1080_out1;

  Logical_Operator_out1577_out1 <= Logical_Operator_out1049_out1 XOR Logical_Operator_out1081_out1;

  Logical_Operator_out1578_out1 <= Logical_Operator_out1050_out1 XOR Logical_Operator_out1082_out1;

  Logical_Operator_out1579_out1 <= Logical_Operator_out1051_out1 XOR Logical_Operator_out1083_out1;

  Logical_Operator_out1580_out1 <= Logical_Operator_out1052_out1 XOR Logical_Operator_out1084_out1;

  Logical_Operator_out1581_out1 <= Logical_Operator_out1053_out1 XOR Logical_Operator_out1085_out1;

  Logical_Operator_out1582_out1 <= Logical_Operator_out1054_out1 XOR Logical_Operator_out1086_out1;

  Logical_Operator_out1583_out1 <= Logical_Operator_out1055_out1 XOR Logical_Operator_out1087_out1;

  Logical_Operator_out1584_out1 <= Logical_Operator_out1056_out1 XOR Logical_Operator_out1088_out1;

  Logical_Operator_out1585_out1 <= Logical_Operator_out793_out1 XOR Logical_Operator_out825_out1;

  Logical_Operator_out1586_out1 <= Logical_Operator_out794_out1 XOR Logical_Operator_out826_out1;

  Logical_Operator_out1587_out1 <= Logical_Operator_out795_out1 XOR Logical_Operator_out827_out1;

  Logical_Operator_out1588_out1 <= Logical_Operator_out796_out1 XOR Logical_Operator_out828_out1;

  Logical_Operator_out1589_out1 <= Logical_Operator_out797_out1 XOR Logical_Operator_out829_out1;

  Logical_Operator_out1590_out1 <= Logical_Operator_out798_out1 XOR Logical_Operator_out830_out1;

  Logical_Operator_out1591_out1 <= Logical_Operator_out799_out1 XOR Logical_Operator_out831_out1;

  Logical_Operator_out1592_out1 <= Logical_Operator_out800_out1 XOR Logical_Operator_out832_out1;

  Logical_Operator_out1593_out1 <= Logical_Operator_out541_out1 XOR Logical_Operator_out573_out1;

  Logical_Operator_out1594_out1 <= Logical_Operator_out542_out1 XOR Logical_Operator_out574_out1;

  Logical_Operator_out1595_out1 <= Logical_Operator_out543_out1 XOR Logical_Operator_out575_out1;

  Logical_Operator_out1596_out1 <= Logical_Operator_out544_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out1597_out1 <= Logical_Operator_out287_out1 XOR Logical_Operator_out319_out1;

  Logical_Operator_out1598_out1 <= Logical_Operator_out288_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out1599_out1 <= Logical_Operator_out32_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out1600_out1 <= in64 XOR in128;

  Logical_Operator_out1601_out1 <= Logical_Operator_out1345_out1 XOR Logical_Operator_out1377_out1;

  Logical_Operator_out1602_out1 <= Logical_Operator_out1346_out1 XOR Logical_Operator_out1378_out1;

  Logical_Operator_out1603_out1 <= Logical_Operator_out1347_out1 XOR Logical_Operator_out1379_out1;

  Logical_Operator_out1604_out1 <= Logical_Operator_out1348_out1 XOR Logical_Operator_out1380_out1;

  Logical_Operator_out1605_out1 <= Logical_Operator_out1349_out1 XOR Logical_Operator_out1381_out1;

  Logical_Operator_out1606_out1 <= Logical_Operator_out1350_out1 XOR Logical_Operator_out1382_out1;

  Logical_Operator_out1607_out1 <= Logical_Operator_out1351_out1 XOR Logical_Operator_out1383_out1;

  Logical_Operator_out1608_out1 <= Logical_Operator_out1352_out1 XOR Logical_Operator_out1384_out1;

  Logical_Operator_out1609_out1 <= Logical_Operator_out1353_out1 XOR Logical_Operator_out1385_out1;

  Logical_Operator_out1610_out1 <= Logical_Operator_out1354_out1 XOR Logical_Operator_out1386_out1;

  Logical_Operator_out1611_out1 <= Logical_Operator_out1355_out1 XOR Logical_Operator_out1387_out1;

  Logical_Operator_out1612_out1 <= Logical_Operator_out1356_out1 XOR Logical_Operator_out1388_out1;

  Logical_Operator_out1613_out1 <= Logical_Operator_out1357_out1 XOR Logical_Operator_out1389_out1;

  Logical_Operator_out1614_out1 <= Logical_Operator_out1358_out1 XOR Logical_Operator_out1390_out1;

  Logical_Operator_out1615_out1 <= Logical_Operator_out1359_out1 XOR Logical_Operator_out1391_out1;

  Logical_Operator_out1616_out1 <= Logical_Operator_out1360_out1 XOR Logical_Operator_out1392_out1;

  Logical_Operator_out1617_out1 <= Logical_Operator_out1361_out1 XOR Logical_Operator_out1393_out1;

  Logical_Operator_out1618_out1 <= Logical_Operator_out1362_out1 XOR Logical_Operator_out1394_out1;

  Logical_Operator_out1619_out1 <= Logical_Operator_out1363_out1 XOR Logical_Operator_out1395_out1;

  Logical_Operator_out1620_out1 <= Logical_Operator_out1364_out1 XOR Logical_Operator_out1396_out1;

  Logical_Operator_out1621_out1 <= Logical_Operator_out1365_out1 XOR Logical_Operator_out1397_out1;

  Logical_Operator_out1622_out1 <= Logical_Operator_out1366_out1 XOR Logical_Operator_out1398_out1;

  Logical_Operator_out1623_out1 <= Logical_Operator_out1367_out1 XOR Logical_Operator_out1399_out1;

  Logical_Operator_out1624_out1 <= Logical_Operator_out1368_out1 XOR Logical_Operator_out1400_out1;

  Logical_Operator_out1625_out1 <= Logical_Operator_out1369_out1 XOR Logical_Operator_out1401_out1;

  Logical_Operator_out1626_out1 <= Logical_Operator_out1370_out1 XOR Logical_Operator_out1402_out1;

  Logical_Operator_out1627_out1 <= Logical_Operator_out1371_out1 XOR Logical_Operator_out1403_out1;

  Logical_Operator_out1628_out1 <= Logical_Operator_out1372_out1 XOR Logical_Operator_out1404_out1;

  Logical_Operator_out1629_out1 <= Logical_Operator_out1373_out1 XOR Logical_Operator_out1405_out1;

  Logical_Operator_out1630_out1 <= Logical_Operator_out1374_out1 XOR Logical_Operator_out1406_out1;

  Logical_Operator_out1631_out1 <= Logical_Operator_out1375_out1 XOR Logical_Operator_out1407_out1;

  Logical_Operator_out1632_out1 <= Logical_Operator_out1376_out1 XOR Logical_Operator_out1408_out1;

  Logical_Operator_out1633_out1 <= Logical_Operator_out1105_out1 XOR Logical_Operator_out1137_out1;

  Logical_Operator_out1634_out1 <= Logical_Operator_out1106_out1 XOR Logical_Operator_out1138_out1;

  Logical_Operator_out1635_out1 <= Logical_Operator_out1107_out1 XOR Logical_Operator_out1139_out1;

  Logical_Operator_out1636_out1 <= Logical_Operator_out1108_out1 XOR Logical_Operator_out1140_out1;

  Logical_Operator_out1637_out1 <= Logical_Operator_out1109_out1 XOR Logical_Operator_out1141_out1;

  Logical_Operator_out1638_out1 <= Logical_Operator_out1110_out1 XOR Logical_Operator_out1142_out1;

  Logical_Operator_out1639_out1 <= Logical_Operator_out1111_out1 XOR Logical_Operator_out1143_out1;

  Logical_Operator_out1640_out1 <= Logical_Operator_out1112_out1 XOR Logical_Operator_out1144_out1;

  Logical_Operator_out1641_out1 <= Logical_Operator_out1113_out1 XOR Logical_Operator_out1145_out1;

  Logical_Operator_out1642_out1 <= Logical_Operator_out1114_out1 XOR Logical_Operator_out1146_out1;

  Logical_Operator_out1643_out1 <= Logical_Operator_out1115_out1 XOR Logical_Operator_out1147_out1;

  Logical_Operator_out1644_out1 <= Logical_Operator_out1116_out1 XOR Logical_Operator_out1148_out1;

  Logical_Operator_out1645_out1 <= Logical_Operator_out1117_out1 XOR Logical_Operator_out1149_out1;

  Logical_Operator_out1646_out1 <= Logical_Operator_out1118_out1 XOR Logical_Operator_out1150_out1;

  Logical_Operator_out1647_out1 <= Logical_Operator_out1119_out1 XOR Logical_Operator_out1151_out1;

  Logical_Operator_out1648_out1 <= Logical_Operator_out1120_out1 XOR Logical_Operator_out1152_out1;

  Logical_Operator_out1649_out1 <= Logical_Operator_out857_out1 XOR Logical_Operator_out889_out1;

  Logical_Operator_out1650_out1 <= Logical_Operator_out858_out1 XOR Logical_Operator_out890_out1;

  Logical_Operator_out1651_out1 <= Logical_Operator_out859_out1 XOR Logical_Operator_out891_out1;

  Logical_Operator_out1652_out1 <= Logical_Operator_out860_out1 XOR Logical_Operator_out892_out1;

  Logical_Operator_out1653_out1 <= Logical_Operator_out861_out1 XOR Logical_Operator_out893_out1;

  Logical_Operator_out1654_out1 <= Logical_Operator_out862_out1 XOR Logical_Operator_out894_out1;

  Logical_Operator_out1655_out1 <= Logical_Operator_out863_out1 XOR Logical_Operator_out895_out1;

  Logical_Operator_out1656_out1 <= Logical_Operator_out864_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out1657_out1 <= Logical_Operator_out605_out1 XOR Logical_Operator_out637_out1;

  Logical_Operator_out1658_out1 <= Logical_Operator_out606_out1 XOR Logical_Operator_out638_out1;

  Logical_Operator_out1659_out1 <= Logical_Operator_out607_out1 XOR Logical_Operator_out639_out1;

  Logical_Operator_out1660_out1 <= Logical_Operator_out608_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out1661_out1 <= Logical_Operator_out351_out1 XOR Logical_Operator_out383_out1;

  Logical_Operator_out1662_out1 <= Logical_Operator_out352_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out1663_out1 <= Logical_Operator_out96_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out1664_out1 <= in192 XOR in256;

  Logical_Operator_out1665_out1 <= Logical_Operator_out1409_out1 XOR Logical_Operator_out1441_out1;

  Logical_Operator_out1666_out1 <= Logical_Operator_out1410_out1 XOR Logical_Operator_out1442_out1;

  Logical_Operator_out1667_out1 <= Logical_Operator_out1411_out1 XOR Logical_Operator_out1443_out1;

  Logical_Operator_out1668_out1 <= Logical_Operator_out1412_out1 XOR Logical_Operator_out1444_out1;

  Logical_Operator_out1669_out1 <= Logical_Operator_out1413_out1 XOR Logical_Operator_out1445_out1;

  Logical_Operator_out1670_out1 <= Logical_Operator_out1414_out1 XOR Logical_Operator_out1446_out1;

  Logical_Operator_out1671_out1 <= Logical_Operator_out1415_out1 XOR Logical_Operator_out1447_out1;

  Logical_Operator_out1672_out1 <= Logical_Operator_out1416_out1 XOR Logical_Operator_out1448_out1;

  Logical_Operator_out1673_out1 <= Logical_Operator_out1417_out1 XOR Logical_Operator_out1449_out1;

  Logical_Operator_out1674_out1 <= Logical_Operator_out1418_out1 XOR Logical_Operator_out1450_out1;

  Logical_Operator_out1675_out1 <= Logical_Operator_out1419_out1 XOR Logical_Operator_out1451_out1;

  Logical_Operator_out1676_out1 <= Logical_Operator_out1420_out1 XOR Logical_Operator_out1452_out1;

  Logical_Operator_out1677_out1 <= Logical_Operator_out1421_out1 XOR Logical_Operator_out1453_out1;

  Logical_Operator_out1678_out1 <= Logical_Operator_out1422_out1 XOR Logical_Operator_out1454_out1;

  Logical_Operator_out1679_out1 <= Logical_Operator_out1423_out1 XOR Logical_Operator_out1455_out1;

  Logical_Operator_out1680_out1 <= Logical_Operator_out1424_out1 XOR Logical_Operator_out1456_out1;

  Logical_Operator_out1681_out1 <= Logical_Operator_out1425_out1 XOR Logical_Operator_out1457_out1;

  Logical_Operator_out1682_out1 <= Logical_Operator_out1426_out1 XOR Logical_Operator_out1458_out1;

  Logical_Operator_out1683_out1 <= Logical_Operator_out1427_out1 XOR Logical_Operator_out1459_out1;

  Logical_Operator_out1684_out1 <= Logical_Operator_out1428_out1 XOR Logical_Operator_out1460_out1;

  Logical_Operator_out1685_out1 <= Logical_Operator_out1429_out1 XOR Logical_Operator_out1461_out1;

  Logical_Operator_out1686_out1 <= Logical_Operator_out1430_out1 XOR Logical_Operator_out1462_out1;

  Logical_Operator_out1687_out1 <= Logical_Operator_out1431_out1 XOR Logical_Operator_out1463_out1;

  Logical_Operator_out1688_out1 <= Logical_Operator_out1432_out1 XOR Logical_Operator_out1464_out1;

  Logical_Operator_out1689_out1 <= Logical_Operator_out1433_out1 XOR Logical_Operator_out1465_out1;

  Logical_Operator_out1690_out1 <= Logical_Operator_out1434_out1 XOR Logical_Operator_out1466_out1;

  Logical_Operator_out1691_out1 <= Logical_Operator_out1435_out1 XOR Logical_Operator_out1467_out1;

  Logical_Operator_out1692_out1 <= Logical_Operator_out1436_out1 XOR Logical_Operator_out1468_out1;

  Logical_Operator_out1693_out1 <= Logical_Operator_out1437_out1 XOR Logical_Operator_out1469_out1;

  Logical_Operator_out1694_out1 <= Logical_Operator_out1438_out1 XOR Logical_Operator_out1470_out1;

  Logical_Operator_out1695_out1 <= Logical_Operator_out1439_out1 XOR Logical_Operator_out1471_out1;

  Logical_Operator_out1696_out1 <= Logical_Operator_out1440_out1 XOR Logical_Operator_out1472_out1;

  Logical_Operator_out1697_out1 <= Logical_Operator_out1169_out1 XOR Logical_Operator_out1201_out1;

  Logical_Operator_out1698_out1 <= Logical_Operator_out1170_out1 XOR Logical_Operator_out1202_out1;

  Logical_Operator_out1699_out1 <= Logical_Operator_out1171_out1 XOR Logical_Operator_out1203_out1;

  Logical_Operator_out1700_out1 <= Logical_Operator_out1172_out1 XOR Logical_Operator_out1204_out1;

  Logical_Operator_out1701_out1 <= Logical_Operator_out1173_out1 XOR Logical_Operator_out1205_out1;

  Logical_Operator_out1702_out1 <= Logical_Operator_out1174_out1 XOR Logical_Operator_out1206_out1;

  Logical_Operator_out1703_out1 <= Logical_Operator_out1175_out1 XOR Logical_Operator_out1207_out1;

  Logical_Operator_out1704_out1 <= Logical_Operator_out1176_out1 XOR Logical_Operator_out1208_out1;

  Logical_Operator_out1705_out1 <= Logical_Operator_out1177_out1 XOR Logical_Operator_out1209_out1;

  Logical_Operator_out1706_out1 <= Logical_Operator_out1178_out1 XOR Logical_Operator_out1210_out1;

  Logical_Operator_out1707_out1 <= Logical_Operator_out1179_out1 XOR Logical_Operator_out1211_out1;

  Logical_Operator_out1708_out1 <= Logical_Operator_out1180_out1 XOR Logical_Operator_out1212_out1;

  Logical_Operator_out1709_out1 <= Logical_Operator_out1181_out1 XOR Logical_Operator_out1213_out1;

  Logical_Operator_out1710_out1 <= Logical_Operator_out1182_out1 XOR Logical_Operator_out1214_out1;

  Logical_Operator_out1711_out1 <= Logical_Operator_out1183_out1 XOR Logical_Operator_out1215_out1;

  Logical_Operator_out1712_out1 <= Logical_Operator_out1184_out1 XOR Logical_Operator_out1216_out1;

  Logical_Operator_out1713_out1 <= Logical_Operator_out921_out1 XOR Logical_Operator_out953_out1;

  Logical_Operator_out1714_out1 <= Logical_Operator_out922_out1 XOR Logical_Operator_out954_out1;

  Logical_Operator_out1715_out1 <= Logical_Operator_out923_out1 XOR Logical_Operator_out955_out1;

  Logical_Operator_out1716_out1 <= Logical_Operator_out924_out1 XOR Logical_Operator_out956_out1;

  Logical_Operator_out1717_out1 <= Logical_Operator_out925_out1 XOR Logical_Operator_out957_out1;

  Logical_Operator_out1718_out1 <= Logical_Operator_out926_out1 XOR Logical_Operator_out958_out1;

  Logical_Operator_out1719_out1 <= Logical_Operator_out927_out1 XOR Logical_Operator_out959_out1;

  Logical_Operator_out1720_out1 <= Logical_Operator_out928_out1 XOR Logical_Operator_out960_out1;

  Logical_Operator_out1721_out1 <= Logical_Operator_out669_out1 XOR Logical_Operator_out701_out1;

  Logical_Operator_out1722_out1 <= Logical_Operator_out670_out1 XOR Logical_Operator_out702_out1;

  Logical_Operator_out1723_out1 <= Logical_Operator_out671_out1 XOR Logical_Operator_out703_out1;

  Logical_Operator_out1724_out1 <= Logical_Operator_out672_out1 XOR Logical_Operator_out704_out1;

  Logical_Operator_out1725_out1 <= Logical_Operator_out415_out1 XOR Logical_Operator_out447_out1;

  Logical_Operator_out1726_out1 <= Logical_Operator_out416_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out1727_out1 <= Logical_Operator_out160_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out1728_out1 <= in320 XOR in384;

  Logical_Operator_out1729_out1 <= Logical_Operator_out1473_out1 XOR Logical_Operator_out1505_out1;

  Logical_Operator_out1730_out1 <= Logical_Operator_out1474_out1 XOR Logical_Operator_out1506_out1;

  Logical_Operator_out1731_out1 <= Logical_Operator_out1475_out1 XOR Logical_Operator_out1507_out1;

  Logical_Operator_out1732_out1 <= Logical_Operator_out1476_out1 XOR Logical_Operator_out1508_out1;

  Logical_Operator_out1733_out1 <= Logical_Operator_out1477_out1 XOR Logical_Operator_out1509_out1;

  Logical_Operator_out1734_out1 <= Logical_Operator_out1478_out1 XOR Logical_Operator_out1510_out1;

  Logical_Operator_out1735_out1 <= Logical_Operator_out1479_out1 XOR Logical_Operator_out1511_out1;

  Logical_Operator_out1736_out1 <= Logical_Operator_out1480_out1 XOR Logical_Operator_out1512_out1;

  Logical_Operator_out1737_out1 <= Logical_Operator_out1481_out1 XOR Logical_Operator_out1513_out1;

  Logical_Operator_out1738_out1 <= Logical_Operator_out1482_out1 XOR Logical_Operator_out1514_out1;

  Logical_Operator_out1739_out1 <= Logical_Operator_out1483_out1 XOR Logical_Operator_out1515_out1;

  Logical_Operator_out1740_out1 <= Logical_Operator_out1484_out1 XOR Logical_Operator_out1516_out1;

  Logical_Operator_out1741_out1 <= Logical_Operator_out1485_out1 XOR Logical_Operator_out1517_out1;

  Logical_Operator_out1742_out1 <= Logical_Operator_out1486_out1 XOR Logical_Operator_out1518_out1;

  Logical_Operator_out1743_out1 <= Logical_Operator_out1487_out1 XOR Logical_Operator_out1519_out1;

  Logical_Operator_out1744_out1 <= Logical_Operator_out1488_out1 XOR Logical_Operator_out1520_out1;

  Logical_Operator_out1745_out1 <= Logical_Operator_out1489_out1 XOR Logical_Operator_out1521_out1;

  Logical_Operator_out1746_out1 <= Logical_Operator_out1490_out1 XOR Logical_Operator_out1522_out1;

  Logical_Operator_out1747_out1 <= Logical_Operator_out1491_out1 XOR Logical_Operator_out1523_out1;

  Logical_Operator_out1748_out1 <= Logical_Operator_out1492_out1 XOR Logical_Operator_out1524_out1;

  Logical_Operator_out1749_out1 <= Logical_Operator_out1493_out1 XOR Logical_Operator_out1525_out1;

  Logical_Operator_out1750_out1 <= Logical_Operator_out1494_out1 XOR Logical_Operator_out1526_out1;

  Logical_Operator_out1751_out1 <= Logical_Operator_out1495_out1 XOR Logical_Operator_out1527_out1;

  Logical_Operator_out1752_out1 <= Logical_Operator_out1496_out1 XOR Logical_Operator_out1528_out1;

  Logical_Operator_out1753_out1 <= Logical_Operator_out1497_out1 XOR Logical_Operator_out1529_out1;

  Logical_Operator_out1754_out1 <= Logical_Operator_out1498_out1 XOR Logical_Operator_out1530_out1;

  Logical_Operator_out1755_out1 <= Logical_Operator_out1499_out1 XOR Logical_Operator_out1531_out1;

  Logical_Operator_out1756_out1 <= Logical_Operator_out1500_out1 XOR Logical_Operator_out1532_out1;

  Logical_Operator_out1757_out1 <= Logical_Operator_out1501_out1 XOR Logical_Operator_out1533_out1;

  Logical_Operator_out1758_out1 <= Logical_Operator_out1502_out1 XOR Logical_Operator_out1534_out1;

  Logical_Operator_out1759_out1 <= Logical_Operator_out1503_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out1760_out1 <= Logical_Operator_out1504_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out1761_out1 <= Logical_Operator_out1233_out1 XOR Logical_Operator_out1265_out1;

  Logical_Operator_out1762_out1 <= Logical_Operator_out1234_out1 XOR Logical_Operator_out1266_out1;

  Logical_Operator_out1763_out1 <= Logical_Operator_out1235_out1 XOR Logical_Operator_out1267_out1;

  Logical_Operator_out1764_out1 <= Logical_Operator_out1236_out1 XOR Logical_Operator_out1268_out1;

  Logical_Operator_out1765_out1 <= Logical_Operator_out1237_out1 XOR Logical_Operator_out1269_out1;

  Logical_Operator_out1766_out1 <= Logical_Operator_out1238_out1 XOR Logical_Operator_out1270_out1;

  Logical_Operator_out1767_out1 <= Logical_Operator_out1239_out1 XOR Logical_Operator_out1271_out1;

  Logical_Operator_out1768_out1 <= Logical_Operator_out1240_out1 XOR Logical_Operator_out1272_out1;

  Logical_Operator_out1769_out1 <= Logical_Operator_out1241_out1 XOR Logical_Operator_out1273_out1;

  Logical_Operator_out1770_out1 <= Logical_Operator_out1242_out1 XOR Logical_Operator_out1274_out1;

  Logical_Operator_out1771_out1 <= Logical_Operator_out1243_out1 XOR Logical_Operator_out1275_out1;

  Logical_Operator_out1772_out1 <= Logical_Operator_out1244_out1 XOR Logical_Operator_out1276_out1;

  Logical_Operator_out1773_out1 <= Logical_Operator_out1245_out1 XOR Logical_Operator_out1277_out1;

  Logical_Operator_out1774_out1 <= Logical_Operator_out1246_out1 XOR Logical_Operator_out1278_out1;

  Logical_Operator_out1775_out1 <= Logical_Operator_out1247_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out1776_out1 <= Logical_Operator_out1248_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out1777_out1 <= Logical_Operator_out985_out1 XOR Logical_Operator_out1017_out1;

  Logical_Operator_out1778_out1 <= Logical_Operator_out986_out1 XOR Logical_Operator_out1018_out1;

  Logical_Operator_out1779_out1 <= Logical_Operator_out987_out1 XOR Logical_Operator_out1019_out1;

  Logical_Operator_out1780_out1 <= Logical_Operator_out988_out1 XOR Logical_Operator_out1020_out1;

  Logical_Operator_out1781_out1 <= Logical_Operator_out989_out1 XOR Logical_Operator_out1021_out1;

  Logical_Operator_out1782_out1 <= Logical_Operator_out990_out1 XOR Logical_Operator_out1022_out1;

  Logical_Operator_out1783_out1 <= Logical_Operator_out991_out1 XOR Logical_Operator_out1023_out1;

  Logical_Operator_out1784_out1 <= Logical_Operator_out992_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out1785_out1 <= Logical_Operator_out733_out1 XOR Logical_Operator_out765_out1;

  Logical_Operator_out1786_out1 <= Logical_Operator_out734_out1 XOR Logical_Operator_out766_out1;

  Logical_Operator_out1787_out1 <= Logical_Operator_out735_out1 XOR Logical_Operator_out767_out1;

  Logical_Operator_out1788_out1 <= Logical_Operator_out736_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out1789_out1 <= Logical_Operator_out479_out1 XOR Logical_Operator_out511_out1;

  Logical_Operator_out1790_out1 <= Logical_Operator_out480_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out1791_out1 <= Logical_Operator_out224_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out1792_out1 <= in448 XOR in512;

  Logical_Operator_out1793_out1 <= Logical_Operator_out1537_out1 XOR Logical_Operator_out1601_out1;

  Logical_Operator_out1794_out1 <= Logical_Operator_out1538_out1 XOR Logical_Operator_out1602_out1;

  Logical_Operator_out1795_out1 <= Logical_Operator_out1539_out1 XOR Logical_Operator_out1603_out1;

  Logical_Operator_out1796_out1 <= Logical_Operator_out1540_out1 XOR Logical_Operator_out1604_out1;

  Logical_Operator_out1797_out1 <= Logical_Operator_out1541_out1 XOR Logical_Operator_out1605_out1;

  Logical_Operator_out1798_out1 <= Logical_Operator_out1542_out1 XOR Logical_Operator_out1606_out1;

  Logical_Operator_out1799_out1 <= Logical_Operator_out1543_out1 XOR Logical_Operator_out1607_out1;

  Logical_Operator_out1800_out1 <= Logical_Operator_out1544_out1 XOR Logical_Operator_out1608_out1;

  Logical_Operator_out1801_out1 <= Logical_Operator_out1545_out1 XOR Logical_Operator_out1609_out1;

  Logical_Operator_out1802_out1 <= Logical_Operator_out1546_out1 XOR Logical_Operator_out1610_out1;

  Logical_Operator_out1803_out1 <= Logical_Operator_out1547_out1 XOR Logical_Operator_out1611_out1;

  Logical_Operator_out1804_out1 <= Logical_Operator_out1548_out1 XOR Logical_Operator_out1612_out1;

  Logical_Operator_out1805_out1 <= Logical_Operator_out1549_out1 XOR Logical_Operator_out1613_out1;

  Logical_Operator_out1806_out1 <= Logical_Operator_out1550_out1 XOR Logical_Operator_out1614_out1;

  Logical_Operator_out1807_out1 <= Logical_Operator_out1551_out1 XOR Logical_Operator_out1615_out1;

  Logical_Operator_out1808_out1 <= Logical_Operator_out1552_out1 XOR Logical_Operator_out1616_out1;

  Logical_Operator_out1809_out1 <= Logical_Operator_out1553_out1 XOR Logical_Operator_out1617_out1;

  Logical_Operator_out1810_out1 <= Logical_Operator_out1554_out1 XOR Logical_Operator_out1618_out1;

  Logical_Operator_out1811_out1 <= Logical_Operator_out1555_out1 XOR Logical_Operator_out1619_out1;

  Logical_Operator_out1812_out1 <= Logical_Operator_out1556_out1 XOR Logical_Operator_out1620_out1;

  Logical_Operator_out1813_out1 <= Logical_Operator_out1557_out1 XOR Logical_Operator_out1621_out1;

  Logical_Operator_out1814_out1 <= Logical_Operator_out1558_out1 XOR Logical_Operator_out1622_out1;

  Logical_Operator_out1815_out1 <= Logical_Operator_out1559_out1 XOR Logical_Operator_out1623_out1;

  Logical_Operator_out1816_out1 <= Logical_Operator_out1560_out1 XOR Logical_Operator_out1624_out1;

  Logical_Operator_out1817_out1 <= Logical_Operator_out1561_out1 XOR Logical_Operator_out1625_out1;

  Logical_Operator_out1818_out1 <= Logical_Operator_out1562_out1 XOR Logical_Operator_out1626_out1;

  Logical_Operator_out1819_out1 <= Logical_Operator_out1563_out1 XOR Logical_Operator_out1627_out1;

  Logical_Operator_out1820_out1 <= Logical_Operator_out1564_out1 XOR Logical_Operator_out1628_out1;

  Logical_Operator_out1821_out1 <= Logical_Operator_out1565_out1 XOR Logical_Operator_out1629_out1;

  Logical_Operator_out1822_out1 <= Logical_Operator_out1566_out1 XOR Logical_Operator_out1630_out1;

  Logical_Operator_out1823_out1 <= Logical_Operator_out1567_out1 XOR Logical_Operator_out1631_out1;

  Logical_Operator_out1824_out1 <= Logical_Operator_out1568_out1 XOR Logical_Operator_out1632_out1;

  Logical_Operator_out1825_out1 <= Logical_Operator_out1569_out1 XOR Logical_Operator_out1633_out1;

  Logical_Operator_out1826_out1 <= Logical_Operator_out1570_out1 XOR Logical_Operator_out1634_out1;

  Logical_Operator_out1827_out1 <= Logical_Operator_out1571_out1 XOR Logical_Operator_out1635_out1;

  Logical_Operator_out1828_out1 <= Logical_Operator_out1572_out1 XOR Logical_Operator_out1636_out1;

  Logical_Operator_out1829_out1 <= Logical_Operator_out1573_out1 XOR Logical_Operator_out1637_out1;

  Logical_Operator_out1830_out1 <= Logical_Operator_out1574_out1 XOR Logical_Operator_out1638_out1;

  Logical_Operator_out1831_out1 <= Logical_Operator_out1575_out1 XOR Logical_Operator_out1639_out1;

  Logical_Operator_out1832_out1 <= Logical_Operator_out1576_out1 XOR Logical_Operator_out1640_out1;

  Logical_Operator_out1833_out1 <= Logical_Operator_out1577_out1 XOR Logical_Operator_out1641_out1;

  Logical_Operator_out1834_out1 <= Logical_Operator_out1578_out1 XOR Logical_Operator_out1642_out1;

  Logical_Operator_out1835_out1 <= Logical_Operator_out1579_out1 XOR Logical_Operator_out1643_out1;

  Logical_Operator_out1836_out1 <= Logical_Operator_out1580_out1 XOR Logical_Operator_out1644_out1;

  Logical_Operator_out1837_out1 <= Logical_Operator_out1581_out1 XOR Logical_Operator_out1645_out1;

  Logical_Operator_out1838_out1 <= Logical_Operator_out1582_out1 XOR Logical_Operator_out1646_out1;

  Logical_Operator_out1839_out1 <= Logical_Operator_out1583_out1 XOR Logical_Operator_out1647_out1;

  Logical_Operator_out1840_out1 <= Logical_Operator_out1584_out1 XOR Logical_Operator_out1648_out1;

  Logical_Operator_out1841_out1 <= Logical_Operator_out1585_out1 XOR Logical_Operator_out1649_out1;

  Logical_Operator_out1842_out1 <= Logical_Operator_out1586_out1 XOR Logical_Operator_out1650_out1;

  Logical_Operator_out1843_out1 <= Logical_Operator_out1587_out1 XOR Logical_Operator_out1651_out1;

  Logical_Operator_out1844_out1 <= Logical_Operator_out1588_out1 XOR Logical_Operator_out1652_out1;

  Logical_Operator_out1845_out1 <= Logical_Operator_out1589_out1 XOR Logical_Operator_out1653_out1;

  Logical_Operator_out1846_out1 <= Logical_Operator_out1590_out1 XOR Logical_Operator_out1654_out1;

  Logical_Operator_out1847_out1 <= Logical_Operator_out1591_out1 XOR Logical_Operator_out1655_out1;

  Logical_Operator_out1848_out1 <= Logical_Operator_out1592_out1 XOR Logical_Operator_out1656_out1;

  Logical_Operator_out1849_out1 <= Logical_Operator_out1593_out1 XOR Logical_Operator_out1657_out1;

  Logical_Operator_out1850_out1 <= Logical_Operator_out1594_out1 XOR Logical_Operator_out1658_out1;

  Logical_Operator_out1851_out1 <= Logical_Operator_out1595_out1 XOR Logical_Operator_out1659_out1;

  Logical_Operator_out1852_out1 <= Logical_Operator_out1596_out1 XOR Logical_Operator_out1660_out1;

  Logical_Operator_out1853_out1 <= Logical_Operator_out1597_out1 XOR Logical_Operator_out1661_out1;

  Logical_Operator_out1854_out1 <= Logical_Operator_out1598_out1 XOR Logical_Operator_out1662_out1;

  Logical_Operator_out1855_out1 <= Logical_Operator_out1599_out1 XOR Logical_Operator_out1663_out1;

  Logical_Operator_out1856_out1 <= Logical_Operator_out1600_out1 XOR Logical_Operator_out1664_out1;

  Logical_Operator_out1857_out1 <= Logical_Operator_out1313_out1 XOR Logical_Operator_out1377_out1;

  Logical_Operator_out1858_out1 <= Logical_Operator_out1314_out1 XOR Logical_Operator_out1378_out1;

  Logical_Operator_out1859_out1 <= Logical_Operator_out1315_out1 XOR Logical_Operator_out1379_out1;

  Logical_Operator_out1860_out1 <= Logical_Operator_out1316_out1 XOR Logical_Operator_out1380_out1;

  Logical_Operator_out1861_out1 <= Logical_Operator_out1317_out1 XOR Logical_Operator_out1381_out1;

  Logical_Operator_out1862_out1 <= Logical_Operator_out1318_out1 XOR Logical_Operator_out1382_out1;

  Logical_Operator_out1863_out1 <= Logical_Operator_out1319_out1 XOR Logical_Operator_out1383_out1;

  Logical_Operator_out1864_out1 <= Logical_Operator_out1320_out1 XOR Logical_Operator_out1384_out1;

  Logical_Operator_out1865_out1 <= Logical_Operator_out1321_out1 XOR Logical_Operator_out1385_out1;

  Logical_Operator_out1866_out1 <= Logical_Operator_out1322_out1 XOR Logical_Operator_out1386_out1;

  Logical_Operator_out1867_out1 <= Logical_Operator_out1323_out1 XOR Logical_Operator_out1387_out1;

  Logical_Operator_out1868_out1 <= Logical_Operator_out1324_out1 XOR Logical_Operator_out1388_out1;

  Logical_Operator_out1869_out1 <= Logical_Operator_out1325_out1 XOR Logical_Operator_out1389_out1;

  Logical_Operator_out1870_out1 <= Logical_Operator_out1326_out1 XOR Logical_Operator_out1390_out1;

  Logical_Operator_out1871_out1 <= Logical_Operator_out1327_out1 XOR Logical_Operator_out1391_out1;

  Logical_Operator_out1872_out1 <= Logical_Operator_out1328_out1 XOR Logical_Operator_out1392_out1;

  Logical_Operator_out1873_out1 <= Logical_Operator_out1329_out1 XOR Logical_Operator_out1393_out1;

  Logical_Operator_out1874_out1 <= Logical_Operator_out1330_out1 XOR Logical_Operator_out1394_out1;

  Logical_Operator_out1875_out1 <= Logical_Operator_out1331_out1 XOR Logical_Operator_out1395_out1;

  Logical_Operator_out1876_out1 <= Logical_Operator_out1332_out1 XOR Logical_Operator_out1396_out1;

  Logical_Operator_out1877_out1 <= Logical_Operator_out1333_out1 XOR Logical_Operator_out1397_out1;

  Logical_Operator_out1878_out1 <= Logical_Operator_out1334_out1 XOR Logical_Operator_out1398_out1;

  Logical_Operator_out1879_out1 <= Logical_Operator_out1335_out1 XOR Logical_Operator_out1399_out1;

  Logical_Operator_out1880_out1 <= Logical_Operator_out1336_out1 XOR Logical_Operator_out1400_out1;

  Logical_Operator_out1881_out1 <= Logical_Operator_out1337_out1 XOR Logical_Operator_out1401_out1;

  Logical_Operator_out1882_out1 <= Logical_Operator_out1338_out1 XOR Logical_Operator_out1402_out1;

  Logical_Operator_out1883_out1 <= Logical_Operator_out1339_out1 XOR Logical_Operator_out1403_out1;

  Logical_Operator_out1884_out1 <= Logical_Operator_out1340_out1 XOR Logical_Operator_out1404_out1;

  Logical_Operator_out1885_out1 <= Logical_Operator_out1341_out1 XOR Logical_Operator_out1405_out1;

  Logical_Operator_out1886_out1 <= Logical_Operator_out1342_out1 XOR Logical_Operator_out1406_out1;

  Logical_Operator_out1887_out1 <= Logical_Operator_out1343_out1 XOR Logical_Operator_out1407_out1;

  Logical_Operator_out1888_out1 <= Logical_Operator_out1344_out1 XOR Logical_Operator_out1408_out1;

  Logical_Operator_out1889_out1 <= Logical_Operator_out1073_out1 XOR Logical_Operator_out1137_out1;

  Logical_Operator_out1890_out1 <= Logical_Operator_out1074_out1 XOR Logical_Operator_out1138_out1;

  Logical_Operator_out1891_out1 <= Logical_Operator_out1075_out1 XOR Logical_Operator_out1139_out1;

  Logical_Operator_out1892_out1 <= Logical_Operator_out1076_out1 XOR Logical_Operator_out1140_out1;

  Logical_Operator_out1893_out1 <= Logical_Operator_out1077_out1 XOR Logical_Operator_out1141_out1;

  Logical_Operator_out1894_out1 <= Logical_Operator_out1078_out1 XOR Logical_Operator_out1142_out1;

  Logical_Operator_out1895_out1 <= Logical_Operator_out1079_out1 XOR Logical_Operator_out1143_out1;

  Logical_Operator_out1896_out1 <= Logical_Operator_out1080_out1 XOR Logical_Operator_out1144_out1;

  Logical_Operator_out1897_out1 <= Logical_Operator_out1081_out1 XOR Logical_Operator_out1145_out1;

  Logical_Operator_out1898_out1 <= Logical_Operator_out1082_out1 XOR Logical_Operator_out1146_out1;

  Logical_Operator_out1899_out1 <= Logical_Operator_out1083_out1 XOR Logical_Operator_out1147_out1;

  Logical_Operator_out1900_out1 <= Logical_Operator_out1084_out1 XOR Logical_Operator_out1148_out1;

  Logical_Operator_out1901_out1 <= Logical_Operator_out1085_out1 XOR Logical_Operator_out1149_out1;

  Logical_Operator_out1902_out1 <= Logical_Operator_out1086_out1 XOR Logical_Operator_out1150_out1;

  Logical_Operator_out1903_out1 <= Logical_Operator_out1087_out1 XOR Logical_Operator_out1151_out1;

  Logical_Operator_out1904_out1 <= Logical_Operator_out1088_out1 XOR Logical_Operator_out1152_out1;

  Logical_Operator_out1905_out1 <= Logical_Operator_out825_out1 XOR Logical_Operator_out889_out1;

  Logical_Operator_out1906_out1 <= Logical_Operator_out826_out1 XOR Logical_Operator_out890_out1;

  Logical_Operator_out1907_out1 <= Logical_Operator_out827_out1 XOR Logical_Operator_out891_out1;

  Logical_Operator_out1908_out1 <= Logical_Operator_out828_out1 XOR Logical_Operator_out892_out1;

  Logical_Operator_out1909_out1 <= Logical_Operator_out829_out1 XOR Logical_Operator_out893_out1;

  Logical_Operator_out1910_out1 <= Logical_Operator_out830_out1 XOR Logical_Operator_out894_out1;

  Logical_Operator_out1911_out1 <= Logical_Operator_out831_out1 XOR Logical_Operator_out895_out1;

  Logical_Operator_out1912_out1 <= Logical_Operator_out832_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out1913_out1 <= Logical_Operator_out573_out1 XOR Logical_Operator_out637_out1;

  Logical_Operator_out1914_out1 <= Logical_Operator_out574_out1 XOR Logical_Operator_out638_out1;

  Logical_Operator_out1915_out1 <= Logical_Operator_out575_out1 XOR Logical_Operator_out639_out1;

  Logical_Operator_out1916_out1 <= Logical_Operator_out576_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out1917_out1 <= Logical_Operator_out319_out1 XOR Logical_Operator_out383_out1;

  Logical_Operator_out1918_out1 <= Logical_Operator_out320_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out1919_out1 <= Logical_Operator_out64_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out1920_out1 <= in128 XOR in256;

  Logical_Operator_out1921_out1 <= Logical_Operator_out1665_out1 XOR Logical_Operator_out1729_out1;

  Logical_Operator_out1922_out1 <= Logical_Operator_out1666_out1 XOR Logical_Operator_out1730_out1;

  Logical_Operator_out1923_out1 <= Logical_Operator_out1667_out1 XOR Logical_Operator_out1731_out1;

  Logical_Operator_out1924_out1 <= Logical_Operator_out1668_out1 XOR Logical_Operator_out1732_out1;

  Logical_Operator_out1925_out1 <= Logical_Operator_out1669_out1 XOR Logical_Operator_out1733_out1;

  Logical_Operator_out1926_out1 <= Logical_Operator_out1670_out1 XOR Logical_Operator_out1734_out1;

  Logical_Operator_out1927_out1 <= Logical_Operator_out1671_out1 XOR Logical_Operator_out1735_out1;

  Logical_Operator_out1928_out1 <= Logical_Operator_out1672_out1 XOR Logical_Operator_out1736_out1;

  Logical_Operator_out1929_out1 <= Logical_Operator_out1673_out1 XOR Logical_Operator_out1737_out1;

  Logical_Operator_out1930_out1 <= Logical_Operator_out1674_out1 XOR Logical_Operator_out1738_out1;

  Logical_Operator_out1931_out1 <= Logical_Operator_out1675_out1 XOR Logical_Operator_out1739_out1;

  Logical_Operator_out1932_out1 <= Logical_Operator_out1676_out1 XOR Logical_Operator_out1740_out1;

  Logical_Operator_out1933_out1 <= Logical_Operator_out1677_out1 XOR Logical_Operator_out1741_out1;

  Logical_Operator_out1934_out1 <= Logical_Operator_out1678_out1 XOR Logical_Operator_out1742_out1;

  Logical_Operator_out1935_out1 <= Logical_Operator_out1679_out1 XOR Logical_Operator_out1743_out1;

  Logical_Operator_out1936_out1 <= Logical_Operator_out1680_out1 XOR Logical_Operator_out1744_out1;

  Logical_Operator_out1937_out1 <= Logical_Operator_out1681_out1 XOR Logical_Operator_out1745_out1;

  Logical_Operator_out1938_out1 <= Logical_Operator_out1682_out1 XOR Logical_Operator_out1746_out1;

  Logical_Operator_out1939_out1 <= Logical_Operator_out1683_out1 XOR Logical_Operator_out1747_out1;

  Logical_Operator_out1940_out1 <= Logical_Operator_out1684_out1 XOR Logical_Operator_out1748_out1;

  Logical_Operator_out1941_out1 <= Logical_Operator_out1685_out1 XOR Logical_Operator_out1749_out1;

  Logical_Operator_out1942_out1 <= Logical_Operator_out1686_out1 XOR Logical_Operator_out1750_out1;

  Logical_Operator_out1943_out1 <= Logical_Operator_out1687_out1 XOR Logical_Operator_out1751_out1;

  Logical_Operator_out1944_out1 <= Logical_Operator_out1688_out1 XOR Logical_Operator_out1752_out1;

  Logical_Operator_out1945_out1 <= Logical_Operator_out1689_out1 XOR Logical_Operator_out1753_out1;

  Logical_Operator_out1946_out1 <= Logical_Operator_out1690_out1 XOR Logical_Operator_out1754_out1;

  Logical_Operator_out1947_out1 <= Logical_Operator_out1691_out1 XOR Logical_Operator_out1755_out1;

  Logical_Operator_out1948_out1 <= Logical_Operator_out1692_out1 XOR Logical_Operator_out1756_out1;

  Logical_Operator_out1949_out1 <= Logical_Operator_out1693_out1 XOR Logical_Operator_out1757_out1;

  Logical_Operator_out1950_out1 <= Logical_Operator_out1694_out1 XOR Logical_Operator_out1758_out1;

  Logical_Operator_out1951_out1 <= Logical_Operator_out1695_out1 XOR Logical_Operator_out1759_out1;

  Logical_Operator_out1952_out1 <= Logical_Operator_out1696_out1 XOR Logical_Operator_out1760_out1;

  Logical_Operator_out1953_out1 <= Logical_Operator_out1697_out1 XOR Logical_Operator_out1761_out1;

  Logical_Operator_out1954_out1 <= Logical_Operator_out1698_out1 XOR Logical_Operator_out1762_out1;

  Logical_Operator_out1955_out1 <= Logical_Operator_out1699_out1 XOR Logical_Operator_out1763_out1;

  Logical_Operator_out1956_out1 <= Logical_Operator_out1700_out1 XOR Logical_Operator_out1764_out1;

  Logical_Operator_out1957_out1 <= Logical_Operator_out1701_out1 XOR Logical_Operator_out1765_out1;

  Logical_Operator_out1958_out1 <= Logical_Operator_out1702_out1 XOR Logical_Operator_out1766_out1;

  Logical_Operator_out1959_out1 <= Logical_Operator_out1703_out1 XOR Logical_Operator_out1767_out1;

  Logical_Operator_out1960_out1 <= Logical_Operator_out1704_out1 XOR Logical_Operator_out1768_out1;

  Logical_Operator_out1961_out1 <= Logical_Operator_out1705_out1 XOR Logical_Operator_out1769_out1;

  Logical_Operator_out1962_out1 <= Logical_Operator_out1706_out1 XOR Logical_Operator_out1770_out1;

  Logical_Operator_out1963_out1 <= Logical_Operator_out1707_out1 XOR Logical_Operator_out1771_out1;

  Logical_Operator_out1964_out1 <= Logical_Operator_out1708_out1 XOR Logical_Operator_out1772_out1;

  Logical_Operator_out1965_out1 <= Logical_Operator_out1709_out1 XOR Logical_Operator_out1773_out1;

  Logical_Operator_out1966_out1 <= Logical_Operator_out1710_out1 XOR Logical_Operator_out1774_out1;

  Logical_Operator_out1967_out1 <= Logical_Operator_out1711_out1 XOR Logical_Operator_out1775_out1;

  Logical_Operator_out1968_out1 <= Logical_Operator_out1712_out1 XOR Logical_Operator_out1776_out1;

  Logical_Operator_out1969_out1 <= Logical_Operator_out1713_out1 XOR Logical_Operator_out1777_out1;

  Logical_Operator_out1970_out1 <= Logical_Operator_out1714_out1 XOR Logical_Operator_out1778_out1;

  Logical_Operator_out1971_out1 <= Logical_Operator_out1715_out1 XOR Logical_Operator_out1779_out1;

  Logical_Operator_out1972_out1 <= Logical_Operator_out1716_out1 XOR Logical_Operator_out1780_out1;

  Logical_Operator_out1973_out1 <= Logical_Operator_out1717_out1 XOR Logical_Operator_out1781_out1;

  Logical_Operator_out1974_out1 <= Logical_Operator_out1718_out1 XOR Logical_Operator_out1782_out1;

  Logical_Operator_out1975_out1 <= Logical_Operator_out1719_out1 XOR Logical_Operator_out1783_out1;

  Logical_Operator_out1976_out1 <= Logical_Operator_out1720_out1 XOR Logical_Operator_out1784_out1;

  Logical_Operator_out1977_out1 <= Logical_Operator_out1721_out1 XOR Logical_Operator_out1785_out1;

  Logical_Operator_out1978_out1 <= Logical_Operator_out1722_out1 XOR Logical_Operator_out1786_out1;

  Logical_Operator_out1979_out1 <= Logical_Operator_out1723_out1 XOR Logical_Operator_out1787_out1;

  Logical_Operator_out1980_out1 <= Logical_Operator_out1724_out1 XOR Logical_Operator_out1788_out1;

  Logical_Operator_out1981_out1 <= Logical_Operator_out1725_out1 XOR Logical_Operator_out1789_out1;

  Logical_Operator_out1982_out1 <= Logical_Operator_out1726_out1 XOR Logical_Operator_out1790_out1;

  Logical_Operator_out1983_out1 <= Logical_Operator_out1727_out1 XOR Logical_Operator_out1791_out1;

  Logical_Operator_out1984_out1 <= Logical_Operator_out1728_out1 XOR Logical_Operator_out1792_out1;

  Logical_Operator_out1985_out1 <= Logical_Operator_out1441_out1 XOR Logical_Operator_out1505_out1;

  Logical_Operator_out1986_out1 <= Logical_Operator_out1442_out1 XOR Logical_Operator_out1506_out1;

  Logical_Operator_out1987_out1 <= Logical_Operator_out1443_out1 XOR Logical_Operator_out1507_out1;

  Logical_Operator_out1988_out1 <= Logical_Operator_out1444_out1 XOR Logical_Operator_out1508_out1;

  Logical_Operator_out1989_out1 <= Logical_Operator_out1445_out1 XOR Logical_Operator_out1509_out1;

  Logical_Operator_out1990_out1 <= Logical_Operator_out1446_out1 XOR Logical_Operator_out1510_out1;

  Logical_Operator_out1991_out1 <= Logical_Operator_out1447_out1 XOR Logical_Operator_out1511_out1;

  Logical_Operator_out1992_out1 <= Logical_Operator_out1448_out1 XOR Logical_Operator_out1512_out1;

  Logical_Operator_out1993_out1 <= Logical_Operator_out1449_out1 XOR Logical_Operator_out1513_out1;

  Logical_Operator_out1994_out1 <= Logical_Operator_out1450_out1 XOR Logical_Operator_out1514_out1;

  Logical_Operator_out1995_out1 <= Logical_Operator_out1451_out1 XOR Logical_Operator_out1515_out1;

  Logical_Operator_out1996_out1 <= Logical_Operator_out1452_out1 XOR Logical_Operator_out1516_out1;

  Logical_Operator_out1997_out1 <= Logical_Operator_out1453_out1 XOR Logical_Operator_out1517_out1;

  Logical_Operator_out1998_out1 <= Logical_Operator_out1454_out1 XOR Logical_Operator_out1518_out1;

  Logical_Operator_out1999_out1 <= Logical_Operator_out1455_out1 XOR Logical_Operator_out1519_out1;

  Logical_Operator_out2000_out1 <= Logical_Operator_out1456_out1 XOR Logical_Operator_out1520_out1;

  Logical_Operator_out2001_out1 <= Logical_Operator_out1457_out1 XOR Logical_Operator_out1521_out1;

  Logical_Operator_out2002_out1 <= Logical_Operator_out1458_out1 XOR Logical_Operator_out1522_out1;

  Logical_Operator_out2003_out1 <= Logical_Operator_out1459_out1 XOR Logical_Operator_out1523_out1;

  Logical_Operator_out2004_out1 <= Logical_Operator_out1460_out1 XOR Logical_Operator_out1524_out1;

  Logical_Operator_out2005_out1 <= Logical_Operator_out1461_out1 XOR Logical_Operator_out1525_out1;

  Logical_Operator_out2006_out1 <= Logical_Operator_out1462_out1 XOR Logical_Operator_out1526_out1;

  Logical_Operator_out2007_out1 <= Logical_Operator_out1463_out1 XOR Logical_Operator_out1527_out1;

  Logical_Operator_out2008_out1 <= Logical_Operator_out1464_out1 XOR Logical_Operator_out1528_out1;

  Logical_Operator_out2009_out1 <= Logical_Operator_out1465_out1 XOR Logical_Operator_out1529_out1;

  Logical_Operator_out2010_out1 <= Logical_Operator_out1466_out1 XOR Logical_Operator_out1530_out1;

  Logical_Operator_out2011_out1 <= Logical_Operator_out1467_out1 XOR Logical_Operator_out1531_out1;

  Logical_Operator_out2012_out1 <= Logical_Operator_out1468_out1 XOR Logical_Operator_out1532_out1;

  Logical_Operator_out2013_out1 <= Logical_Operator_out1469_out1 XOR Logical_Operator_out1533_out1;

  Logical_Operator_out2014_out1 <= Logical_Operator_out1470_out1 XOR Logical_Operator_out1534_out1;

  Logical_Operator_out2015_out1 <= Logical_Operator_out1471_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out2016_out1 <= Logical_Operator_out1472_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out2017_out1 <= Logical_Operator_out1201_out1 XOR Logical_Operator_out1265_out1;

  Logical_Operator_out2018_out1 <= Logical_Operator_out1202_out1 XOR Logical_Operator_out1266_out1;

  Logical_Operator_out2019_out1 <= Logical_Operator_out1203_out1 XOR Logical_Operator_out1267_out1;

  Logical_Operator_out2020_out1 <= Logical_Operator_out1204_out1 XOR Logical_Operator_out1268_out1;

  Logical_Operator_out2021_out1 <= Logical_Operator_out1205_out1 XOR Logical_Operator_out1269_out1;

  Logical_Operator_out2022_out1 <= Logical_Operator_out1206_out1 XOR Logical_Operator_out1270_out1;

  Logical_Operator_out2023_out1 <= Logical_Operator_out1207_out1 XOR Logical_Operator_out1271_out1;

  Logical_Operator_out2024_out1 <= Logical_Operator_out1208_out1 XOR Logical_Operator_out1272_out1;

  Logical_Operator_out2025_out1 <= Logical_Operator_out1209_out1 XOR Logical_Operator_out1273_out1;

  Logical_Operator_out2026_out1 <= Logical_Operator_out1210_out1 XOR Logical_Operator_out1274_out1;

  Logical_Operator_out2027_out1 <= Logical_Operator_out1211_out1 XOR Logical_Operator_out1275_out1;

  Logical_Operator_out2028_out1 <= Logical_Operator_out1212_out1 XOR Logical_Operator_out1276_out1;

  Logical_Operator_out2029_out1 <= Logical_Operator_out1213_out1 XOR Logical_Operator_out1277_out1;

  Logical_Operator_out2030_out1 <= Logical_Operator_out1214_out1 XOR Logical_Operator_out1278_out1;

  Logical_Operator_out2031_out1 <= Logical_Operator_out1215_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out2032_out1 <= Logical_Operator_out1216_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out2033_out1 <= Logical_Operator_out953_out1 XOR Logical_Operator_out1017_out1;

  Logical_Operator_out2034_out1 <= Logical_Operator_out954_out1 XOR Logical_Operator_out1018_out1;

  Logical_Operator_out2035_out1 <= Logical_Operator_out955_out1 XOR Logical_Operator_out1019_out1;

  Logical_Operator_out2036_out1 <= Logical_Operator_out956_out1 XOR Logical_Operator_out1020_out1;

  Logical_Operator_out2037_out1 <= Logical_Operator_out957_out1 XOR Logical_Operator_out1021_out1;

  Logical_Operator_out2038_out1 <= Logical_Operator_out958_out1 XOR Logical_Operator_out1022_out1;

  Logical_Operator_out2039_out1 <= Logical_Operator_out959_out1 XOR Logical_Operator_out1023_out1;

  Logical_Operator_out2040_out1 <= Logical_Operator_out960_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out2041_out1 <= Logical_Operator_out701_out1 XOR Logical_Operator_out765_out1;

  Logical_Operator_out2042_out1 <= Logical_Operator_out702_out1 XOR Logical_Operator_out766_out1;

  Logical_Operator_out2043_out1 <= Logical_Operator_out703_out1 XOR Logical_Operator_out767_out1;

  Logical_Operator_out2044_out1 <= Logical_Operator_out704_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out2045_out1 <= Logical_Operator_out447_out1 XOR Logical_Operator_out511_out1;

  Logical_Operator_out2046_out1 <= Logical_Operator_out448_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out2047_out1 <= Logical_Operator_out192_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out2048_out1 <= in384 XOR in512;

  Logical_Operator_out2049_out1 <= Logical_Operator_out1793_out1 XOR Logical_Operator_out1921_out1;

  Logical_Operator_out2050_out1 <= Logical_Operator_out1794_out1 XOR Logical_Operator_out1922_out1;

  Logical_Operator_out2051_out1 <= Logical_Operator_out1795_out1 XOR Logical_Operator_out1923_out1;

  Logical_Operator_out2052_out1 <= Logical_Operator_out1796_out1 XOR Logical_Operator_out1924_out1;

  Logical_Operator_out2053_out1 <= Logical_Operator_out1797_out1 XOR Logical_Operator_out1925_out1;

  Logical_Operator_out2054_out1 <= Logical_Operator_out1798_out1 XOR Logical_Operator_out1926_out1;

  Logical_Operator_out2055_out1 <= Logical_Operator_out1799_out1 XOR Logical_Operator_out1927_out1;

  Logical_Operator_out2056_out1 <= Logical_Operator_out1800_out1 XOR Logical_Operator_out1928_out1;

  Logical_Operator_out2057_out1 <= Logical_Operator_out1801_out1 XOR Logical_Operator_out1929_out1;

  Logical_Operator_out2058_out1 <= Logical_Operator_out1802_out1 XOR Logical_Operator_out1930_out1;

  Logical_Operator_out2059_out1 <= Logical_Operator_out1803_out1 XOR Logical_Operator_out1931_out1;

  Logical_Operator_out2060_out1 <= Logical_Operator_out1804_out1 XOR Logical_Operator_out1932_out1;

  Logical_Operator_out2061_out1 <= Logical_Operator_out1805_out1 XOR Logical_Operator_out1933_out1;

  Logical_Operator_out2062_out1 <= Logical_Operator_out1806_out1 XOR Logical_Operator_out1934_out1;

  Logical_Operator_out2063_out1 <= Logical_Operator_out1807_out1 XOR Logical_Operator_out1935_out1;

  Logical_Operator_out2064_out1 <= Logical_Operator_out1808_out1 XOR Logical_Operator_out1936_out1;

  Logical_Operator_out2065_out1 <= Logical_Operator_out1809_out1 XOR Logical_Operator_out1937_out1;

  Logical_Operator_out2066_out1 <= Logical_Operator_out1810_out1 XOR Logical_Operator_out1938_out1;

  Logical_Operator_out2067_out1 <= Logical_Operator_out1811_out1 XOR Logical_Operator_out1939_out1;

  Logical_Operator_out2068_out1 <= Logical_Operator_out1812_out1 XOR Logical_Operator_out1940_out1;

  Logical_Operator_out2069_out1 <= Logical_Operator_out1813_out1 XOR Logical_Operator_out1941_out1;

  Logical_Operator_out2070_out1 <= Logical_Operator_out1814_out1 XOR Logical_Operator_out1942_out1;

  Logical_Operator_out2071_out1 <= Logical_Operator_out1815_out1 XOR Logical_Operator_out1943_out1;

  Logical_Operator_out2072_out1 <= Logical_Operator_out1816_out1 XOR Logical_Operator_out1944_out1;

  Logical_Operator_out2073_out1 <= Logical_Operator_out1817_out1 XOR Logical_Operator_out1945_out1;

  Logical_Operator_out2074_out1 <= Logical_Operator_out1818_out1 XOR Logical_Operator_out1946_out1;

  Logical_Operator_out2075_out1 <= Logical_Operator_out1819_out1 XOR Logical_Operator_out1947_out1;

  Logical_Operator_out2076_out1 <= Logical_Operator_out1820_out1 XOR Logical_Operator_out1948_out1;

  Logical_Operator_out2077_out1 <= Logical_Operator_out1821_out1 XOR Logical_Operator_out1949_out1;

  Logical_Operator_out2078_out1 <= Logical_Operator_out1822_out1 XOR Logical_Operator_out1950_out1;

  Logical_Operator_out2079_out1 <= Logical_Operator_out1823_out1 XOR Logical_Operator_out1951_out1;

  Logical_Operator_out2080_out1 <= Logical_Operator_out1824_out1 XOR Logical_Operator_out1952_out1;

  Logical_Operator_out2081_out1 <= Logical_Operator_out1825_out1 XOR Logical_Operator_out1953_out1;

  Logical_Operator_out2082_out1 <= Logical_Operator_out1826_out1 XOR Logical_Operator_out1954_out1;

  Logical_Operator_out2083_out1 <= Logical_Operator_out1827_out1 XOR Logical_Operator_out1955_out1;

  Logical_Operator_out2084_out1 <= Logical_Operator_out1828_out1 XOR Logical_Operator_out1956_out1;

  Logical_Operator_out2085_out1 <= Logical_Operator_out1829_out1 XOR Logical_Operator_out1957_out1;

  Logical_Operator_out2086_out1 <= Logical_Operator_out1830_out1 XOR Logical_Operator_out1958_out1;

  Logical_Operator_out2087_out1 <= Logical_Operator_out1831_out1 XOR Logical_Operator_out1959_out1;

  Logical_Operator_out2088_out1 <= Logical_Operator_out1832_out1 XOR Logical_Operator_out1960_out1;

  Logical_Operator_out2089_out1 <= Logical_Operator_out1833_out1 XOR Logical_Operator_out1961_out1;

  Logical_Operator_out2090_out1 <= Logical_Operator_out1834_out1 XOR Logical_Operator_out1962_out1;

  Logical_Operator_out2091_out1 <= Logical_Operator_out1835_out1 XOR Logical_Operator_out1963_out1;

  Logical_Operator_out2092_out1 <= Logical_Operator_out1836_out1 XOR Logical_Operator_out1964_out1;

  Logical_Operator_out2093_out1 <= Logical_Operator_out1837_out1 XOR Logical_Operator_out1965_out1;

  Logical_Operator_out2094_out1 <= Logical_Operator_out1838_out1 XOR Logical_Operator_out1966_out1;

  Logical_Operator_out2095_out1 <= Logical_Operator_out1839_out1 XOR Logical_Operator_out1967_out1;

  Logical_Operator_out2096_out1 <= Logical_Operator_out1840_out1 XOR Logical_Operator_out1968_out1;

  Logical_Operator_out2097_out1 <= Logical_Operator_out1841_out1 XOR Logical_Operator_out1969_out1;

  Logical_Operator_out2098_out1 <= Logical_Operator_out1842_out1 XOR Logical_Operator_out1970_out1;

  Logical_Operator_out2099_out1 <= Logical_Operator_out1843_out1 XOR Logical_Operator_out1971_out1;

  Logical_Operator_out2100_out1 <= Logical_Operator_out1844_out1 XOR Logical_Operator_out1972_out1;

  Logical_Operator_out2101_out1 <= Logical_Operator_out1845_out1 XOR Logical_Operator_out1973_out1;

  Logical_Operator_out2102_out1 <= Logical_Operator_out1846_out1 XOR Logical_Operator_out1974_out1;

  Logical_Operator_out2103_out1 <= Logical_Operator_out1847_out1 XOR Logical_Operator_out1975_out1;

  Logical_Operator_out2104_out1 <= Logical_Operator_out1848_out1 XOR Logical_Operator_out1976_out1;

  Logical_Operator_out2105_out1 <= Logical_Operator_out1849_out1 XOR Logical_Operator_out1977_out1;

  Logical_Operator_out2106_out1 <= Logical_Operator_out1850_out1 XOR Logical_Operator_out1978_out1;

  Logical_Operator_out2107_out1 <= Logical_Operator_out1851_out1 XOR Logical_Operator_out1979_out1;

  Logical_Operator_out2108_out1 <= Logical_Operator_out1852_out1 XOR Logical_Operator_out1980_out1;

  Logical_Operator_out2109_out1 <= Logical_Operator_out1853_out1 XOR Logical_Operator_out1981_out1;

  Logical_Operator_out2110_out1 <= Logical_Operator_out1854_out1 XOR Logical_Operator_out1982_out1;

  Logical_Operator_out2111_out1 <= Logical_Operator_out1855_out1 XOR Logical_Operator_out1983_out1;

  Logical_Operator_out2112_out1 <= Logical_Operator_out1856_out1 XOR Logical_Operator_out1984_out1;

  Logical_Operator_out2113_out1 <= Logical_Operator_out1857_out1 XOR Logical_Operator_out1985_out1;

  Logical_Operator_out2114_out1 <= Logical_Operator_out1858_out1 XOR Logical_Operator_out1986_out1;

  Logical_Operator_out2115_out1 <= Logical_Operator_out1859_out1 XOR Logical_Operator_out1987_out1;

  Logical_Operator_out2116_out1 <= Logical_Operator_out1860_out1 XOR Logical_Operator_out1988_out1;

  Logical_Operator_out2117_out1 <= Logical_Operator_out1861_out1 XOR Logical_Operator_out1989_out1;

  Logical_Operator_out2118_out1 <= Logical_Operator_out1862_out1 XOR Logical_Operator_out1990_out1;

  Logical_Operator_out2119_out1 <= Logical_Operator_out1863_out1 XOR Logical_Operator_out1991_out1;

  Logical_Operator_out2120_out1 <= Logical_Operator_out1864_out1 XOR Logical_Operator_out1992_out1;

  Logical_Operator_out2121_out1 <= Logical_Operator_out1865_out1 XOR Logical_Operator_out1993_out1;

  Logical_Operator_out2122_out1 <= Logical_Operator_out1866_out1 XOR Logical_Operator_out1994_out1;

  Logical_Operator_out2123_out1 <= Logical_Operator_out1867_out1 XOR Logical_Operator_out1995_out1;

  Logical_Operator_out2124_out1 <= Logical_Operator_out1868_out1 XOR Logical_Operator_out1996_out1;

  Logical_Operator_out2125_out1 <= Logical_Operator_out1869_out1 XOR Logical_Operator_out1997_out1;

  Logical_Operator_out2126_out1 <= Logical_Operator_out1870_out1 XOR Logical_Operator_out1998_out1;

  Logical_Operator_out2127_out1 <= Logical_Operator_out1871_out1 XOR Logical_Operator_out1999_out1;

  Logical_Operator_out2128_out1 <= Logical_Operator_out1872_out1 XOR Logical_Operator_out2000_out1;

  Logical_Operator_out2129_out1 <= Logical_Operator_out1873_out1 XOR Logical_Operator_out2001_out1;

  Logical_Operator_out2130_out1 <= Logical_Operator_out1874_out1 XOR Logical_Operator_out2002_out1;

  Logical_Operator_out2131_out1 <= Logical_Operator_out1875_out1 XOR Logical_Operator_out2003_out1;

  Logical_Operator_out2132_out1 <= Logical_Operator_out1876_out1 XOR Logical_Operator_out2004_out1;

  Logical_Operator_out2133_out1 <= Logical_Operator_out1877_out1 XOR Logical_Operator_out2005_out1;

  Logical_Operator_out2134_out1 <= Logical_Operator_out1878_out1 XOR Logical_Operator_out2006_out1;

  Logical_Operator_out2135_out1 <= Logical_Operator_out1879_out1 XOR Logical_Operator_out2007_out1;

  Logical_Operator_out2136_out1 <= Logical_Operator_out1880_out1 XOR Logical_Operator_out2008_out1;

  Logical_Operator_out2137_out1 <= Logical_Operator_out1881_out1 XOR Logical_Operator_out2009_out1;

  Logical_Operator_out2138_out1 <= Logical_Operator_out1882_out1 XOR Logical_Operator_out2010_out1;

  Logical_Operator_out2139_out1 <= Logical_Operator_out1883_out1 XOR Logical_Operator_out2011_out1;

  Logical_Operator_out2140_out1 <= Logical_Operator_out1884_out1 XOR Logical_Operator_out2012_out1;

  Logical_Operator_out2141_out1 <= Logical_Operator_out1885_out1 XOR Logical_Operator_out2013_out1;

  Logical_Operator_out2142_out1 <= Logical_Operator_out1886_out1 XOR Logical_Operator_out2014_out1;

  Logical_Operator_out2143_out1 <= Logical_Operator_out1887_out1 XOR Logical_Operator_out2015_out1;

  Logical_Operator_out2144_out1 <= Logical_Operator_out1888_out1 XOR Logical_Operator_out2016_out1;

  Logical_Operator_out2145_out1 <= Logical_Operator_out1889_out1 XOR Logical_Operator_out2017_out1;

  Logical_Operator_out2146_out1 <= Logical_Operator_out1890_out1 XOR Logical_Operator_out2018_out1;

  Logical_Operator_out2147_out1 <= Logical_Operator_out1891_out1 XOR Logical_Operator_out2019_out1;

  Logical_Operator_out2148_out1 <= Logical_Operator_out1892_out1 XOR Logical_Operator_out2020_out1;

  Logical_Operator_out2149_out1 <= Logical_Operator_out1893_out1 XOR Logical_Operator_out2021_out1;

  Logical_Operator_out2150_out1 <= Logical_Operator_out1894_out1 XOR Logical_Operator_out2022_out1;

  Logical_Operator_out2151_out1 <= Logical_Operator_out1895_out1 XOR Logical_Operator_out2023_out1;

  Logical_Operator_out2152_out1 <= Logical_Operator_out1896_out1 XOR Logical_Operator_out2024_out1;

  Logical_Operator_out2153_out1 <= Logical_Operator_out1897_out1 XOR Logical_Operator_out2025_out1;

  Logical_Operator_out2154_out1 <= Logical_Operator_out1898_out1 XOR Logical_Operator_out2026_out1;

  Logical_Operator_out2155_out1 <= Logical_Operator_out1899_out1 XOR Logical_Operator_out2027_out1;

  Logical_Operator_out2156_out1 <= Logical_Operator_out1900_out1 XOR Logical_Operator_out2028_out1;

  Logical_Operator_out2157_out1 <= Logical_Operator_out1901_out1 XOR Logical_Operator_out2029_out1;

  Logical_Operator_out2158_out1 <= Logical_Operator_out1902_out1 XOR Logical_Operator_out2030_out1;

  Logical_Operator_out2159_out1 <= Logical_Operator_out1903_out1 XOR Logical_Operator_out2031_out1;

  Logical_Operator_out2160_out1 <= Logical_Operator_out1904_out1 XOR Logical_Operator_out2032_out1;

  Logical_Operator_out2161_out1 <= Logical_Operator_out1905_out1 XOR Logical_Operator_out2033_out1;

  Logical_Operator_out2162_out1 <= Logical_Operator_out1906_out1 XOR Logical_Operator_out2034_out1;

  Logical_Operator_out2163_out1 <= Logical_Operator_out1907_out1 XOR Logical_Operator_out2035_out1;

  Logical_Operator_out2164_out1 <= Logical_Operator_out1908_out1 XOR Logical_Operator_out2036_out1;

  Logical_Operator_out2165_out1 <= Logical_Operator_out1909_out1 XOR Logical_Operator_out2037_out1;

  Logical_Operator_out2166_out1 <= Logical_Operator_out1910_out1 XOR Logical_Operator_out2038_out1;

  Logical_Operator_out2167_out1 <= Logical_Operator_out1911_out1 XOR Logical_Operator_out2039_out1;

  Logical_Operator_out2168_out1 <= Logical_Operator_out1912_out1 XOR Logical_Operator_out2040_out1;

  Logical_Operator_out2169_out1 <= Logical_Operator_out1913_out1 XOR Logical_Operator_out2041_out1;

  Logical_Operator_out2170_out1 <= Logical_Operator_out1914_out1 XOR Logical_Operator_out2042_out1;

  Logical_Operator_out2171_out1 <= Logical_Operator_out1915_out1 XOR Logical_Operator_out2043_out1;

  Logical_Operator_out2172_out1 <= Logical_Operator_out1916_out1 XOR Logical_Operator_out2044_out1;

  Logical_Operator_out2173_out1 <= Logical_Operator_out1917_out1 XOR Logical_Operator_out2045_out1;

  Logical_Operator_out2174_out1 <= Logical_Operator_out1918_out1 XOR Logical_Operator_out2046_out1;

  Logical_Operator_out2175_out1 <= Logical_Operator_out1919_out1 XOR Logical_Operator_out2047_out1;

  Logical_Operator_out2176_out1 <= Logical_Operator_out1920_out1 XOR Logical_Operator_out2048_out1;

  Logical_Operator_out2177_out1 <= Logical_Operator_out1601_out1 XOR Logical_Operator_out1729_out1;

  Logical_Operator_out2178_out1 <= Logical_Operator_out1602_out1 XOR Logical_Operator_out1730_out1;

  Logical_Operator_out2179_out1 <= Logical_Operator_out1603_out1 XOR Logical_Operator_out1731_out1;

  Logical_Operator_out2180_out1 <= Logical_Operator_out1604_out1 XOR Logical_Operator_out1732_out1;

  Logical_Operator_out2181_out1 <= Logical_Operator_out1605_out1 XOR Logical_Operator_out1733_out1;

  Logical_Operator_out2182_out1 <= Logical_Operator_out1606_out1 XOR Logical_Operator_out1734_out1;

  Logical_Operator_out2183_out1 <= Logical_Operator_out1607_out1 XOR Logical_Operator_out1735_out1;

  Logical_Operator_out2184_out1 <= Logical_Operator_out1608_out1 XOR Logical_Operator_out1736_out1;

  Logical_Operator_out2185_out1 <= Logical_Operator_out1609_out1 XOR Logical_Operator_out1737_out1;

  Logical_Operator_out2186_out1 <= Logical_Operator_out1610_out1 XOR Logical_Operator_out1738_out1;

  Logical_Operator_out2187_out1 <= Logical_Operator_out1611_out1 XOR Logical_Operator_out1739_out1;

  Logical_Operator_out2188_out1 <= Logical_Operator_out1612_out1 XOR Logical_Operator_out1740_out1;

  Logical_Operator_out2189_out1 <= Logical_Operator_out1613_out1 XOR Logical_Operator_out1741_out1;

  Logical_Operator_out2190_out1 <= Logical_Operator_out1614_out1 XOR Logical_Operator_out1742_out1;

  Logical_Operator_out2191_out1 <= Logical_Operator_out1615_out1 XOR Logical_Operator_out1743_out1;

  Logical_Operator_out2192_out1 <= Logical_Operator_out1616_out1 XOR Logical_Operator_out1744_out1;

  Logical_Operator_out2193_out1 <= Logical_Operator_out1617_out1 XOR Logical_Operator_out1745_out1;

  Logical_Operator_out2194_out1 <= Logical_Operator_out1618_out1 XOR Logical_Operator_out1746_out1;

  Logical_Operator_out2195_out1 <= Logical_Operator_out1619_out1 XOR Logical_Operator_out1747_out1;

  Logical_Operator_out2196_out1 <= Logical_Operator_out1620_out1 XOR Logical_Operator_out1748_out1;

  Logical_Operator_out2197_out1 <= Logical_Operator_out1621_out1 XOR Logical_Operator_out1749_out1;

  Logical_Operator_out2198_out1 <= Logical_Operator_out1622_out1 XOR Logical_Operator_out1750_out1;

  Logical_Operator_out2199_out1 <= Logical_Operator_out1623_out1 XOR Logical_Operator_out1751_out1;

  Logical_Operator_out2200_out1 <= Logical_Operator_out1624_out1 XOR Logical_Operator_out1752_out1;

  Logical_Operator_out2201_out1 <= Logical_Operator_out1625_out1 XOR Logical_Operator_out1753_out1;

  Logical_Operator_out2202_out1 <= Logical_Operator_out1626_out1 XOR Logical_Operator_out1754_out1;

  Logical_Operator_out2203_out1 <= Logical_Operator_out1627_out1 XOR Logical_Operator_out1755_out1;

  Logical_Operator_out2204_out1 <= Logical_Operator_out1628_out1 XOR Logical_Operator_out1756_out1;

  Logical_Operator_out2205_out1 <= Logical_Operator_out1629_out1 XOR Logical_Operator_out1757_out1;

  Logical_Operator_out2206_out1 <= Logical_Operator_out1630_out1 XOR Logical_Operator_out1758_out1;

  Logical_Operator_out2207_out1 <= Logical_Operator_out1631_out1 XOR Logical_Operator_out1759_out1;

  Logical_Operator_out2208_out1 <= Logical_Operator_out1632_out1 XOR Logical_Operator_out1760_out1;

  Logical_Operator_out2209_out1 <= Logical_Operator_out1633_out1 XOR Logical_Operator_out1761_out1;

  Logical_Operator_out2210_out1 <= Logical_Operator_out1634_out1 XOR Logical_Operator_out1762_out1;

  Logical_Operator_out2211_out1 <= Logical_Operator_out1635_out1 XOR Logical_Operator_out1763_out1;

  Logical_Operator_out2212_out1 <= Logical_Operator_out1636_out1 XOR Logical_Operator_out1764_out1;

  Logical_Operator_out2213_out1 <= Logical_Operator_out1637_out1 XOR Logical_Operator_out1765_out1;

  Logical_Operator_out2214_out1 <= Logical_Operator_out1638_out1 XOR Logical_Operator_out1766_out1;

  Logical_Operator_out2215_out1 <= Logical_Operator_out1639_out1 XOR Logical_Operator_out1767_out1;

  Logical_Operator_out2216_out1 <= Logical_Operator_out1640_out1 XOR Logical_Operator_out1768_out1;

  Logical_Operator_out2217_out1 <= Logical_Operator_out1641_out1 XOR Logical_Operator_out1769_out1;

  Logical_Operator_out2218_out1 <= Logical_Operator_out1642_out1 XOR Logical_Operator_out1770_out1;

  Logical_Operator_out2219_out1 <= Logical_Operator_out1643_out1 XOR Logical_Operator_out1771_out1;

  Logical_Operator_out2220_out1 <= Logical_Operator_out1644_out1 XOR Logical_Operator_out1772_out1;

  Logical_Operator_out2221_out1 <= Logical_Operator_out1645_out1 XOR Logical_Operator_out1773_out1;

  Logical_Operator_out2222_out1 <= Logical_Operator_out1646_out1 XOR Logical_Operator_out1774_out1;

  Logical_Operator_out2223_out1 <= Logical_Operator_out1647_out1 XOR Logical_Operator_out1775_out1;

  Logical_Operator_out2224_out1 <= Logical_Operator_out1648_out1 XOR Logical_Operator_out1776_out1;

  Logical_Operator_out2225_out1 <= Logical_Operator_out1649_out1 XOR Logical_Operator_out1777_out1;

  Logical_Operator_out2226_out1 <= Logical_Operator_out1650_out1 XOR Logical_Operator_out1778_out1;

  Logical_Operator_out2227_out1 <= Logical_Operator_out1651_out1 XOR Logical_Operator_out1779_out1;

  Logical_Operator_out2228_out1 <= Logical_Operator_out1652_out1 XOR Logical_Operator_out1780_out1;

  Logical_Operator_out2229_out1 <= Logical_Operator_out1653_out1 XOR Logical_Operator_out1781_out1;

  Logical_Operator_out2230_out1 <= Logical_Operator_out1654_out1 XOR Logical_Operator_out1782_out1;

  Logical_Operator_out2231_out1 <= Logical_Operator_out1655_out1 XOR Logical_Operator_out1783_out1;

  Logical_Operator_out2232_out1 <= Logical_Operator_out1656_out1 XOR Logical_Operator_out1784_out1;

  Logical_Operator_out2233_out1 <= Logical_Operator_out1657_out1 XOR Logical_Operator_out1785_out1;

  Logical_Operator_out2234_out1 <= Logical_Operator_out1658_out1 XOR Logical_Operator_out1786_out1;

  Logical_Operator_out2235_out1 <= Logical_Operator_out1659_out1 XOR Logical_Operator_out1787_out1;

  Logical_Operator_out2236_out1 <= Logical_Operator_out1660_out1 XOR Logical_Operator_out1788_out1;

  Logical_Operator_out2237_out1 <= Logical_Operator_out1661_out1 XOR Logical_Operator_out1789_out1;

  Logical_Operator_out2238_out1 <= Logical_Operator_out1662_out1 XOR Logical_Operator_out1790_out1;

  Logical_Operator_out2239_out1 <= Logical_Operator_out1663_out1 XOR Logical_Operator_out1791_out1;

  Logical_Operator_out2240_out1 <= Logical_Operator_out1664_out1 XOR Logical_Operator_out1792_out1;

  Logical_Operator_out2241_out1 <= Logical_Operator_out1377_out1 XOR Logical_Operator_out1505_out1;

  Logical_Operator_out2242_out1 <= Logical_Operator_out1378_out1 XOR Logical_Operator_out1506_out1;

  Logical_Operator_out2243_out1 <= Logical_Operator_out1379_out1 XOR Logical_Operator_out1507_out1;

  Logical_Operator_out2244_out1 <= Logical_Operator_out1380_out1 XOR Logical_Operator_out1508_out1;

  Logical_Operator_out2245_out1 <= Logical_Operator_out1381_out1 XOR Logical_Operator_out1509_out1;

  Logical_Operator_out2246_out1 <= Logical_Operator_out1382_out1 XOR Logical_Operator_out1510_out1;

  Logical_Operator_out2247_out1 <= Logical_Operator_out1383_out1 XOR Logical_Operator_out1511_out1;

  Logical_Operator_out2248_out1 <= Logical_Operator_out1384_out1 XOR Logical_Operator_out1512_out1;

  Logical_Operator_out2249_out1 <= Logical_Operator_out1385_out1 XOR Logical_Operator_out1513_out1;

  Logical_Operator_out2250_out1 <= Logical_Operator_out1386_out1 XOR Logical_Operator_out1514_out1;

  Logical_Operator_out2251_out1 <= Logical_Operator_out1387_out1 XOR Logical_Operator_out1515_out1;

  Logical_Operator_out2252_out1 <= Logical_Operator_out1388_out1 XOR Logical_Operator_out1516_out1;

  Logical_Operator_out2253_out1 <= Logical_Operator_out1389_out1 XOR Logical_Operator_out1517_out1;

  Logical_Operator_out2254_out1 <= Logical_Operator_out1390_out1 XOR Logical_Operator_out1518_out1;

  Logical_Operator_out2255_out1 <= Logical_Operator_out1391_out1 XOR Logical_Operator_out1519_out1;

  Logical_Operator_out2256_out1 <= Logical_Operator_out1392_out1 XOR Logical_Operator_out1520_out1;

  Logical_Operator_out2257_out1 <= Logical_Operator_out1393_out1 XOR Logical_Operator_out1521_out1;

  Logical_Operator_out2258_out1 <= Logical_Operator_out1394_out1 XOR Logical_Operator_out1522_out1;

  Logical_Operator_out2259_out1 <= Logical_Operator_out1395_out1 XOR Logical_Operator_out1523_out1;

  Logical_Operator_out2260_out1 <= Logical_Operator_out1396_out1 XOR Logical_Operator_out1524_out1;

  Logical_Operator_out2261_out1 <= Logical_Operator_out1397_out1 XOR Logical_Operator_out1525_out1;

  Logical_Operator_out2262_out1 <= Logical_Operator_out1398_out1 XOR Logical_Operator_out1526_out1;

  Logical_Operator_out2263_out1 <= Logical_Operator_out1399_out1 XOR Logical_Operator_out1527_out1;

  Logical_Operator_out2264_out1 <= Logical_Operator_out1400_out1 XOR Logical_Operator_out1528_out1;

  Logical_Operator_out2265_out1 <= Logical_Operator_out1401_out1 XOR Logical_Operator_out1529_out1;

  Logical_Operator_out2266_out1 <= Logical_Operator_out1402_out1 XOR Logical_Operator_out1530_out1;

  Logical_Operator_out2267_out1 <= Logical_Operator_out1403_out1 XOR Logical_Operator_out1531_out1;

  Logical_Operator_out2268_out1 <= Logical_Operator_out1404_out1 XOR Logical_Operator_out1532_out1;

  Logical_Operator_out2269_out1 <= Logical_Operator_out1405_out1 XOR Logical_Operator_out1533_out1;

  Logical_Operator_out2270_out1 <= Logical_Operator_out1406_out1 XOR Logical_Operator_out1534_out1;

  Logical_Operator_out2271_out1 <= Logical_Operator_out1407_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out2272_out1 <= Logical_Operator_out1408_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out2273_out1 <= Logical_Operator_out1137_out1 XOR Logical_Operator_out1265_out1;

  Logical_Operator_out2274_out1 <= Logical_Operator_out1138_out1 XOR Logical_Operator_out1266_out1;

  Logical_Operator_out2275_out1 <= Logical_Operator_out1139_out1 XOR Logical_Operator_out1267_out1;

  Logical_Operator_out2276_out1 <= Logical_Operator_out1140_out1 XOR Logical_Operator_out1268_out1;

  Logical_Operator_out2277_out1 <= Logical_Operator_out1141_out1 XOR Logical_Operator_out1269_out1;

  Logical_Operator_out2278_out1 <= Logical_Operator_out1142_out1 XOR Logical_Operator_out1270_out1;

  Logical_Operator_out2279_out1 <= Logical_Operator_out1143_out1 XOR Logical_Operator_out1271_out1;

  Logical_Operator_out2280_out1 <= Logical_Operator_out1144_out1 XOR Logical_Operator_out1272_out1;

  Logical_Operator_out2281_out1 <= Logical_Operator_out1145_out1 XOR Logical_Operator_out1273_out1;

  Logical_Operator_out2282_out1 <= Logical_Operator_out1146_out1 XOR Logical_Operator_out1274_out1;

  Logical_Operator_out2283_out1 <= Logical_Operator_out1147_out1 XOR Logical_Operator_out1275_out1;

  Logical_Operator_out2284_out1 <= Logical_Operator_out1148_out1 XOR Logical_Operator_out1276_out1;

  Logical_Operator_out2285_out1 <= Logical_Operator_out1149_out1 XOR Logical_Operator_out1277_out1;

  Logical_Operator_out2286_out1 <= Logical_Operator_out1150_out1 XOR Logical_Operator_out1278_out1;

  Logical_Operator_out2287_out1 <= Logical_Operator_out1151_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out2288_out1 <= Logical_Operator_out1152_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out2289_out1 <= Logical_Operator_out889_out1 XOR Logical_Operator_out1017_out1;

  Logical_Operator_out2290_out1 <= Logical_Operator_out890_out1 XOR Logical_Operator_out1018_out1;

  Logical_Operator_out2291_out1 <= Logical_Operator_out891_out1 XOR Logical_Operator_out1019_out1;

  Logical_Operator_out2292_out1 <= Logical_Operator_out892_out1 XOR Logical_Operator_out1020_out1;

  Logical_Operator_out2293_out1 <= Logical_Operator_out893_out1 XOR Logical_Operator_out1021_out1;

  Logical_Operator_out2294_out1 <= Logical_Operator_out894_out1 XOR Logical_Operator_out1022_out1;

  Logical_Operator_out2295_out1 <= Logical_Operator_out895_out1 XOR Logical_Operator_out1023_out1;

  Logical_Operator_out2296_out1 <= Logical_Operator_out896_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out2297_out1 <= Logical_Operator_out637_out1 XOR Logical_Operator_out765_out1;

  Logical_Operator_out2298_out1 <= Logical_Operator_out638_out1 XOR Logical_Operator_out766_out1;

  Logical_Operator_out2299_out1 <= Logical_Operator_out639_out1 XOR Logical_Operator_out767_out1;

  Logical_Operator_out2300_out1 <= Logical_Operator_out640_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out2301_out1 <= Logical_Operator_out383_out1 XOR Logical_Operator_out511_out1;

  Logical_Operator_out2302_out1 <= Logical_Operator_out384_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out2303_out1 <= Logical_Operator_out128_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out2304_out1 <= in256 XOR in512;

  out1 <= Logical_Operator_out2049_out1;

  out2 <= Logical_Operator_out2050_out1;

  out3 <= Logical_Operator_out2051_out1;

  out4 <= Logical_Operator_out2052_out1;

  out5 <= Logical_Operator_out2053_out1;

  out6 <= Logical_Operator_out2054_out1;

  out7 <= Logical_Operator_out2055_out1;

  out8 <= Logical_Operator_out2056_out1;

  out9 <= Logical_Operator_out2057_out1;

  out10 <= Logical_Operator_out2058_out1;

  out11 <= Logical_Operator_out2059_out1;

  out12 <= Logical_Operator_out2060_out1;

  out13 <= Logical_Operator_out2061_out1;

  out14 <= Logical_Operator_out2062_out1;

  out15 <= Logical_Operator_out2063_out1;

  out16 <= Logical_Operator_out2064_out1;

  out17 <= Logical_Operator_out2065_out1;

  out18 <= Logical_Operator_out2066_out1;

  out19 <= Logical_Operator_out2067_out1;

  out20 <= Logical_Operator_out2068_out1;

  out21 <= Logical_Operator_out2069_out1;

  out22 <= Logical_Operator_out2070_out1;

  out23 <= Logical_Operator_out2071_out1;

  out24 <= Logical_Operator_out2072_out1;

  out25 <= Logical_Operator_out2073_out1;

  out26 <= Logical_Operator_out2074_out1;

  out27 <= Logical_Operator_out2075_out1;

  out28 <= Logical_Operator_out2076_out1;

  out29 <= Logical_Operator_out2077_out1;

  out30 <= Logical_Operator_out2078_out1;

  out31 <= Logical_Operator_out2079_out1;

  out32 <= Logical_Operator_out2080_out1;

  out33 <= Logical_Operator_out2081_out1;

  out34 <= Logical_Operator_out2082_out1;

  out35 <= Logical_Operator_out2083_out1;

  out36 <= Logical_Operator_out2084_out1;

  out37 <= Logical_Operator_out2085_out1;

  out38 <= Logical_Operator_out2086_out1;

  out39 <= Logical_Operator_out2087_out1;

  out40 <= Logical_Operator_out2088_out1;

  out41 <= Logical_Operator_out2089_out1;

  out42 <= Logical_Operator_out2090_out1;

  out43 <= Logical_Operator_out2091_out1;

  out44 <= Logical_Operator_out2092_out1;

  out45 <= Logical_Operator_out2093_out1;

  out46 <= Logical_Operator_out2094_out1;

  out47 <= Logical_Operator_out2095_out1;

  out48 <= Logical_Operator_out2096_out1;

  out49 <= Logical_Operator_out2097_out1;

  out50 <= Logical_Operator_out2098_out1;

  out51 <= Logical_Operator_out2099_out1;

  out52 <= Logical_Operator_out2100_out1;

  out53 <= Logical_Operator_out2101_out1;

  out54 <= Logical_Operator_out2102_out1;

  out55 <= Logical_Operator_out2103_out1;

  out56 <= Logical_Operator_out2104_out1;

  out57 <= Logical_Operator_out2105_out1;

  out58 <= Logical_Operator_out2106_out1;

  out59 <= Logical_Operator_out2107_out1;

  out60 <= Logical_Operator_out2108_out1;

  out61 <= Logical_Operator_out2109_out1;

  out62 <= Logical_Operator_out2110_out1;

  out63 <= Logical_Operator_out2111_out1;

  out64 <= Logical_Operator_out2112_out1;

  out65 <= Logical_Operator_out2113_out1;

  out66 <= Logical_Operator_out2114_out1;

  out67 <= Logical_Operator_out2115_out1;

  out68 <= Logical_Operator_out2116_out1;

  out69 <= Logical_Operator_out2117_out1;

  out70 <= Logical_Operator_out2118_out1;

  out71 <= Logical_Operator_out2119_out1;

  out72 <= Logical_Operator_out2120_out1;

  out73 <= Logical_Operator_out2121_out1;

  out74 <= Logical_Operator_out2122_out1;

  out75 <= Logical_Operator_out2123_out1;

  out76 <= Logical_Operator_out2124_out1;

  out77 <= Logical_Operator_out2125_out1;

  out78 <= Logical_Operator_out2126_out1;

  out79 <= Logical_Operator_out2127_out1;

  out80 <= Logical_Operator_out2128_out1;

  out81 <= Logical_Operator_out2129_out1;

  out82 <= Logical_Operator_out2130_out1;

  out83 <= Logical_Operator_out2131_out1;

  out84 <= Logical_Operator_out2132_out1;

  out85 <= Logical_Operator_out2133_out1;

  out86 <= Logical_Operator_out2134_out1;

  out87 <= Logical_Operator_out2135_out1;

  out88 <= Logical_Operator_out2136_out1;

  out89 <= Logical_Operator_out2137_out1;

  out90 <= Logical_Operator_out2138_out1;

  out91 <= Logical_Operator_out2139_out1;

  out92 <= Logical_Operator_out2140_out1;

  out93 <= Logical_Operator_out2141_out1;

  out94 <= Logical_Operator_out2142_out1;

  out95 <= Logical_Operator_out2143_out1;

  out96 <= Logical_Operator_out2144_out1;

  out97 <= Logical_Operator_out2145_out1;

  out98 <= Logical_Operator_out2146_out1;

  out99 <= Logical_Operator_out2147_out1;

  out100 <= Logical_Operator_out2148_out1;

  out101 <= Logical_Operator_out2149_out1;

  out102 <= Logical_Operator_out2150_out1;

  out103 <= Logical_Operator_out2151_out1;

  out104 <= Logical_Operator_out2152_out1;

  out105 <= Logical_Operator_out2153_out1;

  out106 <= Logical_Operator_out2154_out1;

  out107 <= Logical_Operator_out2155_out1;

  out108 <= Logical_Operator_out2156_out1;

  out109 <= Logical_Operator_out2157_out1;

  out110 <= Logical_Operator_out2158_out1;

  out111 <= Logical_Operator_out2159_out1;

  out112 <= Logical_Operator_out2160_out1;

  out113 <= Logical_Operator_out2161_out1;

  out114 <= Logical_Operator_out2162_out1;

  out115 <= Logical_Operator_out2163_out1;

  out116 <= Logical_Operator_out2164_out1;

  out117 <= Logical_Operator_out2165_out1;

  out118 <= Logical_Operator_out2166_out1;

  out119 <= Logical_Operator_out2167_out1;

  out120 <= Logical_Operator_out2168_out1;

  out121 <= Logical_Operator_out2169_out1;

  out122 <= Logical_Operator_out2170_out1;

  out123 <= Logical_Operator_out2171_out1;

  out124 <= Logical_Operator_out2172_out1;

  out125 <= Logical_Operator_out2173_out1;

  out126 <= Logical_Operator_out2174_out1;

  out127 <= Logical_Operator_out2175_out1;

  out128 <= Logical_Operator_out2176_out1;

  out129 <= Logical_Operator_out2177_out1;

  out130 <= Logical_Operator_out2178_out1;

  out131 <= Logical_Operator_out2179_out1;

  out132 <= Logical_Operator_out2180_out1;

  out133 <= Logical_Operator_out2181_out1;

  out134 <= Logical_Operator_out2182_out1;

  out135 <= Logical_Operator_out2183_out1;

  out136 <= Logical_Operator_out2184_out1;

  out137 <= Logical_Operator_out2185_out1;

  out138 <= Logical_Operator_out2186_out1;

  out139 <= Logical_Operator_out2187_out1;

  out140 <= Logical_Operator_out2188_out1;

  out141 <= Logical_Operator_out2189_out1;

  out142 <= Logical_Operator_out2190_out1;

  out143 <= Logical_Operator_out2191_out1;

  out144 <= Logical_Operator_out2192_out1;

  out145 <= Logical_Operator_out2193_out1;

  out146 <= Logical_Operator_out2194_out1;

  out147 <= Logical_Operator_out2195_out1;

  out148 <= Logical_Operator_out2196_out1;

  out149 <= Logical_Operator_out2197_out1;

  out150 <= Logical_Operator_out2198_out1;

  out151 <= Logical_Operator_out2199_out1;

  out152 <= Logical_Operator_out2200_out1;

  out153 <= Logical_Operator_out2201_out1;

  out154 <= Logical_Operator_out2202_out1;

  out155 <= Logical_Operator_out2203_out1;

  out156 <= Logical_Operator_out2204_out1;

  out157 <= Logical_Operator_out2205_out1;

  out158 <= Logical_Operator_out2206_out1;

  out159 <= Logical_Operator_out2207_out1;

  out160 <= Logical_Operator_out2208_out1;

  out161 <= Logical_Operator_out2209_out1;

  out162 <= Logical_Operator_out2210_out1;

  out163 <= Logical_Operator_out2211_out1;

  out164 <= Logical_Operator_out2212_out1;

  out165 <= Logical_Operator_out2213_out1;

  out166 <= Logical_Operator_out2214_out1;

  out167 <= Logical_Operator_out2215_out1;

  out168 <= Logical_Operator_out2216_out1;

  out169 <= Logical_Operator_out2217_out1;

  out170 <= Logical_Operator_out2218_out1;

  out171 <= Logical_Operator_out2219_out1;

  out172 <= Logical_Operator_out2220_out1;

  out173 <= Logical_Operator_out2221_out1;

  out174 <= Logical_Operator_out2222_out1;

  out175 <= Logical_Operator_out2223_out1;

  out176 <= Logical_Operator_out2224_out1;

  out177 <= Logical_Operator_out2225_out1;

  out178 <= Logical_Operator_out2226_out1;

  out179 <= Logical_Operator_out2227_out1;

  out180 <= Logical_Operator_out2228_out1;

  out181 <= Logical_Operator_out2229_out1;

  out182 <= Logical_Operator_out2230_out1;

  out183 <= Logical_Operator_out2231_out1;

  out184 <= Logical_Operator_out2232_out1;

  out185 <= Logical_Operator_out2233_out1;

  out186 <= Logical_Operator_out2234_out1;

  out187 <= Logical_Operator_out2235_out1;

  out188 <= Logical_Operator_out2236_out1;

  out189 <= Logical_Operator_out2237_out1;

  out190 <= Logical_Operator_out2238_out1;

  out191 <= Logical_Operator_out2239_out1;

  out192 <= Logical_Operator_out2240_out1;

  out193 <= Logical_Operator_out2241_out1;

  out194 <= Logical_Operator_out2242_out1;

  out195 <= Logical_Operator_out2243_out1;

  out196 <= Logical_Operator_out2244_out1;

  out197 <= Logical_Operator_out2245_out1;

  out198 <= Logical_Operator_out2246_out1;

  out199 <= Logical_Operator_out2247_out1;

  out200 <= Logical_Operator_out2248_out1;

  out201 <= Logical_Operator_out2249_out1;

  out202 <= Logical_Operator_out2250_out1;

  out203 <= Logical_Operator_out2251_out1;

  out204 <= Logical_Operator_out2252_out1;

  out205 <= Logical_Operator_out2253_out1;

  out206 <= Logical_Operator_out2254_out1;

  out207 <= Logical_Operator_out2255_out1;

  out208 <= Logical_Operator_out2256_out1;

  out209 <= Logical_Operator_out2257_out1;

  out210 <= Logical_Operator_out2258_out1;

  out211 <= Logical_Operator_out2259_out1;

  out212 <= Logical_Operator_out2260_out1;

  out213 <= Logical_Operator_out2261_out1;

  out214 <= Logical_Operator_out2262_out1;

  out215 <= Logical_Operator_out2263_out1;

  out216 <= Logical_Operator_out2264_out1;

  out217 <= Logical_Operator_out2265_out1;

  out218 <= Logical_Operator_out2266_out1;

  out219 <= Logical_Operator_out2267_out1;

  out220 <= Logical_Operator_out2268_out1;

  out221 <= Logical_Operator_out2269_out1;

  out222 <= Logical_Operator_out2270_out1;

  out223 <= Logical_Operator_out2271_out1;

  out224 <= Logical_Operator_out2272_out1;

  out225 <= Logical_Operator_out2273_out1;

  out226 <= Logical_Operator_out2274_out1;

  out227 <= Logical_Operator_out2275_out1;

  out228 <= Logical_Operator_out2276_out1;

  out229 <= Logical_Operator_out2277_out1;

  out230 <= Logical_Operator_out2278_out1;

  out231 <= Logical_Operator_out2279_out1;

  out232 <= Logical_Operator_out2280_out1;

  out233 <= Logical_Operator_out2281_out1;

  out234 <= Logical_Operator_out2282_out1;

  out235 <= Logical_Operator_out2283_out1;

  out236 <= Logical_Operator_out2284_out1;

  out237 <= Logical_Operator_out2285_out1;

  out238 <= Logical_Operator_out2286_out1;

  out239 <= Logical_Operator_out2287_out1;

  out240 <= Logical_Operator_out2288_out1;

  out241 <= Logical_Operator_out2289_out1;

  out242 <= Logical_Operator_out2290_out1;

  out243 <= Logical_Operator_out2291_out1;

  out244 <= Logical_Operator_out2292_out1;

  out245 <= Logical_Operator_out2293_out1;

  out246 <= Logical_Operator_out2294_out1;

  out247 <= Logical_Operator_out2295_out1;

  out248 <= Logical_Operator_out2296_out1;

  out249 <= Logical_Operator_out2297_out1;

  out250 <= Logical_Operator_out2298_out1;

  out251 <= Logical_Operator_out2299_out1;

  out252 <= Logical_Operator_out2300_out1;

  out253 <= Logical_Operator_out2301_out1;

  out254 <= Logical_Operator_out2302_out1;

  out255 <= Logical_Operator_out2303_out1;

  out256 <= Logical_Operator_out2304_out1;

  out257 <= Logical_Operator_out1921_out1;

  out258 <= Logical_Operator_out1922_out1;

  out259 <= Logical_Operator_out1923_out1;

  out260 <= Logical_Operator_out1924_out1;

  out261 <= Logical_Operator_out1925_out1;

  out262 <= Logical_Operator_out1926_out1;

  out263 <= Logical_Operator_out1927_out1;

  out264 <= Logical_Operator_out1928_out1;

  out265 <= Logical_Operator_out1929_out1;

  out266 <= Logical_Operator_out1930_out1;

  out267 <= Logical_Operator_out1931_out1;

  out268 <= Logical_Operator_out1932_out1;

  out269 <= Logical_Operator_out1933_out1;

  out270 <= Logical_Operator_out1934_out1;

  out271 <= Logical_Operator_out1935_out1;

  out272 <= Logical_Operator_out1936_out1;

  out273 <= Logical_Operator_out1937_out1;

  out274 <= Logical_Operator_out1938_out1;

  out275 <= Logical_Operator_out1939_out1;

  out276 <= Logical_Operator_out1940_out1;

  out277 <= Logical_Operator_out1941_out1;

  out278 <= Logical_Operator_out1942_out1;

  out279 <= Logical_Operator_out1943_out1;

  out280 <= Logical_Operator_out1944_out1;

  out281 <= Logical_Operator_out1945_out1;

  out282 <= Logical_Operator_out1946_out1;

  out283 <= Logical_Operator_out1947_out1;

  out284 <= Logical_Operator_out1948_out1;

  out285 <= Logical_Operator_out1949_out1;

  out286 <= Logical_Operator_out1950_out1;

  out287 <= Logical_Operator_out1951_out1;

  out288 <= Logical_Operator_out1952_out1;

  out289 <= Logical_Operator_out1953_out1;

  out290 <= Logical_Operator_out1954_out1;

  out291 <= Logical_Operator_out1955_out1;

  out292 <= Logical_Operator_out1956_out1;

  out293 <= Logical_Operator_out1957_out1;

  out294 <= Logical_Operator_out1958_out1;

  out295 <= Logical_Operator_out1959_out1;

  out296 <= Logical_Operator_out1960_out1;

  out297 <= Logical_Operator_out1961_out1;

  out298 <= Logical_Operator_out1962_out1;

  out299 <= Logical_Operator_out1963_out1;

  out300 <= Logical_Operator_out1964_out1;

  out301 <= Logical_Operator_out1965_out1;

  out302 <= Logical_Operator_out1966_out1;

  out303 <= Logical_Operator_out1967_out1;

  out304 <= Logical_Operator_out1968_out1;

  out305 <= Logical_Operator_out1969_out1;

  out306 <= Logical_Operator_out1970_out1;

  out307 <= Logical_Operator_out1971_out1;

  out308 <= Logical_Operator_out1972_out1;

  out309 <= Logical_Operator_out1973_out1;

  out310 <= Logical_Operator_out1974_out1;

  out311 <= Logical_Operator_out1975_out1;

  out312 <= Logical_Operator_out1976_out1;

  out313 <= Logical_Operator_out1977_out1;

  out314 <= Logical_Operator_out1978_out1;

  out315 <= Logical_Operator_out1979_out1;

  out316 <= Logical_Operator_out1980_out1;

  out317 <= Logical_Operator_out1981_out1;

  out318 <= Logical_Operator_out1982_out1;

  out319 <= Logical_Operator_out1983_out1;

  out320 <= Logical_Operator_out1984_out1;

  out321 <= Logical_Operator_out1985_out1;

  out322 <= Logical_Operator_out1986_out1;

  out323 <= Logical_Operator_out1987_out1;

  out324 <= Logical_Operator_out1988_out1;

  out325 <= Logical_Operator_out1989_out1;

  out326 <= Logical_Operator_out1990_out1;

  out327 <= Logical_Operator_out1991_out1;

  out328 <= Logical_Operator_out1992_out1;

  out329 <= Logical_Operator_out1993_out1;

  out330 <= Logical_Operator_out1994_out1;

  out331 <= Logical_Operator_out1995_out1;

  out332 <= Logical_Operator_out1996_out1;

  out333 <= Logical_Operator_out1997_out1;

  out334 <= Logical_Operator_out1998_out1;

  out335 <= Logical_Operator_out1999_out1;

  out336 <= Logical_Operator_out2000_out1;

  out337 <= Logical_Operator_out2001_out1;

  out338 <= Logical_Operator_out2002_out1;

  out339 <= Logical_Operator_out2003_out1;

  out340 <= Logical_Operator_out2004_out1;

  out341 <= Logical_Operator_out2005_out1;

  out342 <= Logical_Operator_out2006_out1;

  out343 <= Logical_Operator_out2007_out1;

  out344 <= Logical_Operator_out2008_out1;

  out345 <= Logical_Operator_out2009_out1;

  out346 <= Logical_Operator_out2010_out1;

  out347 <= Logical_Operator_out2011_out1;

  out348 <= Logical_Operator_out2012_out1;

  out349 <= Logical_Operator_out2013_out1;

  out350 <= Logical_Operator_out2014_out1;

  out351 <= Logical_Operator_out2015_out1;

  out352 <= Logical_Operator_out2016_out1;

  out353 <= Logical_Operator_out2017_out1;

  out354 <= Logical_Operator_out2018_out1;

  out355 <= Logical_Operator_out2019_out1;

  out356 <= Logical_Operator_out2020_out1;

  out357 <= Logical_Operator_out2021_out1;

  out358 <= Logical_Operator_out2022_out1;

  out359 <= Logical_Operator_out2023_out1;

  out360 <= Logical_Operator_out2024_out1;

  out361 <= Logical_Operator_out2025_out1;

  out362 <= Logical_Operator_out2026_out1;

  out363 <= Logical_Operator_out2027_out1;

  out364 <= Logical_Operator_out2028_out1;

  out365 <= Logical_Operator_out2029_out1;

  out366 <= Logical_Operator_out2030_out1;

  out367 <= Logical_Operator_out2031_out1;

  out368 <= Logical_Operator_out2032_out1;

  out369 <= Logical_Operator_out2033_out1;

  out370 <= Logical_Operator_out2034_out1;

  out371 <= Logical_Operator_out2035_out1;

  out372 <= Logical_Operator_out2036_out1;

  out373 <= Logical_Operator_out2037_out1;

  out374 <= Logical_Operator_out2038_out1;

  out375 <= Logical_Operator_out2039_out1;

  out376 <= Logical_Operator_out2040_out1;

  out377 <= Logical_Operator_out2041_out1;

  out378 <= Logical_Operator_out2042_out1;

  out379 <= Logical_Operator_out2043_out1;

  out380 <= Logical_Operator_out2044_out1;

  out381 <= Logical_Operator_out2045_out1;

  out382 <= Logical_Operator_out2046_out1;

  out383 <= Logical_Operator_out2047_out1;

  out384 <= Logical_Operator_out2048_out1;

  out385 <= Logical_Operator_out1729_out1;

  out386 <= Logical_Operator_out1730_out1;

  out387 <= Logical_Operator_out1731_out1;

  out388 <= Logical_Operator_out1732_out1;

  out389 <= Logical_Operator_out1733_out1;

  out390 <= Logical_Operator_out1734_out1;

  out391 <= Logical_Operator_out1735_out1;

  out392 <= Logical_Operator_out1736_out1;

  out393 <= Logical_Operator_out1737_out1;

  out394 <= Logical_Operator_out1738_out1;

  out395 <= Logical_Operator_out1739_out1;

  out396 <= Logical_Operator_out1740_out1;

  out397 <= Logical_Operator_out1741_out1;

  out398 <= Logical_Operator_out1742_out1;

  out399 <= Logical_Operator_out1743_out1;

  out400 <= Logical_Operator_out1744_out1;

  out401 <= Logical_Operator_out1745_out1;

  out402 <= Logical_Operator_out1746_out1;

  out403 <= Logical_Operator_out1747_out1;

  out404 <= Logical_Operator_out1748_out1;

  out405 <= Logical_Operator_out1749_out1;

  out406 <= Logical_Operator_out1750_out1;

  out407 <= Logical_Operator_out1751_out1;

  out408 <= Logical_Operator_out1752_out1;

  out409 <= Logical_Operator_out1753_out1;

  out410 <= Logical_Operator_out1754_out1;

  out411 <= Logical_Operator_out1755_out1;

  out412 <= Logical_Operator_out1756_out1;

  out413 <= Logical_Operator_out1757_out1;

  out414 <= Logical_Operator_out1758_out1;

  out415 <= Logical_Operator_out1759_out1;

  out416 <= Logical_Operator_out1760_out1;

  out417 <= Logical_Operator_out1761_out1;

  out418 <= Logical_Operator_out1762_out1;

  out419 <= Logical_Operator_out1763_out1;

  out420 <= Logical_Operator_out1764_out1;

  out421 <= Logical_Operator_out1765_out1;

  out422 <= Logical_Operator_out1766_out1;

  out423 <= Logical_Operator_out1767_out1;

  out424 <= Logical_Operator_out1768_out1;

  out425 <= Logical_Operator_out1769_out1;

  out426 <= Logical_Operator_out1770_out1;

  out427 <= Logical_Operator_out1771_out1;

  out428 <= Logical_Operator_out1772_out1;

  out429 <= Logical_Operator_out1773_out1;

  out430 <= Logical_Operator_out1774_out1;

  out431 <= Logical_Operator_out1775_out1;

  out432 <= Logical_Operator_out1776_out1;

  out433 <= Logical_Operator_out1777_out1;

  out434 <= Logical_Operator_out1778_out1;

  out435 <= Logical_Operator_out1779_out1;

  out436 <= Logical_Operator_out1780_out1;

  out437 <= Logical_Operator_out1781_out1;

  out438 <= Logical_Operator_out1782_out1;

  out439 <= Logical_Operator_out1783_out1;

  out440 <= Logical_Operator_out1784_out1;

  out441 <= Logical_Operator_out1785_out1;

  out442 <= Logical_Operator_out1786_out1;

  out443 <= Logical_Operator_out1787_out1;

  out444 <= Logical_Operator_out1788_out1;

  out445 <= Logical_Operator_out1789_out1;

  out446 <= Logical_Operator_out1790_out1;

  out447 <= Logical_Operator_out1791_out1;

  out448 <= Logical_Operator_out1792_out1;

  out449 <= Logical_Operator_out1505_out1;

  out450 <= Logical_Operator_out1506_out1;

  out451 <= Logical_Operator_out1507_out1;

  out452 <= Logical_Operator_out1508_out1;

  out453 <= Logical_Operator_out1509_out1;

  out454 <= Logical_Operator_out1510_out1;

  out455 <= Logical_Operator_out1511_out1;

  out456 <= Logical_Operator_out1512_out1;

  out457 <= Logical_Operator_out1513_out1;

  out458 <= Logical_Operator_out1514_out1;

  out459 <= Logical_Operator_out1515_out1;

  out460 <= Logical_Operator_out1516_out1;

  out461 <= Logical_Operator_out1517_out1;

  out462 <= Logical_Operator_out1518_out1;

  out463 <= Logical_Operator_out1519_out1;

  out464 <= Logical_Operator_out1520_out1;

  out465 <= Logical_Operator_out1521_out1;

  out466 <= Logical_Operator_out1522_out1;

  out467 <= Logical_Operator_out1523_out1;

  out468 <= Logical_Operator_out1524_out1;

  out469 <= Logical_Operator_out1525_out1;

  out470 <= Logical_Operator_out1526_out1;

  out471 <= Logical_Operator_out1527_out1;

  out472 <= Logical_Operator_out1528_out1;

  out473 <= Logical_Operator_out1529_out1;

  out474 <= Logical_Operator_out1530_out1;

  out475 <= Logical_Operator_out1531_out1;

  out476 <= Logical_Operator_out1532_out1;

  out477 <= Logical_Operator_out1533_out1;

  out478 <= Logical_Operator_out1534_out1;

  out479 <= Logical_Operator_out1535_out1;

  out480 <= Logical_Operator_out1536_out1;

  out481 <= Logical_Operator_out1265_out1;

  out482 <= Logical_Operator_out1266_out1;

  out483 <= Logical_Operator_out1267_out1;

  out484 <= Logical_Operator_out1268_out1;

  out485 <= Logical_Operator_out1269_out1;

  out486 <= Logical_Operator_out1270_out1;

  out487 <= Logical_Operator_out1271_out1;

  out488 <= Logical_Operator_out1272_out1;

  out489 <= Logical_Operator_out1273_out1;

  out490 <= Logical_Operator_out1274_out1;

  out491 <= Logical_Operator_out1275_out1;

  out492 <= Logical_Operator_out1276_out1;

  out493 <= Logical_Operator_out1277_out1;

  out494 <= Logical_Operator_out1278_out1;

  out495 <= Logical_Operator_out1279_out1;

  out496 <= Logical_Operator_out1280_out1;

  out497 <= Logical_Operator_out1017_out1;

  out498 <= Logical_Operator_out1018_out1;

  out499 <= Logical_Operator_out1019_out1;

  out500 <= Logical_Operator_out1020_out1;

  out501 <= Logical_Operator_out1021_out1;

  out502 <= Logical_Operator_out1022_out1;

  out503 <= Logical_Operator_out1023_out1;

  out504 <= Logical_Operator_out1024_out1;

  out505 <= Logical_Operator_out765_out1;

  out506 <= Logical_Operator_out766_out1;

  out507 <= Logical_Operator_out767_out1;

  out508 <= Logical_Operator_out768_out1;

  out509 <= Logical_Operator_out511_out1;

  out510 <= Logical_Operator_out512_out1;

  out511 <= Logical_Operator_out256_out1;

  out512 <= in512;

END rtl;
