LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY encoderN1024 IS
PORT( 
	in1                               :   IN    std_logic;
	in2                               :   IN    std_logic;
	in3                               :   IN    std_logic;
	in4                               :   IN    std_logic;
	in5                               :   IN    std_logic;
	in6                               :   IN    std_logic;
	in7                               :   IN    std_logic;
	in8                               :   IN    std_logic;
	in9                               :   IN    std_logic;
	in10                               :   IN    std_logic;
	in11                               :   IN    std_logic;
	in12                               :   IN    std_logic;
	in13                               :   IN    std_logic;
	in14                               :   IN    std_logic;
	in15                               :   IN    std_logic;
	in16                               :   IN    std_logic;
	in17                               :   IN    std_logic;
	in18                               :   IN    std_logic;
	in19                               :   IN    std_logic;
	in20                               :   IN    std_logic;
	in21                               :   IN    std_logic;
	in22                               :   IN    std_logic;
	in23                               :   IN    std_logic;
	in24                               :   IN    std_logic;
	in25                               :   IN    std_logic;
	in26                               :   IN    std_logic;
	in27                               :   IN    std_logic;
	in28                               :   IN    std_logic;
	in29                               :   IN    std_logic;
	in30                               :   IN    std_logic;
	in31                               :   IN    std_logic;
	in32                               :   IN    std_logic;
	in33                               :   IN    std_logic;
	in34                               :   IN    std_logic;
	in35                               :   IN    std_logic;
	in36                               :   IN    std_logic;
	in37                               :   IN    std_logic;
	in38                               :   IN    std_logic;
	in39                               :   IN    std_logic;
	in40                               :   IN    std_logic;
	in41                               :   IN    std_logic;
	in42                               :   IN    std_logic;
	in43                               :   IN    std_logic;
	in44                               :   IN    std_logic;
	in45                               :   IN    std_logic;
	in46                               :   IN    std_logic;
	in47                               :   IN    std_logic;
	in48                               :   IN    std_logic;
	in49                               :   IN    std_logic;
	in50                               :   IN    std_logic;
	in51                               :   IN    std_logic;
	in52                               :   IN    std_logic;
	in53                               :   IN    std_logic;
	in54                               :   IN    std_logic;
	in55                               :   IN    std_logic;
	in56                               :   IN    std_logic;
	in57                               :   IN    std_logic;
	in58                               :   IN    std_logic;
	in59                               :   IN    std_logic;
	in60                               :   IN    std_logic;
	in61                               :   IN    std_logic;
	in62                               :   IN    std_logic;
	in63                               :   IN    std_logic;
	in64                               :   IN    std_logic;
	in65                               :   IN    std_logic;
	in66                               :   IN    std_logic;
	in67                               :   IN    std_logic;
	in68                               :   IN    std_logic;
	in69                               :   IN    std_logic;
	in70                               :   IN    std_logic;
	in71                               :   IN    std_logic;
	in72                               :   IN    std_logic;
	in73                               :   IN    std_logic;
	in74                               :   IN    std_logic;
	in75                               :   IN    std_logic;
	in76                               :   IN    std_logic;
	in77                               :   IN    std_logic;
	in78                               :   IN    std_logic;
	in79                               :   IN    std_logic;
	in80                               :   IN    std_logic;
	in81                               :   IN    std_logic;
	in82                               :   IN    std_logic;
	in83                               :   IN    std_logic;
	in84                               :   IN    std_logic;
	in85                               :   IN    std_logic;
	in86                               :   IN    std_logic;
	in87                               :   IN    std_logic;
	in88                               :   IN    std_logic;
	in89                               :   IN    std_logic;
	in90                               :   IN    std_logic;
	in91                               :   IN    std_logic;
	in92                               :   IN    std_logic;
	in93                               :   IN    std_logic;
	in94                               :   IN    std_logic;
	in95                               :   IN    std_logic;
	in96                               :   IN    std_logic;
	in97                               :   IN    std_logic;
	in98                               :   IN    std_logic;
	in99                               :   IN    std_logic;
	in100                               :   IN    std_logic;
	in101                               :   IN    std_logic;
	in102                               :   IN    std_logic;
	in103                               :   IN    std_logic;
	in104                               :   IN    std_logic;
	in105                               :   IN    std_logic;
	in106                               :   IN    std_logic;
	in107                               :   IN    std_logic;
	in108                               :   IN    std_logic;
	in109                               :   IN    std_logic;
	in110                               :   IN    std_logic;
	in111                               :   IN    std_logic;
	in112                               :   IN    std_logic;
	in113                               :   IN    std_logic;
	in114                               :   IN    std_logic;
	in115                               :   IN    std_logic;
	in116                               :   IN    std_logic;
	in117                               :   IN    std_logic;
	in118                               :   IN    std_logic;
	in119                               :   IN    std_logic;
	in120                               :   IN    std_logic;
	in121                               :   IN    std_logic;
	in122                               :   IN    std_logic;
	in123                               :   IN    std_logic;
	in124                               :   IN    std_logic;
	in125                               :   IN    std_logic;
	in126                               :   IN    std_logic;
	in127                               :   IN    std_logic;
	in128                               :   IN    std_logic;
	in129                               :   IN    std_logic;
	in130                               :   IN    std_logic;
	in131                               :   IN    std_logic;
	in132                               :   IN    std_logic;
	in133                               :   IN    std_logic;
	in134                               :   IN    std_logic;
	in135                               :   IN    std_logic;
	in136                               :   IN    std_logic;
	in137                               :   IN    std_logic;
	in138                               :   IN    std_logic;
	in139                               :   IN    std_logic;
	in140                               :   IN    std_logic;
	in141                               :   IN    std_logic;
	in142                               :   IN    std_logic;
	in143                               :   IN    std_logic;
	in144                               :   IN    std_logic;
	in145                               :   IN    std_logic;
	in146                               :   IN    std_logic;
	in147                               :   IN    std_logic;
	in148                               :   IN    std_logic;
	in149                               :   IN    std_logic;
	in150                               :   IN    std_logic;
	in151                               :   IN    std_logic;
	in152                               :   IN    std_logic;
	in153                               :   IN    std_logic;
	in154                               :   IN    std_logic;
	in155                               :   IN    std_logic;
	in156                               :   IN    std_logic;
	in157                               :   IN    std_logic;
	in158                               :   IN    std_logic;
	in159                               :   IN    std_logic;
	in160                               :   IN    std_logic;
	in161                               :   IN    std_logic;
	in162                               :   IN    std_logic;
	in163                               :   IN    std_logic;
	in164                               :   IN    std_logic;
	in165                               :   IN    std_logic;
	in166                               :   IN    std_logic;
	in167                               :   IN    std_logic;
	in168                               :   IN    std_logic;
	in169                               :   IN    std_logic;
	in170                               :   IN    std_logic;
	in171                               :   IN    std_logic;
	in172                               :   IN    std_logic;
	in173                               :   IN    std_logic;
	in174                               :   IN    std_logic;
	in175                               :   IN    std_logic;
	in176                               :   IN    std_logic;
	in177                               :   IN    std_logic;
	in178                               :   IN    std_logic;
	in179                               :   IN    std_logic;
	in180                               :   IN    std_logic;
	in181                               :   IN    std_logic;
	in182                               :   IN    std_logic;
	in183                               :   IN    std_logic;
	in184                               :   IN    std_logic;
	in185                               :   IN    std_logic;
	in186                               :   IN    std_logic;
	in187                               :   IN    std_logic;
	in188                               :   IN    std_logic;
	in189                               :   IN    std_logic;
	in190                               :   IN    std_logic;
	in191                               :   IN    std_logic;
	in192                               :   IN    std_logic;
	in193                               :   IN    std_logic;
	in194                               :   IN    std_logic;
	in195                               :   IN    std_logic;
	in196                               :   IN    std_logic;
	in197                               :   IN    std_logic;
	in198                               :   IN    std_logic;
	in199                               :   IN    std_logic;
	in200                               :   IN    std_logic;
	in201                               :   IN    std_logic;
	in202                               :   IN    std_logic;
	in203                               :   IN    std_logic;
	in204                               :   IN    std_logic;
	in205                               :   IN    std_logic;
	in206                               :   IN    std_logic;
	in207                               :   IN    std_logic;
	in208                               :   IN    std_logic;
	in209                               :   IN    std_logic;
	in210                               :   IN    std_logic;
	in211                               :   IN    std_logic;
	in212                               :   IN    std_logic;
	in213                               :   IN    std_logic;
	in214                               :   IN    std_logic;
	in215                               :   IN    std_logic;
	in216                               :   IN    std_logic;
	in217                               :   IN    std_logic;
	in218                               :   IN    std_logic;
	in219                               :   IN    std_logic;
	in220                               :   IN    std_logic;
	in221                               :   IN    std_logic;
	in222                               :   IN    std_logic;
	in223                               :   IN    std_logic;
	in224                               :   IN    std_logic;
	in225                               :   IN    std_logic;
	in226                               :   IN    std_logic;
	in227                               :   IN    std_logic;
	in228                               :   IN    std_logic;
	in229                               :   IN    std_logic;
	in230                               :   IN    std_logic;
	in231                               :   IN    std_logic;
	in232                               :   IN    std_logic;
	in233                               :   IN    std_logic;
	in234                               :   IN    std_logic;
	in235                               :   IN    std_logic;
	in236                               :   IN    std_logic;
	in237                               :   IN    std_logic;
	in238                               :   IN    std_logic;
	in239                               :   IN    std_logic;
	in240                               :   IN    std_logic;
	in241                               :   IN    std_logic;
	in242                               :   IN    std_logic;
	in243                               :   IN    std_logic;
	in244                               :   IN    std_logic;
	in245                               :   IN    std_logic;
	in246                               :   IN    std_logic;
	in247                               :   IN    std_logic;
	in248                               :   IN    std_logic;
	in249                               :   IN    std_logic;
	in250                               :   IN    std_logic;
	in251                               :   IN    std_logic;
	in252                               :   IN    std_logic;
	in253                               :   IN    std_logic;
	in254                               :   IN    std_logic;
	in255                               :   IN    std_logic;
	in256                               :   IN    std_logic;
	in257                               :   IN    std_logic;
	in258                               :   IN    std_logic;
	in259                               :   IN    std_logic;
	in260                               :   IN    std_logic;
	in261                               :   IN    std_logic;
	in262                               :   IN    std_logic;
	in263                               :   IN    std_logic;
	in264                               :   IN    std_logic;
	in265                               :   IN    std_logic;
	in266                               :   IN    std_logic;
	in267                               :   IN    std_logic;
	in268                               :   IN    std_logic;
	in269                               :   IN    std_logic;
	in270                               :   IN    std_logic;
	in271                               :   IN    std_logic;
	in272                               :   IN    std_logic;
	in273                               :   IN    std_logic;
	in274                               :   IN    std_logic;
	in275                               :   IN    std_logic;
	in276                               :   IN    std_logic;
	in277                               :   IN    std_logic;
	in278                               :   IN    std_logic;
	in279                               :   IN    std_logic;
	in280                               :   IN    std_logic;
	in281                               :   IN    std_logic;
	in282                               :   IN    std_logic;
	in283                               :   IN    std_logic;
	in284                               :   IN    std_logic;
	in285                               :   IN    std_logic;
	in286                               :   IN    std_logic;
	in287                               :   IN    std_logic;
	in288                               :   IN    std_logic;
	in289                               :   IN    std_logic;
	in290                               :   IN    std_logic;
	in291                               :   IN    std_logic;
	in292                               :   IN    std_logic;
	in293                               :   IN    std_logic;
	in294                               :   IN    std_logic;
	in295                               :   IN    std_logic;
	in296                               :   IN    std_logic;
	in297                               :   IN    std_logic;
	in298                               :   IN    std_logic;
	in299                               :   IN    std_logic;
	in300                               :   IN    std_logic;
	in301                               :   IN    std_logic;
	in302                               :   IN    std_logic;
	in303                               :   IN    std_logic;
	in304                               :   IN    std_logic;
	in305                               :   IN    std_logic;
	in306                               :   IN    std_logic;
	in307                               :   IN    std_logic;
	in308                               :   IN    std_logic;
	in309                               :   IN    std_logic;
	in310                               :   IN    std_logic;
	in311                               :   IN    std_logic;
	in312                               :   IN    std_logic;
	in313                               :   IN    std_logic;
	in314                               :   IN    std_logic;
	in315                               :   IN    std_logic;
	in316                               :   IN    std_logic;
	in317                               :   IN    std_logic;
	in318                               :   IN    std_logic;
	in319                               :   IN    std_logic;
	in320                               :   IN    std_logic;
	in321                               :   IN    std_logic;
	in322                               :   IN    std_logic;
	in323                               :   IN    std_logic;
	in324                               :   IN    std_logic;
	in325                               :   IN    std_logic;
	in326                               :   IN    std_logic;
	in327                               :   IN    std_logic;
	in328                               :   IN    std_logic;
	in329                               :   IN    std_logic;
	in330                               :   IN    std_logic;
	in331                               :   IN    std_logic;
	in332                               :   IN    std_logic;
	in333                               :   IN    std_logic;
	in334                               :   IN    std_logic;
	in335                               :   IN    std_logic;
	in336                               :   IN    std_logic;
	in337                               :   IN    std_logic;
	in338                               :   IN    std_logic;
	in339                               :   IN    std_logic;
	in340                               :   IN    std_logic;
	in341                               :   IN    std_logic;
	in342                               :   IN    std_logic;
	in343                               :   IN    std_logic;
	in344                               :   IN    std_logic;
	in345                               :   IN    std_logic;
	in346                               :   IN    std_logic;
	in347                               :   IN    std_logic;
	in348                               :   IN    std_logic;
	in349                               :   IN    std_logic;
	in350                               :   IN    std_logic;
	in351                               :   IN    std_logic;
	in352                               :   IN    std_logic;
	in353                               :   IN    std_logic;
	in354                               :   IN    std_logic;
	in355                               :   IN    std_logic;
	in356                               :   IN    std_logic;
	in357                               :   IN    std_logic;
	in358                               :   IN    std_logic;
	in359                               :   IN    std_logic;
	in360                               :   IN    std_logic;
	in361                               :   IN    std_logic;
	in362                               :   IN    std_logic;
	in363                               :   IN    std_logic;
	in364                               :   IN    std_logic;
	in365                               :   IN    std_logic;
	in366                               :   IN    std_logic;
	in367                               :   IN    std_logic;
	in368                               :   IN    std_logic;
	in369                               :   IN    std_logic;
	in370                               :   IN    std_logic;
	in371                               :   IN    std_logic;
	in372                               :   IN    std_logic;
	in373                               :   IN    std_logic;
	in374                               :   IN    std_logic;
	in375                               :   IN    std_logic;
	in376                               :   IN    std_logic;
	in377                               :   IN    std_logic;
	in378                               :   IN    std_logic;
	in379                               :   IN    std_logic;
	in380                               :   IN    std_logic;
	in381                               :   IN    std_logic;
	in382                               :   IN    std_logic;
	in383                               :   IN    std_logic;
	in384                               :   IN    std_logic;
	in385                               :   IN    std_logic;
	in386                               :   IN    std_logic;
	in387                               :   IN    std_logic;
	in388                               :   IN    std_logic;
	in389                               :   IN    std_logic;
	in390                               :   IN    std_logic;
	in391                               :   IN    std_logic;
	in392                               :   IN    std_logic;
	in393                               :   IN    std_logic;
	in394                               :   IN    std_logic;
	in395                               :   IN    std_logic;
	in396                               :   IN    std_logic;
	in397                               :   IN    std_logic;
	in398                               :   IN    std_logic;
	in399                               :   IN    std_logic;
	in400                               :   IN    std_logic;
	in401                               :   IN    std_logic;
	in402                               :   IN    std_logic;
	in403                               :   IN    std_logic;
	in404                               :   IN    std_logic;
	in405                               :   IN    std_logic;
	in406                               :   IN    std_logic;
	in407                               :   IN    std_logic;
	in408                               :   IN    std_logic;
	in409                               :   IN    std_logic;
	in410                               :   IN    std_logic;
	in411                               :   IN    std_logic;
	in412                               :   IN    std_logic;
	in413                               :   IN    std_logic;
	in414                               :   IN    std_logic;
	in415                               :   IN    std_logic;
	in416                               :   IN    std_logic;
	in417                               :   IN    std_logic;
	in418                               :   IN    std_logic;
	in419                               :   IN    std_logic;
	in420                               :   IN    std_logic;
	in421                               :   IN    std_logic;
	in422                               :   IN    std_logic;
	in423                               :   IN    std_logic;
	in424                               :   IN    std_logic;
	in425                               :   IN    std_logic;
	in426                               :   IN    std_logic;
	in427                               :   IN    std_logic;
	in428                               :   IN    std_logic;
	in429                               :   IN    std_logic;
	in430                               :   IN    std_logic;
	in431                               :   IN    std_logic;
	in432                               :   IN    std_logic;
	in433                               :   IN    std_logic;
	in434                               :   IN    std_logic;
	in435                               :   IN    std_logic;
	in436                               :   IN    std_logic;
	in437                               :   IN    std_logic;
	in438                               :   IN    std_logic;
	in439                               :   IN    std_logic;
	in440                               :   IN    std_logic;
	in441                               :   IN    std_logic;
	in442                               :   IN    std_logic;
	in443                               :   IN    std_logic;
	in444                               :   IN    std_logic;
	in445                               :   IN    std_logic;
	in446                               :   IN    std_logic;
	in447                               :   IN    std_logic;
	in448                               :   IN    std_logic;
	in449                               :   IN    std_logic;
	in450                               :   IN    std_logic;
	in451                               :   IN    std_logic;
	in452                               :   IN    std_logic;
	in453                               :   IN    std_logic;
	in454                               :   IN    std_logic;
	in455                               :   IN    std_logic;
	in456                               :   IN    std_logic;
	in457                               :   IN    std_logic;
	in458                               :   IN    std_logic;
	in459                               :   IN    std_logic;
	in460                               :   IN    std_logic;
	in461                               :   IN    std_logic;
	in462                               :   IN    std_logic;
	in463                               :   IN    std_logic;
	in464                               :   IN    std_logic;
	in465                               :   IN    std_logic;
	in466                               :   IN    std_logic;
	in467                               :   IN    std_logic;
	in468                               :   IN    std_logic;
	in469                               :   IN    std_logic;
	in470                               :   IN    std_logic;
	in471                               :   IN    std_logic;
	in472                               :   IN    std_logic;
	in473                               :   IN    std_logic;
	in474                               :   IN    std_logic;
	in475                               :   IN    std_logic;
	in476                               :   IN    std_logic;
	in477                               :   IN    std_logic;
	in478                               :   IN    std_logic;
	in479                               :   IN    std_logic;
	in480                               :   IN    std_logic;
	in481                               :   IN    std_logic;
	in482                               :   IN    std_logic;
	in483                               :   IN    std_logic;
	in484                               :   IN    std_logic;
	in485                               :   IN    std_logic;
	in486                               :   IN    std_logic;
	in487                               :   IN    std_logic;
	in488                               :   IN    std_logic;
	in489                               :   IN    std_logic;
	in490                               :   IN    std_logic;
	in491                               :   IN    std_logic;
	in492                               :   IN    std_logic;
	in493                               :   IN    std_logic;
	in494                               :   IN    std_logic;
	in495                               :   IN    std_logic;
	in496                               :   IN    std_logic;
	in497                               :   IN    std_logic;
	in498                               :   IN    std_logic;
	in499                               :   IN    std_logic;
	in500                               :   IN    std_logic;
	in501                               :   IN    std_logic;
	in502                               :   IN    std_logic;
	in503                               :   IN    std_logic;
	in504                               :   IN    std_logic;
	in505                               :   IN    std_logic;
	in506                               :   IN    std_logic;
	in507                               :   IN    std_logic;
	in508                               :   IN    std_logic;
	in509                               :   IN    std_logic;
	in510                               :   IN    std_logic;
	in511                               :   IN    std_logic;
	in512                               :   IN    std_logic;
	in513                               :   IN    std_logic;
	in514                               :   IN    std_logic;
	in515                               :   IN    std_logic;
	in516                               :   IN    std_logic;
	in517                               :   IN    std_logic;
	in518                               :   IN    std_logic;
	in519                               :   IN    std_logic;
	in520                               :   IN    std_logic;
	in521                               :   IN    std_logic;
	in522                               :   IN    std_logic;
	in523                               :   IN    std_logic;
	in524                               :   IN    std_logic;
	in525                               :   IN    std_logic;
	in526                               :   IN    std_logic;
	in527                               :   IN    std_logic;
	in528                               :   IN    std_logic;
	in529                               :   IN    std_logic;
	in530                               :   IN    std_logic;
	in531                               :   IN    std_logic;
	in532                               :   IN    std_logic;
	in533                               :   IN    std_logic;
	in534                               :   IN    std_logic;
	in535                               :   IN    std_logic;
	in536                               :   IN    std_logic;
	in537                               :   IN    std_logic;
	in538                               :   IN    std_logic;
	in539                               :   IN    std_logic;
	in540                               :   IN    std_logic;
	in541                               :   IN    std_logic;
	in542                               :   IN    std_logic;
	in543                               :   IN    std_logic;
	in544                               :   IN    std_logic;
	in545                               :   IN    std_logic;
	in546                               :   IN    std_logic;
	in547                               :   IN    std_logic;
	in548                               :   IN    std_logic;
	in549                               :   IN    std_logic;
	in550                               :   IN    std_logic;
	in551                               :   IN    std_logic;
	in552                               :   IN    std_logic;
	in553                               :   IN    std_logic;
	in554                               :   IN    std_logic;
	in555                               :   IN    std_logic;
	in556                               :   IN    std_logic;
	in557                               :   IN    std_logic;
	in558                               :   IN    std_logic;
	in559                               :   IN    std_logic;
	in560                               :   IN    std_logic;
	in561                               :   IN    std_logic;
	in562                               :   IN    std_logic;
	in563                               :   IN    std_logic;
	in564                               :   IN    std_logic;
	in565                               :   IN    std_logic;
	in566                               :   IN    std_logic;
	in567                               :   IN    std_logic;
	in568                               :   IN    std_logic;
	in569                               :   IN    std_logic;
	in570                               :   IN    std_logic;
	in571                               :   IN    std_logic;
	in572                               :   IN    std_logic;
	in573                               :   IN    std_logic;
	in574                               :   IN    std_logic;
	in575                               :   IN    std_logic;
	in576                               :   IN    std_logic;
	in577                               :   IN    std_logic;
	in578                               :   IN    std_logic;
	in579                               :   IN    std_logic;
	in580                               :   IN    std_logic;
	in581                               :   IN    std_logic;
	in582                               :   IN    std_logic;
	in583                               :   IN    std_logic;
	in584                               :   IN    std_logic;
	in585                               :   IN    std_logic;
	in586                               :   IN    std_logic;
	in587                               :   IN    std_logic;
	in588                               :   IN    std_logic;
	in589                               :   IN    std_logic;
	in590                               :   IN    std_logic;
	in591                               :   IN    std_logic;
	in592                               :   IN    std_logic;
	in593                               :   IN    std_logic;
	in594                               :   IN    std_logic;
	in595                               :   IN    std_logic;
	in596                               :   IN    std_logic;
	in597                               :   IN    std_logic;
	in598                               :   IN    std_logic;
	in599                               :   IN    std_logic;
	in600                               :   IN    std_logic;
	in601                               :   IN    std_logic;
	in602                               :   IN    std_logic;
	in603                               :   IN    std_logic;
	in604                               :   IN    std_logic;
	in605                               :   IN    std_logic;
	in606                               :   IN    std_logic;
	in607                               :   IN    std_logic;
	in608                               :   IN    std_logic;
	in609                               :   IN    std_logic;
	in610                               :   IN    std_logic;
	in611                               :   IN    std_logic;
	in612                               :   IN    std_logic;
	in613                               :   IN    std_logic;
	in614                               :   IN    std_logic;
	in615                               :   IN    std_logic;
	in616                               :   IN    std_logic;
	in617                               :   IN    std_logic;
	in618                               :   IN    std_logic;
	in619                               :   IN    std_logic;
	in620                               :   IN    std_logic;
	in621                               :   IN    std_logic;
	in622                               :   IN    std_logic;
	in623                               :   IN    std_logic;
	in624                               :   IN    std_logic;
	in625                               :   IN    std_logic;
	in626                               :   IN    std_logic;
	in627                               :   IN    std_logic;
	in628                               :   IN    std_logic;
	in629                               :   IN    std_logic;
	in630                               :   IN    std_logic;
	in631                               :   IN    std_logic;
	in632                               :   IN    std_logic;
	in633                               :   IN    std_logic;
	in634                               :   IN    std_logic;
	in635                               :   IN    std_logic;
	in636                               :   IN    std_logic;
	in637                               :   IN    std_logic;
	in638                               :   IN    std_logic;
	in639                               :   IN    std_logic;
	in640                               :   IN    std_logic;
	in641                               :   IN    std_logic;
	in642                               :   IN    std_logic;
	in643                               :   IN    std_logic;
	in644                               :   IN    std_logic;
	in645                               :   IN    std_logic;
	in646                               :   IN    std_logic;
	in647                               :   IN    std_logic;
	in648                               :   IN    std_logic;
	in649                               :   IN    std_logic;
	in650                               :   IN    std_logic;
	in651                               :   IN    std_logic;
	in652                               :   IN    std_logic;
	in653                               :   IN    std_logic;
	in654                               :   IN    std_logic;
	in655                               :   IN    std_logic;
	in656                               :   IN    std_logic;
	in657                               :   IN    std_logic;
	in658                               :   IN    std_logic;
	in659                               :   IN    std_logic;
	in660                               :   IN    std_logic;
	in661                               :   IN    std_logic;
	in662                               :   IN    std_logic;
	in663                               :   IN    std_logic;
	in664                               :   IN    std_logic;
	in665                               :   IN    std_logic;
	in666                               :   IN    std_logic;
	in667                               :   IN    std_logic;
	in668                               :   IN    std_logic;
	in669                               :   IN    std_logic;
	in670                               :   IN    std_logic;
	in671                               :   IN    std_logic;
	in672                               :   IN    std_logic;
	in673                               :   IN    std_logic;
	in674                               :   IN    std_logic;
	in675                               :   IN    std_logic;
	in676                               :   IN    std_logic;
	in677                               :   IN    std_logic;
	in678                               :   IN    std_logic;
	in679                               :   IN    std_logic;
	in680                               :   IN    std_logic;
	in681                               :   IN    std_logic;
	in682                               :   IN    std_logic;
	in683                               :   IN    std_logic;
	in684                               :   IN    std_logic;
	in685                               :   IN    std_logic;
	in686                               :   IN    std_logic;
	in687                               :   IN    std_logic;
	in688                               :   IN    std_logic;
	in689                               :   IN    std_logic;
	in690                               :   IN    std_logic;
	in691                               :   IN    std_logic;
	in692                               :   IN    std_logic;
	in693                               :   IN    std_logic;
	in694                               :   IN    std_logic;
	in695                               :   IN    std_logic;
	in696                               :   IN    std_logic;
	in697                               :   IN    std_logic;
	in698                               :   IN    std_logic;
	in699                               :   IN    std_logic;
	in700                               :   IN    std_logic;
	in701                               :   IN    std_logic;
	in702                               :   IN    std_logic;
	in703                               :   IN    std_logic;
	in704                               :   IN    std_logic;
	in705                               :   IN    std_logic;
	in706                               :   IN    std_logic;
	in707                               :   IN    std_logic;
	in708                               :   IN    std_logic;
	in709                               :   IN    std_logic;
	in710                               :   IN    std_logic;
	in711                               :   IN    std_logic;
	in712                               :   IN    std_logic;
	in713                               :   IN    std_logic;
	in714                               :   IN    std_logic;
	in715                               :   IN    std_logic;
	in716                               :   IN    std_logic;
	in717                               :   IN    std_logic;
	in718                               :   IN    std_logic;
	in719                               :   IN    std_logic;
	in720                               :   IN    std_logic;
	in721                               :   IN    std_logic;
	in722                               :   IN    std_logic;
	in723                               :   IN    std_logic;
	in724                               :   IN    std_logic;
	in725                               :   IN    std_logic;
	in726                               :   IN    std_logic;
	in727                               :   IN    std_logic;
	in728                               :   IN    std_logic;
	in729                               :   IN    std_logic;
	in730                               :   IN    std_logic;
	in731                               :   IN    std_logic;
	in732                               :   IN    std_logic;
	in733                               :   IN    std_logic;
	in734                               :   IN    std_logic;
	in735                               :   IN    std_logic;
	in736                               :   IN    std_logic;
	in737                               :   IN    std_logic;
	in738                               :   IN    std_logic;
	in739                               :   IN    std_logic;
	in740                               :   IN    std_logic;
	in741                               :   IN    std_logic;
	in742                               :   IN    std_logic;
	in743                               :   IN    std_logic;
	in744                               :   IN    std_logic;
	in745                               :   IN    std_logic;
	in746                               :   IN    std_logic;
	in747                               :   IN    std_logic;
	in748                               :   IN    std_logic;
	in749                               :   IN    std_logic;
	in750                               :   IN    std_logic;
	in751                               :   IN    std_logic;
	in752                               :   IN    std_logic;
	in753                               :   IN    std_logic;
	in754                               :   IN    std_logic;
	in755                               :   IN    std_logic;
	in756                               :   IN    std_logic;
	in757                               :   IN    std_logic;
	in758                               :   IN    std_logic;
	in759                               :   IN    std_logic;
	in760                               :   IN    std_logic;
	in761                               :   IN    std_logic;
	in762                               :   IN    std_logic;
	in763                               :   IN    std_logic;
	in764                               :   IN    std_logic;
	in765                               :   IN    std_logic;
	in766                               :   IN    std_logic;
	in767                               :   IN    std_logic;
	in768                               :   IN    std_logic;
	in769                               :   IN    std_logic;
	in770                               :   IN    std_logic;
	in771                               :   IN    std_logic;
	in772                               :   IN    std_logic;
	in773                               :   IN    std_logic;
	in774                               :   IN    std_logic;
	in775                               :   IN    std_logic;
	in776                               :   IN    std_logic;
	in777                               :   IN    std_logic;
	in778                               :   IN    std_logic;
	in779                               :   IN    std_logic;
	in780                               :   IN    std_logic;
	in781                               :   IN    std_logic;
	in782                               :   IN    std_logic;
	in783                               :   IN    std_logic;
	in784                               :   IN    std_logic;
	in785                               :   IN    std_logic;
	in786                               :   IN    std_logic;
	in787                               :   IN    std_logic;
	in788                               :   IN    std_logic;
	in789                               :   IN    std_logic;
	in790                               :   IN    std_logic;
	in791                               :   IN    std_logic;
	in792                               :   IN    std_logic;
	in793                               :   IN    std_logic;
	in794                               :   IN    std_logic;
	in795                               :   IN    std_logic;
	in796                               :   IN    std_logic;
	in797                               :   IN    std_logic;
	in798                               :   IN    std_logic;
	in799                               :   IN    std_logic;
	in800                               :   IN    std_logic;
	in801                               :   IN    std_logic;
	in802                               :   IN    std_logic;
	in803                               :   IN    std_logic;
	in804                               :   IN    std_logic;
	in805                               :   IN    std_logic;
	in806                               :   IN    std_logic;
	in807                               :   IN    std_logic;
	in808                               :   IN    std_logic;
	in809                               :   IN    std_logic;
	in810                               :   IN    std_logic;
	in811                               :   IN    std_logic;
	in812                               :   IN    std_logic;
	in813                               :   IN    std_logic;
	in814                               :   IN    std_logic;
	in815                               :   IN    std_logic;
	in816                               :   IN    std_logic;
	in817                               :   IN    std_logic;
	in818                               :   IN    std_logic;
	in819                               :   IN    std_logic;
	in820                               :   IN    std_logic;
	in821                               :   IN    std_logic;
	in822                               :   IN    std_logic;
	in823                               :   IN    std_logic;
	in824                               :   IN    std_logic;
	in825                               :   IN    std_logic;
	in826                               :   IN    std_logic;
	in827                               :   IN    std_logic;
	in828                               :   IN    std_logic;
	in829                               :   IN    std_logic;
	in830                               :   IN    std_logic;
	in831                               :   IN    std_logic;
	in832                               :   IN    std_logic;
	in833                               :   IN    std_logic;
	in834                               :   IN    std_logic;
	in835                               :   IN    std_logic;
	in836                               :   IN    std_logic;
	in837                               :   IN    std_logic;
	in838                               :   IN    std_logic;
	in839                               :   IN    std_logic;
	in840                               :   IN    std_logic;
	in841                               :   IN    std_logic;
	in842                               :   IN    std_logic;
	in843                               :   IN    std_logic;
	in844                               :   IN    std_logic;
	in845                               :   IN    std_logic;
	in846                               :   IN    std_logic;
	in847                               :   IN    std_logic;
	in848                               :   IN    std_logic;
	in849                               :   IN    std_logic;
	in850                               :   IN    std_logic;
	in851                               :   IN    std_logic;
	in852                               :   IN    std_logic;
	in853                               :   IN    std_logic;
	in854                               :   IN    std_logic;
	in855                               :   IN    std_logic;
	in856                               :   IN    std_logic;
	in857                               :   IN    std_logic;
	in858                               :   IN    std_logic;
	in859                               :   IN    std_logic;
	in860                               :   IN    std_logic;
	in861                               :   IN    std_logic;
	in862                               :   IN    std_logic;
	in863                               :   IN    std_logic;
	in864                               :   IN    std_logic;
	in865                               :   IN    std_logic;
	in866                               :   IN    std_logic;
	in867                               :   IN    std_logic;
	in868                               :   IN    std_logic;
	in869                               :   IN    std_logic;
	in870                               :   IN    std_logic;
	in871                               :   IN    std_logic;
	in872                               :   IN    std_logic;
	in873                               :   IN    std_logic;
	in874                               :   IN    std_logic;
	in875                               :   IN    std_logic;
	in876                               :   IN    std_logic;
	in877                               :   IN    std_logic;
	in878                               :   IN    std_logic;
	in879                               :   IN    std_logic;
	in880                               :   IN    std_logic;
	in881                               :   IN    std_logic;
	in882                               :   IN    std_logic;
	in883                               :   IN    std_logic;
	in884                               :   IN    std_logic;
	in885                               :   IN    std_logic;
	in886                               :   IN    std_logic;
	in887                               :   IN    std_logic;
	in888                               :   IN    std_logic;
	in889                               :   IN    std_logic;
	in890                               :   IN    std_logic;
	in891                               :   IN    std_logic;
	in892                               :   IN    std_logic;
	in893                               :   IN    std_logic;
	in894                               :   IN    std_logic;
	in895                               :   IN    std_logic;
	in896                               :   IN    std_logic;
	in897                               :   IN    std_logic;
	in898                               :   IN    std_logic;
	in899                               :   IN    std_logic;
	in900                               :   IN    std_logic;
	in901                               :   IN    std_logic;
	in902                               :   IN    std_logic;
	in903                               :   IN    std_logic;
	in904                               :   IN    std_logic;
	in905                               :   IN    std_logic;
	in906                               :   IN    std_logic;
	in907                               :   IN    std_logic;
	in908                               :   IN    std_logic;
	in909                               :   IN    std_logic;
	in910                               :   IN    std_logic;
	in911                               :   IN    std_logic;
	in912                               :   IN    std_logic;
	in913                               :   IN    std_logic;
	in914                               :   IN    std_logic;
	in915                               :   IN    std_logic;
	in916                               :   IN    std_logic;
	in917                               :   IN    std_logic;
	in918                               :   IN    std_logic;
	in919                               :   IN    std_logic;
	in920                               :   IN    std_logic;
	in921                               :   IN    std_logic;
	in922                               :   IN    std_logic;
	in923                               :   IN    std_logic;
	in924                               :   IN    std_logic;
	in925                               :   IN    std_logic;
	in926                               :   IN    std_logic;
	in927                               :   IN    std_logic;
	in928                               :   IN    std_logic;
	in929                               :   IN    std_logic;
	in930                               :   IN    std_logic;
	in931                               :   IN    std_logic;
	in932                               :   IN    std_logic;
	in933                               :   IN    std_logic;
	in934                               :   IN    std_logic;
	in935                               :   IN    std_logic;
	in936                               :   IN    std_logic;
	in937                               :   IN    std_logic;
	in938                               :   IN    std_logic;
	in939                               :   IN    std_logic;
	in940                               :   IN    std_logic;
	in941                               :   IN    std_logic;
	in942                               :   IN    std_logic;
	in943                               :   IN    std_logic;
	in944                               :   IN    std_logic;
	in945                               :   IN    std_logic;
	in946                               :   IN    std_logic;
	in947                               :   IN    std_logic;
	in948                               :   IN    std_logic;
	in949                               :   IN    std_logic;
	in950                               :   IN    std_logic;
	in951                               :   IN    std_logic;
	in952                               :   IN    std_logic;
	in953                               :   IN    std_logic;
	in954                               :   IN    std_logic;
	in955                               :   IN    std_logic;
	in956                               :   IN    std_logic;
	in957                               :   IN    std_logic;
	in958                               :   IN    std_logic;
	in959                               :   IN    std_logic;
	in960                               :   IN    std_logic;
	in961                               :   IN    std_logic;
	in962                               :   IN    std_logic;
	in963                               :   IN    std_logic;
	in964                               :   IN    std_logic;
	in965                               :   IN    std_logic;
	in966                               :   IN    std_logic;
	in967                               :   IN    std_logic;
	in968                               :   IN    std_logic;
	in969                               :   IN    std_logic;
	in970                               :   IN    std_logic;
	in971                               :   IN    std_logic;
	in972                               :   IN    std_logic;
	in973                               :   IN    std_logic;
	in974                               :   IN    std_logic;
	in975                               :   IN    std_logic;
	in976                               :   IN    std_logic;
	in977                               :   IN    std_logic;
	in978                               :   IN    std_logic;
	in979                               :   IN    std_logic;
	in980                               :   IN    std_logic;
	in981                               :   IN    std_logic;
	in982                               :   IN    std_logic;
	in983                               :   IN    std_logic;
	in984                               :   IN    std_logic;
	in985                               :   IN    std_logic;
	in986                               :   IN    std_logic;
	in987                               :   IN    std_logic;
	in988                               :   IN    std_logic;
	in989                               :   IN    std_logic;
	in990                               :   IN    std_logic;
	in991                               :   IN    std_logic;
	in992                               :   IN    std_logic;
	in993                               :   IN    std_logic;
	in994                               :   IN    std_logic;
	in995                               :   IN    std_logic;
	in996                               :   IN    std_logic;
	in997                               :   IN    std_logic;
	in998                               :   IN    std_logic;
	in999                               :   IN    std_logic;
	in1000                               :   IN    std_logic;
	in1001                               :   IN    std_logic;
	in1002                               :   IN    std_logic;
	in1003                               :   IN    std_logic;
	in1004                               :   IN    std_logic;
	in1005                               :   IN    std_logic;
	in1006                               :   IN    std_logic;
	in1007                               :   IN    std_logic;
	in1008                               :   IN    std_logic;
	in1009                               :   IN    std_logic;
	in1010                               :   IN    std_logic;
	in1011                               :   IN    std_logic;
	in1012                               :   IN    std_logic;
	in1013                               :   IN    std_logic;
	in1014                               :   IN    std_logic;
	in1015                               :   IN    std_logic;
	in1016                               :   IN    std_logic;
	in1017                               :   IN    std_logic;
	in1018                               :   IN    std_logic;
	in1019                               :   IN    std_logic;
	in1020                               :   IN    std_logic;
	in1021                               :   IN    std_logic;
	in1022                               :   IN    std_logic;
	in1023                               :   IN    std_logic;
	in1024                               :   IN    std_logic;
	out1                               :   OUT    std_logic;
	out2                               :   OUT    std_logic;
	out3                               :   OUT    std_logic;
	out4                               :   OUT    std_logic;
	out5                               :   OUT    std_logic;
	out6                               :   OUT    std_logic;
	out7                               :   OUT    std_logic;
	out8                               :   OUT    std_logic;
	out9                               :   OUT    std_logic;
	out10                               :   OUT    std_logic;
	out11                               :   OUT    std_logic;
	out12                               :   OUT    std_logic;
	out13                               :   OUT    std_logic;
	out14                               :   OUT    std_logic;
	out15                               :   OUT    std_logic;
	out16                               :   OUT    std_logic;
	out17                               :   OUT    std_logic;
	out18                               :   OUT    std_logic;
	out19                               :   OUT    std_logic;
	out20                               :   OUT    std_logic;
	out21                               :   OUT    std_logic;
	out22                               :   OUT    std_logic;
	out23                               :   OUT    std_logic;
	out24                               :   OUT    std_logic;
	out25                               :   OUT    std_logic;
	out26                               :   OUT    std_logic;
	out27                               :   OUT    std_logic;
	out28                               :   OUT    std_logic;
	out29                               :   OUT    std_logic;
	out30                               :   OUT    std_logic;
	out31                               :   OUT    std_logic;
	out32                               :   OUT    std_logic;
	out33                               :   OUT    std_logic;
	out34                               :   OUT    std_logic;
	out35                               :   OUT    std_logic;
	out36                               :   OUT    std_logic;
	out37                               :   OUT    std_logic;
	out38                               :   OUT    std_logic;
	out39                               :   OUT    std_logic;
	out40                               :   OUT    std_logic;
	out41                               :   OUT    std_logic;
	out42                               :   OUT    std_logic;
	out43                               :   OUT    std_logic;
	out44                               :   OUT    std_logic;
	out45                               :   OUT    std_logic;
	out46                               :   OUT    std_logic;
	out47                               :   OUT    std_logic;
	out48                               :   OUT    std_logic;
	out49                               :   OUT    std_logic;
	out50                               :   OUT    std_logic;
	out51                               :   OUT    std_logic;
	out52                               :   OUT    std_logic;
	out53                               :   OUT    std_logic;
	out54                               :   OUT    std_logic;
	out55                               :   OUT    std_logic;
	out56                               :   OUT    std_logic;
	out57                               :   OUT    std_logic;
	out58                               :   OUT    std_logic;
	out59                               :   OUT    std_logic;
	out60                               :   OUT    std_logic;
	out61                               :   OUT    std_logic;
	out62                               :   OUT    std_logic;
	out63                               :   OUT    std_logic;
	out64                               :   OUT    std_logic;
	out65                               :   OUT    std_logic;
	out66                               :   OUT    std_logic;
	out67                               :   OUT    std_logic;
	out68                               :   OUT    std_logic;
	out69                               :   OUT    std_logic;
	out70                               :   OUT    std_logic;
	out71                               :   OUT    std_logic;
	out72                               :   OUT    std_logic;
	out73                               :   OUT    std_logic;
	out74                               :   OUT    std_logic;
	out75                               :   OUT    std_logic;
	out76                               :   OUT    std_logic;
	out77                               :   OUT    std_logic;
	out78                               :   OUT    std_logic;
	out79                               :   OUT    std_logic;
	out80                               :   OUT    std_logic;
	out81                               :   OUT    std_logic;
	out82                               :   OUT    std_logic;
	out83                               :   OUT    std_logic;
	out84                               :   OUT    std_logic;
	out85                               :   OUT    std_logic;
	out86                               :   OUT    std_logic;
	out87                               :   OUT    std_logic;
	out88                               :   OUT    std_logic;
	out89                               :   OUT    std_logic;
	out90                               :   OUT    std_logic;
	out91                               :   OUT    std_logic;
	out92                               :   OUT    std_logic;
	out93                               :   OUT    std_logic;
	out94                               :   OUT    std_logic;
	out95                               :   OUT    std_logic;
	out96                               :   OUT    std_logic;
	out97                               :   OUT    std_logic;
	out98                               :   OUT    std_logic;
	out99                               :   OUT    std_logic;
	out100                               :   OUT    std_logic;
	out101                               :   OUT    std_logic;
	out102                               :   OUT    std_logic;
	out103                               :   OUT    std_logic;
	out104                               :   OUT    std_logic;
	out105                               :   OUT    std_logic;
	out106                               :   OUT    std_logic;
	out107                               :   OUT    std_logic;
	out108                               :   OUT    std_logic;
	out109                               :   OUT    std_logic;
	out110                               :   OUT    std_logic;
	out111                               :   OUT    std_logic;
	out112                               :   OUT    std_logic;
	out113                               :   OUT    std_logic;
	out114                               :   OUT    std_logic;
	out115                               :   OUT    std_logic;
	out116                               :   OUT    std_logic;
	out117                               :   OUT    std_logic;
	out118                               :   OUT    std_logic;
	out119                               :   OUT    std_logic;
	out120                               :   OUT    std_logic;
	out121                               :   OUT    std_logic;
	out122                               :   OUT    std_logic;
	out123                               :   OUT    std_logic;
	out124                               :   OUT    std_logic;
	out125                               :   OUT    std_logic;
	out126                               :   OUT    std_logic;
	out127                               :   OUT    std_logic;
	out128                               :   OUT    std_logic;
	out129                               :   OUT    std_logic;
	out130                               :   OUT    std_logic;
	out131                               :   OUT    std_logic;
	out132                               :   OUT    std_logic;
	out133                               :   OUT    std_logic;
	out134                               :   OUT    std_logic;
	out135                               :   OUT    std_logic;
	out136                               :   OUT    std_logic;
	out137                               :   OUT    std_logic;
	out138                               :   OUT    std_logic;
	out139                               :   OUT    std_logic;
	out140                               :   OUT    std_logic;
	out141                               :   OUT    std_logic;
	out142                               :   OUT    std_logic;
	out143                               :   OUT    std_logic;
	out144                               :   OUT    std_logic;
	out145                               :   OUT    std_logic;
	out146                               :   OUT    std_logic;
	out147                               :   OUT    std_logic;
	out148                               :   OUT    std_logic;
	out149                               :   OUT    std_logic;
	out150                               :   OUT    std_logic;
	out151                               :   OUT    std_logic;
	out152                               :   OUT    std_logic;
	out153                               :   OUT    std_logic;
	out154                               :   OUT    std_logic;
	out155                               :   OUT    std_logic;
	out156                               :   OUT    std_logic;
	out157                               :   OUT    std_logic;
	out158                               :   OUT    std_logic;
	out159                               :   OUT    std_logic;
	out160                               :   OUT    std_logic;
	out161                               :   OUT    std_logic;
	out162                               :   OUT    std_logic;
	out163                               :   OUT    std_logic;
	out164                               :   OUT    std_logic;
	out165                               :   OUT    std_logic;
	out166                               :   OUT    std_logic;
	out167                               :   OUT    std_logic;
	out168                               :   OUT    std_logic;
	out169                               :   OUT    std_logic;
	out170                               :   OUT    std_logic;
	out171                               :   OUT    std_logic;
	out172                               :   OUT    std_logic;
	out173                               :   OUT    std_logic;
	out174                               :   OUT    std_logic;
	out175                               :   OUT    std_logic;
	out176                               :   OUT    std_logic;
	out177                               :   OUT    std_logic;
	out178                               :   OUT    std_logic;
	out179                               :   OUT    std_logic;
	out180                               :   OUT    std_logic;
	out181                               :   OUT    std_logic;
	out182                               :   OUT    std_logic;
	out183                               :   OUT    std_logic;
	out184                               :   OUT    std_logic;
	out185                               :   OUT    std_logic;
	out186                               :   OUT    std_logic;
	out187                               :   OUT    std_logic;
	out188                               :   OUT    std_logic;
	out189                               :   OUT    std_logic;
	out190                               :   OUT    std_logic;
	out191                               :   OUT    std_logic;
	out192                               :   OUT    std_logic;
	out193                               :   OUT    std_logic;
	out194                               :   OUT    std_logic;
	out195                               :   OUT    std_logic;
	out196                               :   OUT    std_logic;
	out197                               :   OUT    std_logic;
	out198                               :   OUT    std_logic;
	out199                               :   OUT    std_logic;
	out200                               :   OUT    std_logic;
	out201                               :   OUT    std_logic;
	out202                               :   OUT    std_logic;
	out203                               :   OUT    std_logic;
	out204                               :   OUT    std_logic;
	out205                               :   OUT    std_logic;
	out206                               :   OUT    std_logic;
	out207                               :   OUT    std_logic;
	out208                               :   OUT    std_logic;
	out209                               :   OUT    std_logic;
	out210                               :   OUT    std_logic;
	out211                               :   OUT    std_logic;
	out212                               :   OUT    std_logic;
	out213                               :   OUT    std_logic;
	out214                               :   OUT    std_logic;
	out215                               :   OUT    std_logic;
	out216                               :   OUT    std_logic;
	out217                               :   OUT    std_logic;
	out218                               :   OUT    std_logic;
	out219                               :   OUT    std_logic;
	out220                               :   OUT    std_logic;
	out221                               :   OUT    std_logic;
	out222                               :   OUT    std_logic;
	out223                               :   OUT    std_logic;
	out224                               :   OUT    std_logic;
	out225                               :   OUT    std_logic;
	out226                               :   OUT    std_logic;
	out227                               :   OUT    std_logic;
	out228                               :   OUT    std_logic;
	out229                               :   OUT    std_logic;
	out230                               :   OUT    std_logic;
	out231                               :   OUT    std_logic;
	out232                               :   OUT    std_logic;
	out233                               :   OUT    std_logic;
	out234                               :   OUT    std_logic;
	out235                               :   OUT    std_logic;
	out236                               :   OUT    std_logic;
	out237                               :   OUT    std_logic;
	out238                               :   OUT    std_logic;
	out239                               :   OUT    std_logic;
	out240                               :   OUT    std_logic;
	out241                               :   OUT    std_logic;
	out242                               :   OUT    std_logic;
	out243                               :   OUT    std_logic;
	out244                               :   OUT    std_logic;
	out245                               :   OUT    std_logic;
	out246                               :   OUT    std_logic;
	out247                               :   OUT    std_logic;
	out248                               :   OUT    std_logic;
	out249                               :   OUT    std_logic;
	out250                               :   OUT    std_logic;
	out251                               :   OUT    std_logic;
	out252                               :   OUT    std_logic;
	out253                               :   OUT    std_logic;
	out254                               :   OUT    std_logic;
	out255                               :   OUT    std_logic;
	out256                               :   OUT    std_logic;
	out257                               :   OUT    std_logic;
	out258                               :   OUT    std_logic;
	out259                               :   OUT    std_logic;
	out260                               :   OUT    std_logic;
	out261                               :   OUT    std_logic;
	out262                               :   OUT    std_logic;
	out263                               :   OUT    std_logic;
	out264                               :   OUT    std_logic;
	out265                               :   OUT    std_logic;
	out266                               :   OUT    std_logic;
	out267                               :   OUT    std_logic;
	out268                               :   OUT    std_logic;
	out269                               :   OUT    std_logic;
	out270                               :   OUT    std_logic;
	out271                               :   OUT    std_logic;
	out272                               :   OUT    std_logic;
	out273                               :   OUT    std_logic;
	out274                               :   OUT    std_logic;
	out275                               :   OUT    std_logic;
	out276                               :   OUT    std_logic;
	out277                               :   OUT    std_logic;
	out278                               :   OUT    std_logic;
	out279                               :   OUT    std_logic;
	out280                               :   OUT    std_logic;
	out281                               :   OUT    std_logic;
	out282                               :   OUT    std_logic;
	out283                               :   OUT    std_logic;
	out284                               :   OUT    std_logic;
	out285                               :   OUT    std_logic;
	out286                               :   OUT    std_logic;
	out287                               :   OUT    std_logic;
	out288                               :   OUT    std_logic;
	out289                               :   OUT    std_logic;
	out290                               :   OUT    std_logic;
	out291                               :   OUT    std_logic;
	out292                               :   OUT    std_logic;
	out293                               :   OUT    std_logic;
	out294                               :   OUT    std_logic;
	out295                               :   OUT    std_logic;
	out296                               :   OUT    std_logic;
	out297                               :   OUT    std_logic;
	out298                               :   OUT    std_logic;
	out299                               :   OUT    std_logic;
	out300                               :   OUT    std_logic;
	out301                               :   OUT    std_logic;
	out302                               :   OUT    std_logic;
	out303                               :   OUT    std_logic;
	out304                               :   OUT    std_logic;
	out305                               :   OUT    std_logic;
	out306                               :   OUT    std_logic;
	out307                               :   OUT    std_logic;
	out308                               :   OUT    std_logic;
	out309                               :   OUT    std_logic;
	out310                               :   OUT    std_logic;
	out311                               :   OUT    std_logic;
	out312                               :   OUT    std_logic;
	out313                               :   OUT    std_logic;
	out314                               :   OUT    std_logic;
	out315                               :   OUT    std_logic;
	out316                               :   OUT    std_logic;
	out317                               :   OUT    std_logic;
	out318                               :   OUT    std_logic;
	out319                               :   OUT    std_logic;
	out320                               :   OUT    std_logic;
	out321                               :   OUT    std_logic;
	out322                               :   OUT    std_logic;
	out323                               :   OUT    std_logic;
	out324                               :   OUT    std_logic;
	out325                               :   OUT    std_logic;
	out326                               :   OUT    std_logic;
	out327                               :   OUT    std_logic;
	out328                               :   OUT    std_logic;
	out329                               :   OUT    std_logic;
	out330                               :   OUT    std_logic;
	out331                               :   OUT    std_logic;
	out332                               :   OUT    std_logic;
	out333                               :   OUT    std_logic;
	out334                               :   OUT    std_logic;
	out335                               :   OUT    std_logic;
	out336                               :   OUT    std_logic;
	out337                               :   OUT    std_logic;
	out338                               :   OUT    std_logic;
	out339                               :   OUT    std_logic;
	out340                               :   OUT    std_logic;
	out341                               :   OUT    std_logic;
	out342                               :   OUT    std_logic;
	out343                               :   OUT    std_logic;
	out344                               :   OUT    std_logic;
	out345                               :   OUT    std_logic;
	out346                               :   OUT    std_logic;
	out347                               :   OUT    std_logic;
	out348                               :   OUT    std_logic;
	out349                               :   OUT    std_logic;
	out350                               :   OUT    std_logic;
	out351                               :   OUT    std_logic;
	out352                               :   OUT    std_logic;
	out353                               :   OUT    std_logic;
	out354                               :   OUT    std_logic;
	out355                               :   OUT    std_logic;
	out356                               :   OUT    std_logic;
	out357                               :   OUT    std_logic;
	out358                               :   OUT    std_logic;
	out359                               :   OUT    std_logic;
	out360                               :   OUT    std_logic;
	out361                               :   OUT    std_logic;
	out362                               :   OUT    std_logic;
	out363                               :   OUT    std_logic;
	out364                               :   OUT    std_logic;
	out365                               :   OUT    std_logic;
	out366                               :   OUT    std_logic;
	out367                               :   OUT    std_logic;
	out368                               :   OUT    std_logic;
	out369                               :   OUT    std_logic;
	out370                               :   OUT    std_logic;
	out371                               :   OUT    std_logic;
	out372                               :   OUT    std_logic;
	out373                               :   OUT    std_logic;
	out374                               :   OUT    std_logic;
	out375                               :   OUT    std_logic;
	out376                               :   OUT    std_logic;
	out377                               :   OUT    std_logic;
	out378                               :   OUT    std_logic;
	out379                               :   OUT    std_logic;
	out380                               :   OUT    std_logic;
	out381                               :   OUT    std_logic;
	out382                               :   OUT    std_logic;
	out383                               :   OUT    std_logic;
	out384                               :   OUT    std_logic;
	out385                               :   OUT    std_logic;
	out386                               :   OUT    std_logic;
	out387                               :   OUT    std_logic;
	out388                               :   OUT    std_logic;
	out389                               :   OUT    std_logic;
	out390                               :   OUT    std_logic;
	out391                               :   OUT    std_logic;
	out392                               :   OUT    std_logic;
	out393                               :   OUT    std_logic;
	out394                               :   OUT    std_logic;
	out395                               :   OUT    std_logic;
	out396                               :   OUT    std_logic;
	out397                               :   OUT    std_logic;
	out398                               :   OUT    std_logic;
	out399                               :   OUT    std_logic;
	out400                               :   OUT    std_logic;
	out401                               :   OUT    std_logic;
	out402                               :   OUT    std_logic;
	out403                               :   OUT    std_logic;
	out404                               :   OUT    std_logic;
	out405                               :   OUT    std_logic;
	out406                               :   OUT    std_logic;
	out407                               :   OUT    std_logic;
	out408                               :   OUT    std_logic;
	out409                               :   OUT    std_logic;
	out410                               :   OUT    std_logic;
	out411                               :   OUT    std_logic;
	out412                               :   OUT    std_logic;
	out413                               :   OUT    std_logic;
	out414                               :   OUT    std_logic;
	out415                               :   OUT    std_logic;
	out416                               :   OUT    std_logic;
	out417                               :   OUT    std_logic;
	out418                               :   OUT    std_logic;
	out419                               :   OUT    std_logic;
	out420                               :   OUT    std_logic;
	out421                               :   OUT    std_logic;
	out422                               :   OUT    std_logic;
	out423                               :   OUT    std_logic;
	out424                               :   OUT    std_logic;
	out425                               :   OUT    std_logic;
	out426                               :   OUT    std_logic;
	out427                               :   OUT    std_logic;
	out428                               :   OUT    std_logic;
	out429                               :   OUT    std_logic;
	out430                               :   OUT    std_logic;
	out431                               :   OUT    std_logic;
	out432                               :   OUT    std_logic;
	out433                               :   OUT    std_logic;
	out434                               :   OUT    std_logic;
	out435                               :   OUT    std_logic;
	out436                               :   OUT    std_logic;
	out437                               :   OUT    std_logic;
	out438                               :   OUT    std_logic;
	out439                               :   OUT    std_logic;
	out440                               :   OUT    std_logic;
	out441                               :   OUT    std_logic;
	out442                               :   OUT    std_logic;
	out443                               :   OUT    std_logic;
	out444                               :   OUT    std_logic;
	out445                               :   OUT    std_logic;
	out446                               :   OUT    std_logic;
	out447                               :   OUT    std_logic;
	out448                               :   OUT    std_logic;
	out449                               :   OUT    std_logic;
	out450                               :   OUT    std_logic;
	out451                               :   OUT    std_logic;
	out452                               :   OUT    std_logic;
	out453                               :   OUT    std_logic;
	out454                               :   OUT    std_logic;
	out455                               :   OUT    std_logic;
	out456                               :   OUT    std_logic;
	out457                               :   OUT    std_logic;
	out458                               :   OUT    std_logic;
	out459                               :   OUT    std_logic;
	out460                               :   OUT    std_logic;
	out461                               :   OUT    std_logic;
	out462                               :   OUT    std_logic;
	out463                               :   OUT    std_logic;
	out464                               :   OUT    std_logic;
	out465                               :   OUT    std_logic;
	out466                               :   OUT    std_logic;
	out467                               :   OUT    std_logic;
	out468                               :   OUT    std_logic;
	out469                               :   OUT    std_logic;
	out470                               :   OUT    std_logic;
	out471                               :   OUT    std_logic;
	out472                               :   OUT    std_logic;
	out473                               :   OUT    std_logic;
	out474                               :   OUT    std_logic;
	out475                               :   OUT    std_logic;
	out476                               :   OUT    std_logic;
	out477                               :   OUT    std_logic;
	out478                               :   OUT    std_logic;
	out479                               :   OUT    std_logic;
	out480                               :   OUT    std_logic;
	out481                               :   OUT    std_logic;
	out482                               :   OUT    std_logic;
	out483                               :   OUT    std_logic;
	out484                               :   OUT    std_logic;
	out485                               :   OUT    std_logic;
	out486                               :   OUT    std_logic;
	out487                               :   OUT    std_logic;
	out488                               :   OUT    std_logic;
	out489                               :   OUT    std_logic;
	out490                               :   OUT    std_logic;
	out491                               :   OUT    std_logic;
	out492                               :   OUT    std_logic;
	out493                               :   OUT    std_logic;
	out494                               :   OUT    std_logic;
	out495                               :   OUT    std_logic;
	out496                               :   OUT    std_logic;
	out497                               :   OUT    std_logic;
	out498                               :   OUT    std_logic;
	out499                               :   OUT    std_logic;
	out500                               :   OUT    std_logic;
	out501                               :   OUT    std_logic;
	out502                               :   OUT    std_logic;
	out503                               :   OUT    std_logic;
	out504                               :   OUT    std_logic;
	out505                               :   OUT    std_logic;
	out506                               :   OUT    std_logic;
	out507                               :   OUT    std_logic;
	out508                               :   OUT    std_logic;
	out509                               :   OUT    std_logic;
	out510                               :   OUT    std_logic;
	out511                               :   OUT    std_logic;
	out512                               :   OUT    std_logic;
	out513                               :   OUT    std_logic;
	out514                               :   OUT    std_logic;
	out515                               :   OUT    std_logic;
	out516                               :   OUT    std_logic;
	out517                               :   OUT    std_logic;
	out518                               :   OUT    std_logic;
	out519                               :   OUT    std_logic;
	out520                               :   OUT    std_logic;
	out521                               :   OUT    std_logic;
	out522                               :   OUT    std_logic;
	out523                               :   OUT    std_logic;
	out524                               :   OUT    std_logic;
	out525                               :   OUT    std_logic;
	out526                               :   OUT    std_logic;
	out527                               :   OUT    std_logic;
	out528                               :   OUT    std_logic;
	out529                               :   OUT    std_logic;
	out530                               :   OUT    std_logic;
	out531                               :   OUT    std_logic;
	out532                               :   OUT    std_logic;
	out533                               :   OUT    std_logic;
	out534                               :   OUT    std_logic;
	out535                               :   OUT    std_logic;
	out536                               :   OUT    std_logic;
	out537                               :   OUT    std_logic;
	out538                               :   OUT    std_logic;
	out539                               :   OUT    std_logic;
	out540                               :   OUT    std_logic;
	out541                               :   OUT    std_logic;
	out542                               :   OUT    std_logic;
	out543                               :   OUT    std_logic;
	out544                               :   OUT    std_logic;
	out545                               :   OUT    std_logic;
	out546                               :   OUT    std_logic;
	out547                               :   OUT    std_logic;
	out548                               :   OUT    std_logic;
	out549                               :   OUT    std_logic;
	out550                               :   OUT    std_logic;
	out551                               :   OUT    std_logic;
	out552                               :   OUT    std_logic;
	out553                               :   OUT    std_logic;
	out554                               :   OUT    std_logic;
	out555                               :   OUT    std_logic;
	out556                               :   OUT    std_logic;
	out557                               :   OUT    std_logic;
	out558                               :   OUT    std_logic;
	out559                               :   OUT    std_logic;
	out560                               :   OUT    std_logic;
	out561                               :   OUT    std_logic;
	out562                               :   OUT    std_logic;
	out563                               :   OUT    std_logic;
	out564                               :   OUT    std_logic;
	out565                               :   OUT    std_logic;
	out566                               :   OUT    std_logic;
	out567                               :   OUT    std_logic;
	out568                               :   OUT    std_logic;
	out569                               :   OUT    std_logic;
	out570                               :   OUT    std_logic;
	out571                               :   OUT    std_logic;
	out572                               :   OUT    std_logic;
	out573                               :   OUT    std_logic;
	out574                               :   OUT    std_logic;
	out575                               :   OUT    std_logic;
	out576                               :   OUT    std_logic;
	out577                               :   OUT    std_logic;
	out578                               :   OUT    std_logic;
	out579                               :   OUT    std_logic;
	out580                               :   OUT    std_logic;
	out581                               :   OUT    std_logic;
	out582                               :   OUT    std_logic;
	out583                               :   OUT    std_logic;
	out584                               :   OUT    std_logic;
	out585                               :   OUT    std_logic;
	out586                               :   OUT    std_logic;
	out587                               :   OUT    std_logic;
	out588                               :   OUT    std_logic;
	out589                               :   OUT    std_logic;
	out590                               :   OUT    std_logic;
	out591                               :   OUT    std_logic;
	out592                               :   OUT    std_logic;
	out593                               :   OUT    std_logic;
	out594                               :   OUT    std_logic;
	out595                               :   OUT    std_logic;
	out596                               :   OUT    std_logic;
	out597                               :   OUT    std_logic;
	out598                               :   OUT    std_logic;
	out599                               :   OUT    std_logic;
	out600                               :   OUT    std_logic;
	out601                               :   OUT    std_logic;
	out602                               :   OUT    std_logic;
	out603                               :   OUT    std_logic;
	out604                               :   OUT    std_logic;
	out605                               :   OUT    std_logic;
	out606                               :   OUT    std_logic;
	out607                               :   OUT    std_logic;
	out608                               :   OUT    std_logic;
	out609                               :   OUT    std_logic;
	out610                               :   OUT    std_logic;
	out611                               :   OUT    std_logic;
	out612                               :   OUT    std_logic;
	out613                               :   OUT    std_logic;
	out614                               :   OUT    std_logic;
	out615                               :   OUT    std_logic;
	out616                               :   OUT    std_logic;
	out617                               :   OUT    std_logic;
	out618                               :   OUT    std_logic;
	out619                               :   OUT    std_logic;
	out620                               :   OUT    std_logic;
	out621                               :   OUT    std_logic;
	out622                               :   OUT    std_logic;
	out623                               :   OUT    std_logic;
	out624                               :   OUT    std_logic;
	out625                               :   OUT    std_logic;
	out626                               :   OUT    std_logic;
	out627                               :   OUT    std_logic;
	out628                               :   OUT    std_logic;
	out629                               :   OUT    std_logic;
	out630                               :   OUT    std_logic;
	out631                               :   OUT    std_logic;
	out632                               :   OUT    std_logic;
	out633                               :   OUT    std_logic;
	out634                               :   OUT    std_logic;
	out635                               :   OUT    std_logic;
	out636                               :   OUT    std_logic;
	out637                               :   OUT    std_logic;
	out638                               :   OUT    std_logic;
	out639                               :   OUT    std_logic;
	out640                               :   OUT    std_logic;
	out641                               :   OUT    std_logic;
	out642                               :   OUT    std_logic;
	out643                               :   OUT    std_logic;
	out644                               :   OUT    std_logic;
	out645                               :   OUT    std_logic;
	out646                               :   OUT    std_logic;
	out647                               :   OUT    std_logic;
	out648                               :   OUT    std_logic;
	out649                               :   OUT    std_logic;
	out650                               :   OUT    std_logic;
	out651                               :   OUT    std_logic;
	out652                               :   OUT    std_logic;
	out653                               :   OUT    std_logic;
	out654                               :   OUT    std_logic;
	out655                               :   OUT    std_logic;
	out656                               :   OUT    std_logic;
	out657                               :   OUT    std_logic;
	out658                               :   OUT    std_logic;
	out659                               :   OUT    std_logic;
	out660                               :   OUT    std_logic;
	out661                               :   OUT    std_logic;
	out662                               :   OUT    std_logic;
	out663                               :   OUT    std_logic;
	out664                               :   OUT    std_logic;
	out665                               :   OUT    std_logic;
	out666                               :   OUT    std_logic;
	out667                               :   OUT    std_logic;
	out668                               :   OUT    std_logic;
	out669                               :   OUT    std_logic;
	out670                               :   OUT    std_logic;
	out671                               :   OUT    std_logic;
	out672                               :   OUT    std_logic;
	out673                               :   OUT    std_logic;
	out674                               :   OUT    std_logic;
	out675                               :   OUT    std_logic;
	out676                               :   OUT    std_logic;
	out677                               :   OUT    std_logic;
	out678                               :   OUT    std_logic;
	out679                               :   OUT    std_logic;
	out680                               :   OUT    std_logic;
	out681                               :   OUT    std_logic;
	out682                               :   OUT    std_logic;
	out683                               :   OUT    std_logic;
	out684                               :   OUT    std_logic;
	out685                               :   OUT    std_logic;
	out686                               :   OUT    std_logic;
	out687                               :   OUT    std_logic;
	out688                               :   OUT    std_logic;
	out689                               :   OUT    std_logic;
	out690                               :   OUT    std_logic;
	out691                               :   OUT    std_logic;
	out692                               :   OUT    std_logic;
	out693                               :   OUT    std_logic;
	out694                               :   OUT    std_logic;
	out695                               :   OUT    std_logic;
	out696                               :   OUT    std_logic;
	out697                               :   OUT    std_logic;
	out698                               :   OUT    std_logic;
	out699                               :   OUT    std_logic;
	out700                               :   OUT    std_logic;
	out701                               :   OUT    std_logic;
	out702                               :   OUT    std_logic;
	out703                               :   OUT    std_logic;
	out704                               :   OUT    std_logic;
	out705                               :   OUT    std_logic;
	out706                               :   OUT    std_logic;
	out707                               :   OUT    std_logic;
	out708                               :   OUT    std_logic;
	out709                               :   OUT    std_logic;
	out710                               :   OUT    std_logic;
	out711                               :   OUT    std_logic;
	out712                               :   OUT    std_logic;
	out713                               :   OUT    std_logic;
	out714                               :   OUT    std_logic;
	out715                               :   OUT    std_logic;
	out716                               :   OUT    std_logic;
	out717                               :   OUT    std_logic;
	out718                               :   OUT    std_logic;
	out719                               :   OUT    std_logic;
	out720                               :   OUT    std_logic;
	out721                               :   OUT    std_logic;
	out722                               :   OUT    std_logic;
	out723                               :   OUT    std_logic;
	out724                               :   OUT    std_logic;
	out725                               :   OUT    std_logic;
	out726                               :   OUT    std_logic;
	out727                               :   OUT    std_logic;
	out728                               :   OUT    std_logic;
	out729                               :   OUT    std_logic;
	out730                               :   OUT    std_logic;
	out731                               :   OUT    std_logic;
	out732                               :   OUT    std_logic;
	out733                               :   OUT    std_logic;
	out734                               :   OUT    std_logic;
	out735                               :   OUT    std_logic;
	out736                               :   OUT    std_logic;
	out737                               :   OUT    std_logic;
	out738                               :   OUT    std_logic;
	out739                               :   OUT    std_logic;
	out740                               :   OUT    std_logic;
	out741                               :   OUT    std_logic;
	out742                               :   OUT    std_logic;
	out743                               :   OUT    std_logic;
	out744                               :   OUT    std_logic;
	out745                               :   OUT    std_logic;
	out746                               :   OUT    std_logic;
	out747                               :   OUT    std_logic;
	out748                               :   OUT    std_logic;
	out749                               :   OUT    std_logic;
	out750                               :   OUT    std_logic;
	out751                               :   OUT    std_logic;
	out752                               :   OUT    std_logic;
	out753                               :   OUT    std_logic;
	out754                               :   OUT    std_logic;
	out755                               :   OUT    std_logic;
	out756                               :   OUT    std_logic;
	out757                               :   OUT    std_logic;
	out758                               :   OUT    std_logic;
	out759                               :   OUT    std_logic;
	out760                               :   OUT    std_logic;
	out761                               :   OUT    std_logic;
	out762                               :   OUT    std_logic;
	out763                               :   OUT    std_logic;
	out764                               :   OUT    std_logic;
	out765                               :   OUT    std_logic;
	out766                               :   OUT    std_logic;
	out767                               :   OUT    std_logic;
	out768                               :   OUT    std_logic;
	out769                               :   OUT    std_logic;
	out770                               :   OUT    std_logic;
	out771                               :   OUT    std_logic;
	out772                               :   OUT    std_logic;
	out773                               :   OUT    std_logic;
	out774                               :   OUT    std_logic;
	out775                               :   OUT    std_logic;
	out776                               :   OUT    std_logic;
	out777                               :   OUT    std_logic;
	out778                               :   OUT    std_logic;
	out779                               :   OUT    std_logic;
	out780                               :   OUT    std_logic;
	out781                               :   OUT    std_logic;
	out782                               :   OUT    std_logic;
	out783                               :   OUT    std_logic;
	out784                               :   OUT    std_logic;
	out785                               :   OUT    std_logic;
	out786                               :   OUT    std_logic;
	out787                               :   OUT    std_logic;
	out788                               :   OUT    std_logic;
	out789                               :   OUT    std_logic;
	out790                               :   OUT    std_logic;
	out791                               :   OUT    std_logic;
	out792                               :   OUT    std_logic;
	out793                               :   OUT    std_logic;
	out794                               :   OUT    std_logic;
	out795                               :   OUT    std_logic;
	out796                               :   OUT    std_logic;
	out797                               :   OUT    std_logic;
	out798                               :   OUT    std_logic;
	out799                               :   OUT    std_logic;
	out800                               :   OUT    std_logic;
	out801                               :   OUT    std_logic;
	out802                               :   OUT    std_logic;
	out803                               :   OUT    std_logic;
	out804                               :   OUT    std_logic;
	out805                               :   OUT    std_logic;
	out806                               :   OUT    std_logic;
	out807                               :   OUT    std_logic;
	out808                               :   OUT    std_logic;
	out809                               :   OUT    std_logic;
	out810                               :   OUT    std_logic;
	out811                               :   OUT    std_logic;
	out812                               :   OUT    std_logic;
	out813                               :   OUT    std_logic;
	out814                               :   OUT    std_logic;
	out815                               :   OUT    std_logic;
	out816                               :   OUT    std_logic;
	out817                               :   OUT    std_logic;
	out818                               :   OUT    std_logic;
	out819                               :   OUT    std_logic;
	out820                               :   OUT    std_logic;
	out821                               :   OUT    std_logic;
	out822                               :   OUT    std_logic;
	out823                               :   OUT    std_logic;
	out824                               :   OUT    std_logic;
	out825                               :   OUT    std_logic;
	out826                               :   OUT    std_logic;
	out827                               :   OUT    std_logic;
	out828                               :   OUT    std_logic;
	out829                               :   OUT    std_logic;
	out830                               :   OUT    std_logic;
	out831                               :   OUT    std_logic;
	out832                               :   OUT    std_logic;
	out833                               :   OUT    std_logic;
	out834                               :   OUT    std_logic;
	out835                               :   OUT    std_logic;
	out836                               :   OUT    std_logic;
	out837                               :   OUT    std_logic;
	out838                               :   OUT    std_logic;
	out839                               :   OUT    std_logic;
	out840                               :   OUT    std_logic;
	out841                               :   OUT    std_logic;
	out842                               :   OUT    std_logic;
	out843                               :   OUT    std_logic;
	out844                               :   OUT    std_logic;
	out845                               :   OUT    std_logic;
	out846                               :   OUT    std_logic;
	out847                               :   OUT    std_logic;
	out848                               :   OUT    std_logic;
	out849                               :   OUT    std_logic;
	out850                               :   OUT    std_logic;
	out851                               :   OUT    std_logic;
	out852                               :   OUT    std_logic;
	out853                               :   OUT    std_logic;
	out854                               :   OUT    std_logic;
	out855                               :   OUT    std_logic;
	out856                               :   OUT    std_logic;
	out857                               :   OUT    std_logic;
	out858                               :   OUT    std_logic;
	out859                               :   OUT    std_logic;
	out860                               :   OUT    std_logic;
	out861                               :   OUT    std_logic;
	out862                               :   OUT    std_logic;
	out863                               :   OUT    std_logic;
	out864                               :   OUT    std_logic;
	out865                               :   OUT    std_logic;
	out866                               :   OUT    std_logic;
	out867                               :   OUT    std_logic;
	out868                               :   OUT    std_logic;
	out869                               :   OUT    std_logic;
	out870                               :   OUT    std_logic;
	out871                               :   OUT    std_logic;
	out872                               :   OUT    std_logic;
	out873                               :   OUT    std_logic;
	out874                               :   OUT    std_logic;
	out875                               :   OUT    std_logic;
	out876                               :   OUT    std_logic;
	out877                               :   OUT    std_logic;
	out878                               :   OUT    std_logic;
	out879                               :   OUT    std_logic;
	out880                               :   OUT    std_logic;
	out881                               :   OUT    std_logic;
	out882                               :   OUT    std_logic;
	out883                               :   OUT    std_logic;
	out884                               :   OUT    std_logic;
	out885                               :   OUT    std_logic;
	out886                               :   OUT    std_logic;
	out887                               :   OUT    std_logic;
	out888                               :   OUT    std_logic;
	out889                               :   OUT    std_logic;
	out890                               :   OUT    std_logic;
	out891                               :   OUT    std_logic;
	out892                               :   OUT    std_logic;
	out893                               :   OUT    std_logic;
	out894                               :   OUT    std_logic;
	out895                               :   OUT    std_logic;
	out896                               :   OUT    std_logic;
	out897                               :   OUT    std_logic;
	out898                               :   OUT    std_logic;
	out899                               :   OUT    std_logic;
	out900                               :   OUT    std_logic;
	out901                               :   OUT    std_logic;
	out902                               :   OUT    std_logic;
	out903                               :   OUT    std_logic;
	out904                               :   OUT    std_logic;
	out905                               :   OUT    std_logic;
	out906                               :   OUT    std_logic;
	out907                               :   OUT    std_logic;
	out908                               :   OUT    std_logic;
	out909                               :   OUT    std_logic;
	out910                               :   OUT    std_logic;
	out911                               :   OUT    std_logic;
	out912                               :   OUT    std_logic;
	out913                               :   OUT    std_logic;
	out914                               :   OUT    std_logic;
	out915                               :   OUT    std_logic;
	out916                               :   OUT    std_logic;
	out917                               :   OUT    std_logic;
	out918                               :   OUT    std_logic;
	out919                               :   OUT    std_logic;
	out920                               :   OUT    std_logic;
	out921                               :   OUT    std_logic;
	out922                               :   OUT    std_logic;
	out923                               :   OUT    std_logic;
	out924                               :   OUT    std_logic;
	out925                               :   OUT    std_logic;
	out926                               :   OUT    std_logic;
	out927                               :   OUT    std_logic;
	out928                               :   OUT    std_logic;
	out929                               :   OUT    std_logic;
	out930                               :   OUT    std_logic;
	out931                               :   OUT    std_logic;
	out932                               :   OUT    std_logic;
	out933                               :   OUT    std_logic;
	out934                               :   OUT    std_logic;
	out935                               :   OUT    std_logic;
	out936                               :   OUT    std_logic;
	out937                               :   OUT    std_logic;
	out938                               :   OUT    std_logic;
	out939                               :   OUT    std_logic;
	out940                               :   OUT    std_logic;
	out941                               :   OUT    std_logic;
	out942                               :   OUT    std_logic;
	out943                               :   OUT    std_logic;
	out944                               :   OUT    std_logic;
	out945                               :   OUT    std_logic;
	out946                               :   OUT    std_logic;
	out947                               :   OUT    std_logic;
	out948                               :   OUT    std_logic;
	out949                               :   OUT    std_logic;
	out950                               :   OUT    std_logic;
	out951                               :   OUT    std_logic;
	out952                               :   OUT    std_logic;
	out953                               :   OUT    std_logic;
	out954                               :   OUT    std_logic;
	out955                               :   OUT    std_logic;
	out956                               :   OUT    std_logic;
	out957                               :   OUT    std_logic;
	out958                               :   OUT    std_logic;
	out959                               :   OUT    std_logic;
	out960                               :   OUT    std_logic;
	out961                               :   OUT    std_logic;
	out962                               :   OUT    std_logic;
	out963                               :   OUT    std_logic;
	out964                               :   OUT    std_logic;
	out965                               :   OUT    std_logic;
	out966                               :   OUT    std_logic;
	out967                               :   OUT    std_logic;
	out968                               :   OUT    std_logic;
	out969                               :   OUT    std_logic;
	out970                               :   OUT    std_logic;
	out971                               :   OUT    std_logic;
	out972                               :   OUT    std_logic;
	out973                               :   OUT    std_logic;
	out974                               :   OUT    std_logic;
	out975                               :   OUT    std_logic;
	out976                               :   OUT    std_logic;
	out977                               :   OUT    std_logic;
	out978                               :   OUT    std_logic;
	out979                               :   OUT    std_logic;
	out980                               :   OUT    std_logic;
	out981                               :   OUT    std_logic;
	out982                               :   OUT    std_logic;
	out983                               :   OUT    std_logic;
	out984                               :   OUT    std_logic;
	out985                               :   OUT    std_logic;
	out986                               :   OUT    std_logic;
	out987                               :   OUT    std_logic;
	out988                               :   OUT    std_logic;
	out989                               :   OUT    std_logic;
	out990                               :   OUT    std_logic;
	out991                               :   OUT    std_logic;
	out992                               :   OUT    std_logic;
	out993                               :   OUT    std_logic;
	out994                               :   OUT    std_logic;
	out995                               :   OUT    std_logic;
	out996                               :   OUT    std_logic;
	out997                               :   OUT    std_logic;
	out998                               :   OUT    std_logic;
	out999                               :   OUT    std_logic;
	out1000                               :   OUT    std_logic;
	out1001                               :   OUT    std_logic;
	out1002                               :   OUT    std_logic;
	out1003                               :   OUT    std_logic;
	out1004                               :   OUT    std_logic;
	out1005                               :   OUT    std_logic;
	out1006                               :   OUT    std_logic;
	out1007                               :   OUT    std_logic;
	out1008                               :   OUT    std_logic;
	out1009                               :   OUT    std_logic;
	out1010                               :   OUT    std_logic;
	out1011                               :   OUT    std_logic;
	out1012                               :   OUT    std_logic;
	out1013                               :   OUT    std_logic;
	out1014                               :   OUT    std_logic;
	out1015                               :   OUT    std_logic;
	out1016                               :   OUT    std_logic;
	out1017                               :   OUT    std_logic;
	out1018                               :   OUT    std_logic;
	out1019                               :   OUT    std_logic;
	out1020                               :   OUT    std_logic;
	out1021                               :   OUT    std_logic;
	out1022                               :   OUT    std_logic;
	out1023                               :   OUT    std_logic;
	out1024                               :   OUT    std_logic
	);
END encoderN1024;

ARCHITECTURE rtl OF encoderN1024 IS

  SIGNAL Logical_Operator_out1_out1            : std_logic;
  SIGNAL Logical_Operator_out2_out1            : std_logic;
  SIGNAL Logical_Operator_out3_out1            : std_logic;
  SIGNAL Logical_Operator_out4_out1            : std_logic;
  SIGNAL Logical_Operator_out5_out1            : std_logic;
  SIGNAL Logical_Operator_out6_out1            : std_logic;
  SIGNAL Logical_Operator_out7_out1            : std_logic;
  SIGNAL Logical_Operator_out8_out1            : std_logic;
  SIGNAL Logical_Operator_out9_out1            : std_logic;
  SIGNAL Logical_Operator_out10_out1            : std_logic;
  SIGNAL Logical_Operator_out11_out1            : std_logic;
  SIGNAL Logical_Operator_out12_out1            : std_logic;
  SIGNAL Logical_Operator_out13_out1            : std_logic;
  SIGNAL Logical_Operator_out14_out1            : std_logic;
  SIGNAL Logical_Operator_out15_out1            : std_logic;
  SIGNAL Logical_Operator_out16_out1            : std_logic;
  SIGNAL Logical_Operator_out17_out1            : std_logic;
  SIGNAL Logical_Operator_out18_out1            : std_logic;
  SIGNAL Logical_Operator_out19_out1            : std_logic;
  SIGNAL Logical_Operator_out20_out1            : std_logic;
  SIGNAL Logical_Operator_out21_out1            : std_logic;
  SIGNAL Logical_Operator_out22_out1            : std_logic;
  SIGNAL Logical_Operator_out23_out1            : std_logic;
  SIGNAL Logical_Operator_out24_out1            : std_logic;
  SIGNAL Logical_Operator_out25_out1            : std_logic;
  SIGNAL Logical_Operator_out26_out1            : std_logic;
  SIGNAL Logical_Operator_out27_out1            : std_logic;
  SIGNAL Logical_Operator_out28_out1            : std_logic;
  SIGNAL Logical_Operator_out29_out1            : std_logic;
  SIGNAL Logical_Operator_out30_out1            : std_logic;
  SIGNAL Logical_Operator_out31_out1            : std_logic;
  SIGNAL Logical_Operator_out32_out1            : std_logic;
  SIGNAL Logical_Operator_out33_out1            : std_logic;
  SIGNAL Logical_Operator_out34_out1            : std_logic;
  SIGNAL Logical_Operator_out35_out1            : std_logic;
  SIGNAL Logical_Operator_out36_out1            : std_logic;
  SIGNAL Logical_Operator_out37_out1            : std_logic;
  SIGNAL Logical_Operator_out38_out1            : std_logic;
  SIGNAL Logical_Operator_out39_out1            : std_logic;
  SIGNAL Logical_Operator_out40_out1            : std_logic;
  SIGNAL Logical_Operator_out41_out1            : std_logic;
  SIGNAL Logical_Operator_out42_out1            : std_logic;
  SIGNAL Logical_Operator_out43_out1            : std_logic;
  SIGNAL Logical_Operator_out44_out1            : std_logic;
  SIGNAL Logical_Operator_out45_out1            : std_logic;
  SIGNAL Logical_Operator_out46_out1            : std_logic;
  SIGNAL Logical_Operator_out47_out1            : std_logic;
  SIGNAL Logical_Operator_out48_out1            : std_logic;
  SIGNAL Logical_Operator_out49_out1            : std_logic;
  SIGNAL Logical_Operator_out50_out1            : std_logic;
  SIGNAL Logical_Operator_out51_out1            : std_logic;
  SIGNAL Logical_Operator_out52_out1            : std_logic;
  SIGNAL Logical_Operator_out53_out1            : std_logic;
  SIGNAL Logical_Operator_out54_out1            : std_logic;
  SIGNAL Logical_Operator_out55_out1            : std_logic;
  SIGNAL Logical_Operator_out56_out1            : std_logic;
  SIGNAL Logical_Operator_out57_out1            : std_logic;
  SIGNAL Logical_Operator_out58_out1            : std_logic;
  SIGNAL Logical_Operator_out59_out1            : std_logic;
  SIGNAL Logical_Operator_out60_out1            : std_logic;
  SIGNAL Logical_Operator_out61_out1            : std_logic;
  SIGNAL Logical_Operator_out62_out1            : std_logic;
  SIGNAL Logical_Operator_out63_out1            : std_logic;
  SIGNAL Logical_Operator_out64_out1            : std_logic;
  SIGNAL Logical_Operator_out65_out1            : std_logic;
  SIGNAL Logical_Operator_out66_out1            : std_logic;
  SIGNAL Logical_Operator_out67_out1            : std_logic;
  SIGNAL Logical_Operator_out68_out1            : std_logic;
  SIGNAL Logical_Operator_out69_out1            : std_logic;
  SIGNAL Logical_Operator_out70_out1            : std_logic;
  SIGNAL Logical_Operator_out71_out1            : std_logic;
  SIGNAL Logical_Operator_out72_out1            : std_logic;
  SIGNAL Logical_Operator_out73_out1            : std_logic;
  SIGNAL Logical_Operator_out74_out1            : std_logic;
  SIGNAL Logical_Operator_out75_out1            : std_logic;
  SIGNAL Logical_Operator_out76_out1            : std_logic;
  SIGNAL Logical_Operator_out77_out1            : std_logic;
  SIGNAL Logical_Operator_out78_out1            : std_logic;
  SIGNAL Logical_Operator_out79_out1            : std_logic;
  SIGNAL Logical_Operator_out80_out1            : std_logic;
  SIGNAL Logical_Operator_out81_out1            : std_logic;
  SIGNAL Logical_Operator_out82_out1            : std_logic;
  SIGNAL Logical_Operator_out83_out1            : std_logic;
  SIGNAL Logical_Operator_out84_out1            : std_logic;
  SIGNAL Logical_Operator_out85_out1            : std_logic;
  SIGNAL Logical_Operator_out86_out1            : std_logic;
  SIGNAL Logical_Operator_out87_out1            : std_logic;
  SIGNAL Logical_Operator_out88_out1            : std_logic;
  SIGNAL Logical_Operator_out89_out1            : std_logic;
  SIGNAL Logical_Operator_out90_out1            : std_logic;
  SIGNAL Logical_Operator_out91_out1            : std_logic;
  SIGNAL Logical_Operator_out92_out1            : std_logic;
  SIGNAL Logical_Operator_out93_out1            : std_logic;
  SIGNAL Logical_Operator_out94_out1            : std_logic;
  SIGNAL Logical_Operator_out95_out1            : std_logic;
  SIGNAL Logical_Operator_out96_out1            : std_logic;
  SIGNAL Logical_Operator_out97_out1            : std_logic;
  SIGNAL Logical_Operator_out98_out1            : std_logic;
  SIGNAL Logical_Operator_out99_out1            : std_logic;
  SIGNAL Logical_Operator_out100_out1            : std_logic;
  SIGNAL Logical_Operator_out101_out1            : std_logic;
  SIGNAL Logical_Operator_out102_out1            : std_logic;
  SIGNAL Logical_Operator_out103_out1            : std_logic;
  SIGNAL Logical_Operator_out104_out1            : std_logic;
  SIGNAL Logical_Operator_out105_out1            : std_logic;
  SIGNAL Logical_Operator_out106_out1            : std_logic;
  SIGNAL Logical_Operator_out107_out1            : std_logic;
  SIGNAL Logical_Operator_out108_out1            : std_logic;
  SIGNAL Logical_Operator_out109_out1            : std_logic;
  SIGNAL Logical_Operator_out110_out1            : std_logic;
  SIGNAL Logical_Operator_out111_out1            : std_logic;
  SIGNAL Logical_Operator_out112_out1            : std_logic;
  SIGNAL Logical_Operator_out113_out1            : std_logic;
  SIGNAL Logical_Operator_out114_out1            : std_logic;
  SIGNAL Logical_Operator_out115_out1            : std_logic;
  SIGNAL Logical_Operator_out116_out1            : std_logic;
  SIGNAL Logical_Operator_out117_out1            : std_logic;
  SIGNAL Logical_Operator_out118_out1            : std_logic;
  SIGNAL Logical_Operator_out119_out1            : std_logic;
  SIGNAL Logical_Operator_out120_out1            : std_logic;
  SIGNAL Logical_Operator_out121_out1            : std_logic;
  SIGNAL Logical_Operator_out122_out1            : std_logic;
  SIGNAL Logical_Operator_out123_out1            : std_logic;
  SIGNAL Logical_Operator_out124_out1            : std_logic;
  SIGNAL Logical_Operator_out125_out1            : std_logic;
  SIGNAL Logical_Operator_out126_out1            : std_logic;
  SIGNAL Logical_Operator_out127_out1            : std_logic;
  SIGNAL Logical_Operator_out128_out1            : std_logic;
  SIGNAL Logical_Operator_out129_out1            : std_logic;
  SIGNAL Logical_Operator_out130_out1            : std_logic;
  SIGNAL Logical_Operator_out131_out1            : std_logic;
  SIGNAL Logical_Operator_out132_out1            : std_logic;
  SIGNAL Logical_Operator_out133_out1            : std_logic;
  SIGNAL Logical_Operator_out134_out1            : std_logic;
  SIGNAL Logical_Operator_out135_out1            : std_logic;
  SIGNAL Logical_Operator_out136_out1            : std_logic;
  SIGNAL Logical_Operator_out137_out1            : std_logic;
  SIGNAL Logical_Operator_out138_out1            : std_logic;
  SIGNAL Logical_Operator_out139_out1            : std_logic;
  SIGNAL Logical_Operator_out140_out1            : std_logic;
  SIGNAL Logical_Operator_out141_out1            : std_logic;
  SIGNAL Logical_Operator_out142_out1            : std_logic;
  SIGNAL Logical_Operator_out143_out1            : std_logic;
  SIGNAL Logical_Operator_out144_out1            : std_logic;
  SIGNAL Logical_Operator_out145_out1            : std_logic;
  SIGNAL Logical_Operator_out146_out1            : std_logic;
  SIGNAL Logical_Operator_out147_out1            : std_logic;
  SIGNAL Logical_Operator_out148_out1            : std_logic;
  SIGNAL Logical_Operator_out149_out1            : std_logic;
  SIGNAL Logical_Operator_out150_out1            : std_logic;
  SIGNAL Logical_Operator_out151_out1            : std_logic;
  SIGNAL Logical_Operator_out152_out1            : std_logic;
  SIGNAL Logical_Operator_out153_out1            : std_logic;
  SIGNAL Logical_Operator_out154_out1            : std_logic;
  SIGNAL Logical_Operator_out155_out1            : std_logic;
  SIGNAL Logical_Operator_out156_out1            : std_logic;
  SIGNAL Logical_Operator_out157_out1            : std_logic;
  SIGNAL Logical_Operator_out158_out1            : std_logic;
  SIGNAL Logical_Operator_out159_out1            : std_logic;
  SIGNAL Logical_Operator_out160_out1            : std_logic;
  SIGNAL Logical_Operator_out161_out1            : std_logic;
  SIGNAL Logical_Operator_out162_out1            : std_logic;
  SIGNAL Logical_Operator_out163_out1            : std_logic;
  SIGNAL Logical_Operator_out164_out1            : std_logic;
  SIGNAL Logical_Operator_out165_out1            : std_logic;
  SIGNAL Logical_Operator_out166_out1            : std_logic;
  SIGNAL Logical_Operator_out167_out1            : std_logic;
  SIGNAL Logical_Operator_out168_out1            : std_logic;
  SIGNAL Logical_Operator_out169_out1            : std_logic;
  SIGNAL Logical_Operator_out170_out1            : std_logic;
  SIGNAL Logical_Operator_out171_out1            : std_logic;
  SIGNAL Logical_Operator_out172_out1            : std_logic;
  SIGNAL Logical_Operator_out173_out1            : std_logic;
  SIGNAL Logical_Operator_out174_out1            : std_logic;
  SIGNAL Logical_Operator_out175_out1            : std_logic;
  SIGNAL Logical_Operator_out176_out1            : std_logic;
  SIGNAL Logical_Operator_out177_out1            : std_logic;
  SIGNAL Logical_Operator_out178_out1            : std_logic;
  SIGNAL Logical_Operator_out179_out1            : std_logic;
  SIGNAL Logical_Operator_out180_out1            : std_logic;
  SIGNAL Logical_Operator_out181_out1            : std_logic;
  SIGNAL Logical_Operator_out182_out1            : std_logic;
  SIGNAL Logical_Operator_out183_out1            : std_logic;
  SIGNAL Logical_Operator_out184_out1            : std_logic;
  SIGNAL Logical_Operator_out185_out1            : std_logic;
  SIGNAL Logical_Operator_out186_out1            : std_logic;
  SIGNAL Logical_Operator_out187_out1            : std_logic;
  SIGNAL Logical_Operator_out188_out1            : std_logic;
  SIGNAL Logical_Operator_out189_out1            : std_logic;
  SIGNAL Logical_Operator_out190_out1            : std_logic;
  SIGNAL Logical_Operator_out191_out1            : std_logic;
  SIGNAL Logical_Operator_out192_out1            : std_logic;
  SIGNAL Logical_Operator_out193_out1            : std_logic;
  SIGNAL Logical_Operator_out194_out1            : std_logic;
  SIGNAL Logical_Operator_out195_out1            : std_logic;
  SIGNAL Logical_Operator_out196_out1            : std_logic;
  SIGNAL Logical_Operator_out197_out1            : std_logic;
  SIGNAL Logical_Operator_out198_out1            : std_logic;
  SIGNAL Logical_Operator_out199_out1            : std_logic;
  SIGNAL Logical_Operator_out200_out1            : std_logic;
  SIGNAL Logical_Operator_out201_out1            : std_logic;
  SIGNAL Logical_Operator_out202_out1            : std_logic;
  SIGNAL Logical_Operator_out203_out1            : std_logic;
  SIGNAL Logical_Operator_out204_out1            : std_logic;
  SIGNAL Logical_Operator_out205_out1            : std_logic;
  SIGNAL Logical_Operator_out206_out1            : std_logic;
  SIGNAL Logical_Operator_out207_out1            : std_logic;
  SIGNAL Logical_Operator_out208_out1            : std_logic;
  SIGNAL Logical_Operator_out209_out1            : std_logic;
  SIGNAL Logical_Operator_out210_out1            : std_logic;
  SIGNAL Logical_Operator_out211_out1            : std_logic;
  SIGNAL Logical_Operator_out212_out1            : std_logic;
  SIGNAL Logical_Operator_out213_out1            : std_logic;
  SIGNAL Logical_Operator_out214_out1            : std_logic;
  SIGNAL Logical_Operator_out215_out1            : std_logic;
  SIGNAL Logical_Operator_out216_out1            : std_logic;
  SIGNAL Logical_Operator_out217_out1            : std_logic;
  SIGNAL Logical_Operator_out218_out1            : std_logic;
  SIGNAL Logical_Operator_out219_out1            : std_logic;
  SIGNAL Logical_Operator_out220_out1            : std_logic;
  SIGNAL Logical_Operator_out221_out1            : std_logic;
  SIGNAL Logical_Operator_out222_out1            : std_logic;
  SIGNAL Logical_Operator_out223_out1            : std_logic;
  SIGNAL Logical_Operator_out224_out1            : std_logic;
  SIGNAL Logical_Operator_out225_out1            : std_logic;
  SIGNAL Logical_Operator_out226_out1            : std_logic;
  SIGNAL Logical_Operator_out227_out1            : std_logic;
  SIGNAL Logical_Operator_out228_out1            : std_logic;
  SIGNAL Logical_Operator_out229_out1            : std_logic;
  SIGNAL Logical_Operator_out230_out1            : std_logic;
  SIGNAL Logical_Operator_out231_out1            : std_logic;
  SIGNAL Logical_Operator_out232_out1            : std_logic;
  SIGNAL Logical_Operator_out233_out1            : std_logic;
  SIGNAL Logical_Operator_out234_out1            : std_logic;
  SIGNAL Logical_Operator_out235_out1            : std_logic;
  SIGNAL Logical_Operator_out236_out1            : std_logic;
  SIGNAL Logical_Operator_out237_out1            : std_logic;
  SIGNAL Logical_Operator_out238_out1            : std_logic;
  SIGNAL Logical_Operator_out239_out1            : std_logic;
  SIGNAL Logical_Operator_out240_out1            : std_logic;
  SIGNAL Logical_Operator_out241_out1            : std_logic;
  SIGNAL Logical_Operator_out242_out1            : std_logic;
  SIGNAL Logical_Operator_out243_out1            : std_logic;
  SIGNAL Logical_Operator_out244_out1            : std_logic;
  SIGNAL Logical_Operator_out245_out1            : std_logic;
  SIGNAL Logical_Operator_out246_out1            : std_logic;
  SIGNAL Logical_Operator_out247_out1            : std_logic;
  SIGNAL Logical_Operator_out248_out1            : std_logic;
  SIGNAL Logical_Operator_out249_out1            : std_logic;
  SIGNAL Logical_Operator_out250_out1            : std_logic;
  SIGNAL Logical_Operator_out251_out1            : std_logic;
  SIGNAL Logical_Operator_out252_out1            : std_logic;
  SIGNAL Logical_Operator_out253_out1            : std_logic;
  SIGNAL Logical_Operator_out254_out1            : std_logic;
  SIGNAL Logical_Operator_out255_out1            : std_logic;
  SIGNAL Logical_Operator_out256_out1            : std_logic;
  SIGNAL Logical_Operator_out257_out1            : std_logic;
  SIGNAL Logical_Operator_out258_out1            : std_logic;
  SIGNAL Logical_Operator_out259_out1            : std_logic;
  SIGNAL Logical_Operator_out260_out1            : std_logic;
  SIGNAL Logical_Operator_out261_out1            : std_logic;
  SIGNAL Logical_Operator_out262_out1            : std_logic;
  SIGNAL Logical_Operator_out263_out1            : std_logic;
  SIGNAL Logical_Operator_out264_out1            : std_logic;
  SIGNAL Logical_Operator_out265_out1            : std_logic;
  SIGNAL Logical_Operator_out266_out1            : std_logic;
  SIGNAL Logical_Operator_out267_out1            : std_logic;
  SIGNAL Logical_Operator_out268_out1            : std_logic;
  SIGNAL Logical_Operator_out269_out1            : std_logic;
  SIGNAL Logical_Operator_out270_out1            : std_logic;
  SIGNAL Logical_Operator_out271_out1            : std_logic;
  SIGNAL Logical_Operator_out272_out1            : std_logic;
  SIGNAL Logical_Operator_out273_out1            : std_logic;
  SIGNAL Logical_Operator_out274_out1            : std_logic;
  SIGNAL Logical_Operator_out275_out1            : std_logic;
  SIGNAL Logical_Operator_out276_out1            : std_logic;
  SIGNAL Logical_Operator_out277_out1            : std_logic;
  SIGNAL Logical_Operator_out278_out1            : std_logic;
  SIGNAL Logical_Operator_out279_out1            : std_logic;
  SIGNAL Logical_Operator_out280_out1            : std_logic;
  SIGNAL Logical_Operator_out281_out1            : std_logic;
  SIGNAL Logical_Operator_out282_out1            : std_logic;
  SIGNAL Logical_Operator_out283_out1            : std_logic;
  SIGNAL Logical_Operator_out284_out1            : std_logic;
  SIGNAL Logical_Operator_out285_out1            : std_logic;
  SIGNAL Logical_Operator_out286_out1            : std_logic;
  SIGNAL Logical_Operator_out287_out1            : std_logic;
  SIGNAL Logical_Operator_out288_out1            : std_logic;
  SIGNAL Logical_Operator_out289_out1            : std_logic;
  SIGNAL Logical_Operator_out290_out1            : std_logic;
  SIGNAL Logical_Operator_out291_out1            : std_logic;
  SIGNAL Logical_Operator_out292_out1            : std_logic;
  SIGNAL Logical_Operator_out293_out1            : std_logic;
  SIGNAL Logical_Operator_out294_out1            : std_logic;
  SIGNAL Logical_Operator_out295_out1            : std_logic;
  SIGNAL Logical_Operator_out296_out1            : std_logic;
  SIGNAL Logical_Operator_out297_out1            : std_logic;
  SIGNAL Logical_Operator_out298_out1            : std_logic;
  SIGNAL Logical_Operator_out299_out1            : std_logic;
  SIGNAL Logical_Operator_out300_out1            : std_logic;
  SIGNAL Logical_Operator_out301_out1            : std_logic;
  SIGNAL Logical_Operator_out302_out1            : std_logic;
  SIGNAL Logical_Operator_out303_out1            : std_logic;
  SIGNAL Logical_Operator_out304_out1            : std_logic;
  SIGNAL Logical_Operator_out305_out1            : std_logic;
  SIGNAL Logical_Operator_out306_out1            : std_logic;
  SIGNAL Logical_Operator_out307_out1            : std_logic;
  SIGNAL Logical_Operator_out308_out1            : std_logic;
  SIGNAL Logical_Operator_out309_out1            : std_logic;
  SIGNAL Logical_Operator_out310_out1            : std_logic;
  SIGNAL Logical_Operator_out311_out1            : std_logic;
  SIGNAL Logical_Operator_out312_out1            : std_logic;
  SIGNAL Logical_Operator_out313_out1            : std_logic;
  SIGNAL Logical_Operator_out314_out1            : std_logic;
  SIGNAL Logical_Operator_out315_out1            : std_logic;
  SIGNAL Logical_Operator_out316_out1            : std_logic;
  SIGNAL Logical_Operator_out317_out1            : std_logic;
  SIGNAL Logical_Operator_out318_out1            : std_logic;
  SIGNAL Logical_Operator_out319_out1            : std_logic;
  SIGNAL Logical_Operator_out320_out1            : std_logic;
  SIGNAL Logical_Operator_out321_out1            : std_logic;
  SIGNAL Logical_Operator_out322_out1            : std_logic;
  SIGNAL Logical_Operator_out323_out1            : std_logic;
  SIGNAL Logical_Operator_out324_out1            : std_logic;
  SIGNAL Logical_Operator_out325_out1            : std_logic;
  SIGNAL Logical_Operator_out326_out1            : std_logic;
  SIGNAL Logical_Operator_out327_out1            : std_logic;
  SIGNAL Logical_Operator_out328_out1            : std_logic;
  SIGNAL Logical_Operator_out329_out1            : std_logic;
  SIGNAL Logical_Operator_out330_out1            : std_logic;
  SIGNAL Logical_Operator_out331_out1            : std_logic;
  SIGNAL Logical_Operator_out332_out1            : std_logic;
  SIGNAL Logical_Operator_out333_out1            : std_logic;
  SIGNAL Logical_Operator_out334_out1            : std_logic;
  SIGNAL Logical_Operator_out335_out1            : std_logic;
  SIGNAL Logical_Operator_out336_out1            : std_logic;
  SIGNAL Logical_Operator_out337_out1            : std_logic;
  SIGNAL Logical_Operator_out338_out1            : std_logic;
  SIGNAL Logical_Operator_out339_out1            : std_logic;
  SIGNAL Logical_Operator_out340_out1            : std_logic;
  SIGNAL Logical_Operator_out341_out1            : std_logic;
  SIGNAL Logical_Operator_out342_out1            : std_logic;
  SIGNAL Logical_Operator_out343_out1            : std_logic;
  SIGNAL Logical_Operator_out344_out1            : std_logic;
  SIGNAL Logical_Operator_out345_out1            : std_logic;
  SIGNAL Logical_Operator_out346_out1            : std_logic;
  SIGNAL Logical_Operator_out347_out1            : std_logic;
  SIGNAL Logical_Operator_out348_out1            : std_logic;
  SIGNAL Logical_Operator_out349_out1            : std_logic;
  SIGNAL Logical_Operator_out350_out1            : std_logic;
  SIGNAL Logical_Operator_out351_out1            : std_logic;
  SIGNAL Logical_Operator_out352_out1            : std_logic;
  SIGNAL Logical_Operator_out353_out1            : std_logic;
  SIGNAL Logical_Operator_out354_out1            : std_logic;
  SIGNAL Logical_Operator_out355_out1            : std_logic;
  SIGNAL Logical_Operator_out356_out1            : std_logic;
  SIGNAL Logical_Operator_out357_out1            : std_logic;
  SIGNAL Logical_Operator_out358_out1            : std_logic;
  SIGNAL Logical_Operator_out359_out1            : std_logic;
  SIGNAL Logical_Operator_out360_out1            : std_logic;
  SIGNAL Logical_Operator_out361_out1            : std_logic;
  SIGNAL Logical_Operator_out362_out1            : std_logic;
  SIGNAL Logical_Operator_out363_out1            : std_logic;
  SIGNAL Logical_Operator_out364_out1            : std_logic;
  SIGNAL Logical_Operator_out365_out1            : std_logic;
  SIGNAL Logical_Operator_out366_out1            : std_logic;
  SIGNAL Logical_Operator_out367_out1            : std_logic;
  SIGNAL Logical_Operator_out368_out1            : std_logic;
  SIGNAL Logical_Operator_out369_out1            : std_logic;
  SIGNAL Logical_Operator_out370_out1            : std_logic;
  SIGNAL Logical_Operator_out371_out1            : std_logic;
  SIGNAL Logical_Operator_out372_out1            : std_logic;
  SIGNAL Logical_Operator_out373_out1            : std_logic;
  SIGNAL Logical_Operator_out374_out1            : std_logic;
  SIGNAL Logical_Operator_out375_out1            : std_logic;
  SIGNAL Logical_Operator_out376_out1            : std_logic;
  SIGNAL Logical_Operator_out377_out1            : std_logic;
  SIGNAL Logical_Operator_out378_out1            : std_logic;
  SIGNAL Logical_Operator_out379_out1            : std_logic;
  SIGNAL Logical_Operator_out380_out1            : std_logic;
  SIGNAL Logical_Operator_out381_out1            : std_logic;
  SIGNAL Logical_Operator_out382_out1            : std_logic;
  SIGNAL Logical_Operator_out383_out1            : std_logic;
  SIGNAL Logical_Operator_out384_out1            : std_logic;
  SIGNAL Logical_Operator_out385_out1            : std_logic;
  SIGNAL Logical_Operator_out386_out1            : std_logic;
  SIGNAL Logical_Operator_out387_out1            : std_logic;
  SIGNAL Logical_Operator_out388_out1            : std_logic;
  SIGNAL Logical_Operator_out389_out1            : std_logic;
  SIGNAL Logical_Operator_out390_out1            : std_logic;
  SIGNAL Logical_Operator_out391_out1            : std_logic;
  SIGNAL Logical_Operator_out392_out1            : std_logic;
  SIGNAL Logical_Operator_out393_out1            : std_logic;
  SIGNAL Logical_Operator_out394_out1            : std_logic;
  SIGNAL Logical_Operator_out395_out1            : std_logic;
  SIGNAL Logical_Operator_out396_out1            : std_logic;
  SIGNAL Logical_Operator_out397_out1            : std_logic;
  SIGNAL Logical_Operator_out398_out1            : std_logic;
  SIGNAL Logical_Operator_out399_out1            : std_logic;
  SIGNAL Logical_Operator_out400_out1            : std_logic;
  SIGNAL Logical_Operator_out401_out1            : std_logic;
  SIGNAL Logical_Operator_out402_out1            : std_logic;
  SIGNAL Logical_Operator_out403_out1            : std_logic;
  SIGNAL Logical_Operator_out404_out1            : std_logic;
  SIGNAL Logical_Operator_out405_out1            : std_logic;
  SIGNAL Logical_Operator_out406_out1            : std_logic;
  SIGNAL Logical_Operator_out407_out1            : std_logic;
  SIGNAL Logical_Operator_out408_out1            : std_logic;
  SIGNAL Logical_Operator_out409_out1            : std_logic;
  SIGNAL Logical_Operator_out410_out1            : std_logic;
  SIGNAL Logical_Operator_out411_out1            : std_logic;
  SIGNAL Logical_Operator_out412_out1            : std_logic;
  SIGNAL Logical_Operator_out413_out1            : std_logic;
  SIGNAL Logical_Operator_out414_out1            : std_logic;
  SIGNAL Logical_Operator_out415_out1            : std_logic;
  SIGNAL Logical_Operator_out416_out1            : std_logic;
  SIGNAL Logical_Operator_out417_out1            : std_logic;
  SIGNAL Logical_Operator_out418_out1            : std_logic;
  SIGNAL Logical_Operator_out419_out1            : std_logic;
  SIGNAL Logical_Operator_out420_out1            : std_logic;
  SIGNAL Logical_Operator_out421_out1            : std_logic;
  SIGNAL Logical_Operator_out422_out1            : std_logic;
  SIGNAL Logical_Operator_out423_out1            : std_logic;
  SIGNAL Logical_Operator_out424_out1            : std_logic;
  SIGNAL Logical_Operator_out425_out1            : std_logic;
  SIGNAL Logical_Operator_out426_out1            : std_logic;
  SIGNAL Logical_Operator_out427_out1            : std_logic;
  SIGNAL Logical_Operator_out428_out1            : std_logic;
  SIGNAL Logical_Operator_out429_out1            : std_logic;
  SIGNAL Logical_Operator_out430_out1            : std_logic;
  SIGNAL Logical_Operator_out431_out1            : std_logic;
  SIGNAL Logical_Operator_out432_out1            : std_logic;
  SIGNAL Logical_Operator_out433_out1            : std_logic;
  SIGNAL Logical_Operator_out434_out1            : std_logic;
  SIGNAL Logical_Operator_out435_out1            : std_logic;
  SIGNAL Logical_Operator_out436_out1            : std_logic;
  SIGNAL Logical_Operator_out437_out1            : std_logic;
  SIGNAL Logical_Operator_out438_out1            : std_logic;
  SIGNAL Logical_Operator_out439_out1            : std_logic;
  SIGNAL Logical_Operator_out440_out1            : std_logic;
  SIGNAL Logical_Operator_out441_out1            : std_logic;
  SIGNAL Logical_Operator_out442_out1            : std_logic;
  SIGNAL Logical_Operator_out443_out1            : std_logic;
  SIGNAL Logical_Operator_out444_out1            : std_logic;
  SIGNAL Logical_Operator_out445_out1            : std_logic;
  SIGNAL Logical_Operator_out446_out1            : std_logic;
  SIGNAL Logical_Operator_out447_out1            : std_logic;
  SIGNAL Logical_Operator_out448_out1            : std_logic;
  SIGNAL Logical_Operator_out449_out1            : std_logic;
  SIGNAL Logical_Operator_out450_out1            : std_logic;
  SIGNAL Logical_Operator_out451_out1            : std_logic;
  SIGNAL Logical_Operator_out452_out1            : std_logic;
  SIGNAL Logical_Operator_out453_out1            : std_logic;
  SIGNAL Logical_Operator_out454_out1            : std_logic;
  SIGNAL Logical_Operator_out455_out1            : std_logic;
  SIGNAL Logical_Operator_out456_out1            : std_logic;
  SIGNAL Logical_Operator_out457_out1            : std_logic;
  SIGNAL Logical_Operator_out458_out1            : std_logic;
  SIGNAL Logical_Operator_out459_out1            : std_logic;
  SIGNAL Logical_Operator_out460_out1            : std_logic;
  SIGNAL Logical_Operator_out461_out1            : std_logic;
  SIGNAL Logical_Operator_out462_out1            : std_logic;
  SIGNAL Logical_Operator_out463_out1            : std_logic;
  SIGNAL Logical_Operator_out464_out1            : std_logic;
  SIGNAL Logical_Operator_out465_out1            : std_logic;
  SIGNAL Logical_Operator_out466_out1            : std_logic;
  SIGNAL Logical_Operator_out467_out1            : std_logic;
  SIGNAL Logical_Operator_out468_out1            : std_logic;
  SIGNAL Logical_Operator_out469_out1            : std_logic;
  SIGNAL Logical_Operator_out470_out1            : std_logic;
  SIGNAL Logical_Operator_out471_out1            : std_logic;
  SIGNAL Logical_Operator_out472_out1            : std_logic;
  SIGNAL Logical_Operator_out473_out1            : std_logic;
  SIGNAL Logical_Operator_out474_out1            : std_logic;
  SIGNAL Logical_Operator_out475_out1            : std_logic;
  SIGNAL Logical_Operator_out476_out1            : std_logic;
  SIGNAL Logical_Operator_out477_out1            : std_logic;
  SIGNAL Logical_Operator_out478_out1            : std_logic;
  SIGNAL Logical_Operator_out479_out1            : std_logic;
  SIGNAL Logical_Operator_out480_out1            : std_logic;
  SIGNAL Logical_Operator_out481_out1            : std_logic;
  SIGNAL Logical_Operator_out482_out1            : std_logic;
  SIGNAL Logical_Operator_out483_out1            : std_logic;
  SIGNAL Logical_Operator_out484_out1            : std_logic;
  SIGNAL Logical_Operator_out485_out1            : std_logic;
  SIGNAL Logical_Operator_out486_out1            : std_logic;
  SIGNAL Logical_Operator_out487_out1            : std_logic;
  SIGNAL Logical_Operator_out488_out1            : std_logic;
  SIGNAL Logical_Operator_out489_out1            : std_logic;
  SIGNAL Logical_Operator_out490_out1            : std_logic;
  SIGNAL Logical_Operator_out491_out1            : std_logic;
  SIGNAL Logical_Operator_out492_out1            : std_logic;
  SIGNAL Logical_Operator_out493_out1            : std_logic;
  SIGNAL Logical_Operator_out494_out1            : std_logic;
  SIGNAL Logical_Operator_out495_out1            : std_logic;
  SIGNAL Logical_Operator_out496_out1            : std_logic;
  SIGNAL Logical_Operator_out497_out1            : std_logic;
  SIGNAL Logical_Operator_out498_out1            : std_logic;
  SIGNAL Logical_Operator_out499_out1            : std_logic;
  SIGNAL Logical_Operator_out500_out1            : std_logic;
  SIGNAL Logical_Operator_out501_out1            : std_logic;
  SIGNAL Logical_Operator_out502_out1            : std_logic;
  SIGNAL Logical_Operator_out503_out1            : std_logic;
  SIGNAL Logical_Operator_out504_out1            : std_logic;
  SIGNAL Logical_Operator_out505_out1            : std_logic;
  SIGNAL Logical_Operator_out506_out1            : std_logic;
  SIGNAL Logical_Operator_out507_out1            : std_logic;
  SIGNAL Logical_Operator_out508_out1            : std_logic;
  SIGNAL Logical_Operator_out509_out1            : std_logic;
  SIGNAL Logical_Operator_out510_out1            : std_logic;
  SIGNAL Logical_Operator_out511_out1            : std_logic;
  SIGNAL Logical_Operator_out512_out1            : std_logic;
  SIGNAL Logical_Operator_out513_out1            : std_logic;
  SIGNAL Logical_Operator_out514_out1            : std_logic;
  SIGNAL Logical_Operator_out515_out1            : std_logic;
  SIGNAL Logical_Operator_out516_out1            : std_logic;
  SIGNAL Logical_Operator_out517_out1            : std_logic;
  SIGNAL Logical_Operator_out518_out1            : std_logic;
  SIGNAL Logical_Operator_out519_out1            : std_logic;
  SIGNAL Logical_Operator_out520_out1            : std_logic;
  SIGNAL Logical_Operator_out521_out1            : std_logic;
  SIGNAL Logical_Operator_out522_out1            : std_logic;
  SIGNAL Logical_Operator_out523_out1            : std_logic;
  SIGNAL Logical_Operator_out524_out1            : std_logic;
  SIGNAL Logical_Operator_out525_out1            : std_logic;
  SIGNAL Logical_Operator_out526_out1            : std_logic;
  SIGNAL Logical_Operator_out527_out1            : std_logic;
  SIGNAL Logical_Operator_out528_out1            : std_logic;
  SIGNAL Logical_Operator_out529_out1            : std_logic;
  SIGNAL Logical_Operator_out530_out1            : std_logic;
  SIGNAL Logical_Operator_out531_out1            : std_logic;
  SIGNAL Logical_Operator_out532_out1            : std_logic;
  SIGNAL Logical_Operator_out533_out1            : std_logic;
  SIGNAL Logical_Operator_out534_out1            : std_logic;
  SIGNAL Logical_Operator_out535_out1            : std_logic;
  SIGNAL Logical_Operator_out536_out1            : std_logic;
  SIGNAL Logical_Operator_out537_out1            : std_logic;
  SIGNAL Logical_Operator_out538_out1            : std_logic;
  SIGNAL Logical_Operator_out539_out1            : std_logic;
  SIGNAL Logical_Operator_out540_out1            : std_logic;
  SIGNAL Logical_Operator_out541_out1            : std_logic;
  SIGNAL Logical_Operator_out542_out1            : std_logic;
  SIGNAL Logical_Operator_out543_out1            : std_logic;
  SIGNAL Logical_Operator_out544_out1            : std_logic;
  SIGNAL Logical_Operator_out545_out1            : std_logic;
  SIGNAL Logical_Operator_out546_out1            : std_logic;
  SIGNAL Logical_Operator_out547_out1            : std_logic;
  SIGNAL Logical_Operator_out548_out1            : std_logic;
  SIGNAL Logical_Operator_out549_out1            : std_logic;
  SIGNAL Logical_Operator_out550_out1            : std_logic;
  SIGNAL Logical_Operator_out551_out1            : std_logic;
  SIGNAL Logical_Operator_out552_out1            : std_logic;
  SIGNAL Logical_Operator_out553_out1            : std_logic;
  SIGNAL Logical_Operator_out554_out1            : std_logic;
  SIGNAL Logical_Operator_out555_out1            : std_logic;
  SIGNAL Logical_Operator_out556_out1            : std_logic;
  SIGNAL Logical_Operator_out557_out1            : std_logic;
  SIGNAL Logical_Operator_out558_out1            : std_logic;
  SIGNAL Logical_Operator_out559_out1            : std_logic;
  SIGNAL Logical_Operator_out560_out1            : std_logic;
  SIGNAL Logical_Operator_out561_out1            : std_logic;
  SIGNAL Logical_Operator_out562_out1            : std_logic;
  SIGNAL Logical_Operator_out563_out1            : std_logic;
  SIGNAL Logical_Operator_out564_out1            : std_logic;
  SIGNAL Logical_Operator_out565_out1            : std_logic;
  SIGNAL Logical_Operator_out566_out1            : std_logic;
  SIGNAL Logical_Operator_out567_out1            : std_logic;
  SIGNAL Logical_Operator_out568_out1            : std_logic;
  SIGNAL Logical_Operator_out569_out1            : std_logic;
  SIGNAL Logical_Operator_out570_out1            : std_logic;
  SIGNAL Logical_Operator_out571_out1            : std_logic;
  SIGNAL Logical_Operator_out572_out1            : std_logic;
  SIGNAL Logical_Operator_out573_out1            : std_logic;
  SIGNAL Logical_Operator_out574_out1            : std_logic;
  SIGNAL Logical_Operator_out575_out1            : std_logic;
  SIGNAL Logical_Operator_out576_out1            : std_logic;
  SIGNAL Logical_Operator_out577_out1            : std_logic;
  SIGNAL Logical_Operator_out578_out1            : std_logic;
  SIGNAL Logical_Operator_out579_out1            : std_logic;
  SIGNAL Logical_Operator_out580_out1            : std_logic;
  SIGNAL Logical_Operator_out581_out1            : std_logic;
  SIGNAL Logical_Operator_out582_out1            : std_logic;
  SIGNAL Logical_Operator_out583_out1            : std_logic;
  SIGNAL Logical_Operator_out584_out1            : std_logic;
  SIGNAL Logical_Operator_out585_out1            : std_logic;
  SIGNAL Logical_Operator_out586_out1            : std_logic;
  SIGNAL Logical_Operator_out587_out1            : std_logic;
  SIGNAL Logical_Operator_out588_out1            : std_logic;
  SIGNAL Logical_Operator_out589_out1            : std_logic;
  SIGNAL Logical_Operator_out590_out1            : std_logic;
  SIGNAL Logical_Operator_out591_out1            : std_logic;
  SIGNAL Logical_Operator_out592_out1            : std_logic;
  SIGNAL Logical_Operator_out593_out1            : std_logic;
  SIGNAL Logical_Operator_out594_out1            : std_logic;
  SIGNAL Logical_Operator_out595_out1            : std_logic;
  SIGNAL Logical_Operator_out596_out1            : std_logic;
  SIGNAL Logical_Operator_out597_out1            : std_logic;
  SIGNAL Logical_Operator_out598_out1            : std_logic;
  SIGNAL Logical_Operator_out599_out1            : std_logic;
  SIGNAL Logical_Operator_out600_out1            : std_logic;
  SIGNAL Logical_Operator_out601_out1            : std_logic;
  SIGNAL Logical_Operator_out602_out1            : std_logic;
  SIGNAL Logical_Operator_out603_out1            : std_logic;
  SIGNAL Logical_Operator_out604_out1            : std_logic;
  SIGNAL Logical_Operator_out605_out1            : std_logic;
  SIGNAL Logical_Operator_out606_out1            : std_logic;
  SIGNAL Logical_Operator_out607_out1            : std_logic;
  SIGNAL Logical_Operator_out608_out1            : std_logic;
  SIGNAL Logical_Operator_out609_out1            : std_logic;
  SIGNAL Logical_Operator_out610_out1            : std_logic;
  SIGNAL Logical_Operator_out611_out1            : std_logic;
  SIGNAL Logical_Operator_out612_out1            : std_logic;
  SIGNAL Logical_Operator_out613_out1            : std_logic;
  SIGNAL Logical_Operator_out614_out1            : std_logic;
  SIGNAL Logical_Operator_out615_out1            : std_logic;
  SIGNAL Logical_Operator_out616_out1            : std_logic;
  SIGNAL Logical_Operator_out617_out1            : std_logic;
  SIGNAL Logical_Operator_out618_out1            : std_logic;
  SIGNAL Logical_Operator_out619_out1            : std_logic;
  SIGNAL Logical_Operator_out620_out1            : std_logic;
  SIGNAL Logical_Operator_out621_out1            : std_logic;
  SIGNAL Logical_Operator_out622_out1            : std_logic;
  SIGNAL Logical_Operator_out623_out1            : std_logic;
  SIGNAL Logical_Operator_out624_out1            : std_logic;
  SIGNAL Logical_Operator_out625_out1            : std_logic;
  SIGNAL Logical_Operator_out626_out1            : std_logic;
  SIGNAL Logical_Operator_out627_out1            : std_logic;
  SIGNAL Logical_Operator_out628_out1            : std_logic;
  SIGNAL Logical_Operator_out629_out1            : std_logic;
  SIGNAL Logical_Operator_out630_out1            : std_logic;
  SIGNAL Logical_Operator_out631_out1            : std_logic;
  SIGNAL Logical_Operator_out632_out1            : std_logic;
  SIGNAL Logical_Operator_out633_out1            : std_logic;
  SIGNAL Logical_Operator_out634_out1            : std_logic;
  SIGNAL Logical_Operator_out635_out1            : std_logic;
  SIGNAL Logical_Operator_out636_out1            : std_logic;
  SIGNAL Logical_Operator_out637_out1            : std_logic;
  SIGNAL Logical_Operator_out638_out1            : std_logic;
  SIGNAL Logical_Operator_out639_out1            : std_logic;
  SIGNAL Logical_Operator_out640_out1            : std_logic;
  SIGNAL Logical_Operator_out641_out1            : std_logic;
  SIGNAL Logical_Operator_out642_out1            : std_logic;
  SIGNAL Logical_Operator_out643_out1            : std_logic;
  SIGNAL Logical_Operator_out644_out1            : std_logic;
  SIGNAL Logical_Operator_out645_out1            : std_logic;
  SIGNAL Logical_Operator_out646_out1            : std_logic;
  SIGNAL Logical_Operator_out647_out1            : std_logic;
  SIGNAL Logical_Operator_out648_out1            : std_logic;
  SIGNAL Logical_Operator_out649_out1            : std_logic;
  SIGNAL Logical_Operator_out650_out1            : std_logic;
  SIGNAL Logical_Operator_out651_out1            : std_logic;
  SIGNAL Logical_Operator_out652_out1            : std_logic;
  SIGNAL Logical_Operator_out653_out1            : std_logic;
  SIGNAL Logical_Operator_out654_out1            : std_logic;
  SIGNAL Logical_Operator_out655_out1            : std_logic;
  SIGNAL Logical_Operator_out656_out1            : std_logic;
  SIGNAL Logical_Operator_out657_out1            : std_logic;
  SIGNAL Logical_Operator_out658_out1            : std_logic;
  SIGNAL Logical_Operator_out659_out1            : std_logic;
  SIGNAL Logical_Operator_out660_out1            : std_logic;
  SIGNAL Logical_Operator_out661_out1            : std_logic;
  SIGNAL Logical_Operator_out662_out1            : std_logic;
  SIGNAL Logical_Operator_out663_out1            : std_logic;
  SIGNAL Logical_Operator_out664_out1            : std_logic;
  SIGNAL Logical_Operator_out665_out1            : std_logic;
  SIGNAL Logical_Operator_out666_out1            : std_logic;
  SIGNAL Logical_Operator_out667_out1            : std_logic;
  SIGNAL Logical_Operator_out668_out1            : std_logic;
  SIGNAL Logical_Operator_out669_out1            : std_logic;
  SIGNAL Logical_Operator_out670_out1            : std_logic;
  SIGNAL Logical_Operator_out671_out1            : std_logic;
  SIGNAL Logical_Operator_out672_out1            : std_logic;
  SIGNAL Logical_Operator_out673_out1            : std_logic;
  SIGNAL Logical_Operator_out674_out1            : std_logic;
  SIGNAL Logical_Operator_out675_out1            : std_logic;
  SIGNAL Logical_Operator_out676_out1            : std_logic;
  SIGNAL Logical_Operator_out677_out1            : std_logic;
  SIGNAL Logical_Operator_out678_out1            : std_logic;
  SIGNAL Logical_Operator_out679_out1            : std_logic;
  SIGNAL Logical_Operator_out680_out1            : std_logic;
  SIGNAL Logical_Operator_out681_out1            : std_logic;
  SIGNAL Logical_Operator_out682_out1            : std_logic;
  SIGNAL Logical_Operator_out683_out1            : std_logic;
  SIGNAL Logical_Operator_out684_out1            : std_logic;
  SIGNAL Logical_Operator_out685_out1            : std_logic;
  SIGNAL Logical_Operator_out686_out1            : std_logic;
  SIGNAL Logical_Operator_out687_out1            : std_logic;
  SIGNAL Logical_Operator_out688_out1            : std_logic;
  SIGNAL Logical_Operator_out689_out1            : std_logic;
  SIGNAL Logical_Operator_out690_out1            : std_logic;
  SIGNAL Logical_Operator_out691_out1            : std_logic;
  SIGNAL Logical_Operator_out692_out1            : std_logic;
  SIGNAL Logical_Operator_out693_out1            : std_logic;
  SIGNAL Logical_Operator_out694_out1            : std_logic;
  SIGNAL Logical_Operator_out695_out1            : std_logic;
  SIGNAL Logical_Operator_out696_out1            : std_logic;
  SIGNAL Logical_Operator_out697_out1            : std_logic;
  SIGNAL Logical_Operator_out698_out1            : std_logic;
  SIGNAL Logical_Operator_out699_out1            : std_logic;
  SIGNAL Logical_Operator_out700_out1            : std_logic;
  SIGNAL Logical_Operator_out701_out1            : std_logic;
  SIGNAL Logical_Operator_out702_out1            : std_logic;
  SIGNAL Logical_Operator_out703_out1            : std_logic;
  SIGNAL Logical_Operator_out704_out1            : std_logic;
  SIGNAL Logical_Operator_out705_out1            : std_logic;
  SIGNAL Logical_Operator_out706_out1            : std_logic;
  SIGNAL Logical_Operator_out707_out1            : std_logic;
  SIGNAL Logical_Operator_out708_out1            : std_logic;
  SIGNAL Logical_Operator_out709_out1            : std_logic;
  SIGNAL Logical_Operator_out710_out1            : std_logic;
  SIGNAL Logical_Operator_out711_out1            : std_logic;
  SIGNAL Logical_Operator_out712_out1            : std_logic;
  SIGNAL Logical_Operator_out713_out1            : std_logic;
  SIGNAL Logical_Operator_out714_out1            : std_logic;
  SIGNAL Logical_Operator_out715_out1            : std_logic;
  SIGNAL Logical_Operator_out716_out1            : std_logic;
  SIGNAL Logical_Operator_out717_out1            : std_logic;
  SIGNAL Logical_Operator_out718_out1            : std_logic;
  SIGNAL Logical_Operator_out719_out1            : std_logic;
  SIGNAL Logical_Operator_out720_out1            : std_logic;
  SIGNAL Logical_Operator_out721_out1            : std_logic;
  SIGNAL Logical_Operator_out722_out1            : std_logic;
  SIGNAL Logical_Operator_out723_out1            : std_logic;
  SIGNAL Logical_Operator_out724_out1            : std_logic;
  SIGNAL Logical_Operator_out725_out1            : std_logic;
  SIGNAL Logical_Operator_out726_out1            : std_logic;
  SIGNAL Logical_Operator_out727_out1            : std_logic;
  SIGNAL Logical_Operator_out728_out1            : std_logic;
  SIGNAL Logical_Operator_out729_out1            : std_logic;
  SIGNAL Logical_Operator_out730_out1            : std_logic;
  SIGNAL Logical_Operator_out731_out1            : std_logic;
  SIGNAL Logical_Operator_out732_out1            : std_logic;
  SIGNAL Logical_Operator_out733_out1            : std_logic;
  SIGNAL Logical_Operator_out734_out1            : std_logic;
  SIGNAL Logical_Operator_out735_out1            : std_logic;
  SIGNAL Logical_Operator_out736_out1            : std_logic;
  SIGNAL Logical_Operator_out737_out1            : std_logic;
  SIGNAL Logical_Operator_out738_out1            : std_logic;
  SIGNAL Logical_Operator_out739_out1            : std_logic;
  SIGNAL Logical_Operator_out740_out1            : std_logic;
  SIGNAL Logical_Operator_out741_out1            : std_logic;
  SIGNAL Logical_Operator_out742_out1            : std_logic;
  SIGNAL Logical_Operator_out743_out1            : std_logic;
  SIGNAL Logical_Operator_out744_out1            : std_logic;
  SIGNAL Logical_Operator_out745_out1            : std_logic;
  SIGNAL Logical_Operator_out746_out1            : std_logic;
  SIGNAL Logical_Operator_out747_out1            : std_logic;
  SIGNAL Logical_Operator_out748_out1            : std_logic;
  SIGNAL Logical_Operator_out749_out1            : std_logic;
  SIGNAL Logical_Operator_out750_out1            : std_logic;
  SIGNAL Logical_Operator_out751_out1            : std_logic;
  SIGNAL Logical_Operator_out752_out1            : std_logic;
  SIGNAL Logical_Operator_out753_out1            : std_logic;
  SIGNAL Logical_Operator_out754_out1            : std_logic;
  SIGNAL Logical_Operator_out755_out1            : std_logic;
  SIGNAL Logical_Operator_out756_out1            : std_logic;
  SIGNAL Logical_Operator_out757_out1            : std_logic;
  SIGNAL Logical_Operator_out758_out1            : std_logic;
  SIGNAL Logical_Operator_out759_out1            : std_logic;
  SIGNAL Logical_Operator_out760_out1            : std_logic;
  SIGNAL Logical_Operator_out761_out1            : std_logic;
  SIGNAL Logical_Operator_out762_out1            : std_logic;
  SIGNAL Logical_Operator_out763_out1            : std_logic;
  SIGNAL Logical_Operator_out764_out1            : std_logic;
  SIGNAL Logical_Operator_out765_out1            : std_logic;
  SIGNAL Logical_Operator_out766_out1            : std_logic;
  SIGNAL Logical_Operator_out767_out1            : std_logic;
  SIGNAL Logical_Operator_out768_out1            : std_logic;
  SIGNAL Logical_Operator_out769_out1            : std_logic;
  SIGNAL Logical_Operator_out770_out1            : std_logic;
  SIGNAL Logical_Operator_out771_out1            : std_logic;
  SIGNAL Logical_Operator_out772_out1            : std_logic;
  SIGNAL Logical_Operator_out773_out1            : std_logic;
  SIGNAL Logical_Operator_out774_out1            : std_logic;
  SIGNAL Logical_Operator_out775_out1            : std_logic;
  SIGNAL Logical_Operator_out776_out1            : std_logic;
  SIGNAL Logical_Operator_out777_out1            : std_logic;
  SIGNAL Logical_Operator_out778_out1            : std_logic;
  SIGNAL Logical_Operator_out779_out1            : std_logic;
  SIGNAL Logical_Operator_out780_out1            : std_logic;
  SIGNAL Logical_Operator_out781_out1            : std_logic;
  SIGNAL Logical_Operator_out782_out1            : std_logic;
  SIGNAL Logical_Operator_out783_out1            : std_logic;
  SIGNAL Logical_Operator_out784_out1            : std_logic;
  SIGNAL Logical_Operator_out785_out1            : std_logic;
  SIGNAL Logical_Operator_out786_out1            : std_logic;
  SIGNAL Logical_Operator_out787_out1            : std_logic;
  SIGNAL Logical_Operator_out788_out1            : std_logic;
  SIGNAL Logical_Operator_out789_out1            : std_logic;
  SIGNAL Logical_Operator_out790_out1            : std_logic;
  SIGNAL Logical_Operator_out791_out1            : std_logic;
  SIGNAL Logical_Operator_out792_out1            : std_logic;
  SIGNAL Logical_Operator_out793_out1            : std_logic;
  SIGNAL Logical_Operator_out794_out1            : std_logic;
  SIGNAL Logical_Operator_out795_out1            : std_logic;
  SIGNAL Logical_Operator_out796_out1            : std_logic;
  SIGNAL Logical_Operator_out797_out1            : std_logic;
  SIGNAL Logical_Operator_out798_out1            : std_logic;
  SIGNAL Logical_Operator_out799_out1            : std_logic;
  SIGNAL Logical_Operator_out800_out1            : std_logic;
  SIGNAL Logical_Operator_out801_out1            : std_logic;
  SIGNAL Logical_Operator_out802_out1            : std_logic;
  SIGNAL Logical_Operator_out803_out1            : std_logic;
  SIGNAL Logical_Operator_out804_out1            : std_logic;
  SIGNAL Logical_Operator_out805_out1            : std_logic;
  SIGNAL Logical_Operator_out806_out1            : std_logic;
  SIGNAL Logical_Operator_out807_out1            : std_logic;
  SIGNAL Logical_Operator_out808_out1            : std_logic;
  SIGNAL Logical_Operator_out809_out1            : std_logic;
  SIGNAL Logical_Operator_out810_out1            : std_logic;
  SIGNAL Logical_Operator_out811_out1            : std_logic;
  SIGNAL Logical_Operator_out812_out1            : std_logic;
  SIGNAL Logical_Operator_out813_out1            : std_logic;
  SIGNAL Logical_Operator_out814_out1            : std_logic;
  SIGNAL Logical_Operator_out815_out1            : std_logic;
  SIGNAL Logical_Operator_out816_out1            : std_logic;
  SIGNAL Logical_Operator_out817_out1            : std_logic;
  SIGNAL Logical_Operator_out818_out1            : std_logic;
  SIGNAL Logical_Operator_out819_out1            : std_logic;
  SIGNAL Logical_Operator_out820_out1            : std_logic;
  SIGNAL Logical_Operator_out821_out1            : std_logic;
  SIGNAL Logical_Operator_out822_out1            : std_logic;
  SIGNAL Logical_Operator_out823_out1            : std_logic;
  SIGNAL Logical_Operator_out824_out1            : std_logic;
  SIGNAL Logical_Operator_out825_out1            : std_logic;
  SIGNAL Logical_Operator_out826_out1            : std_logic;
  SIGNAL Logical_Operator_out827_out1            : std_logic;
  SIGNAL Logical_Operator_out828_out1            : std_logic;
  SIGNAL Logical_Operator_out829_out1            : std_logic;
  SIGNAL Logical_Operator_out830_out1            : std_logic;
  SIGNAL Logical_Operator_out831_out1            : std_logic;
  SIGNAL Logical_Operator_out832_out1            : std_logic;
  SIGNAL Logical_Operator_out833_out1            : std_logic;
  SIGNAL Logical_Operator_out834_out1            : std_logic;
  SIGNAL Logical_Operator_out835_out1            : std_logic;
  SIGNAL Logical_Operator_out836_out1            : std_logic;
  SIGNAL Logical_Operator_out837_out1            : std_logic;
  SIGNAL Logical_Operator_out838_out1            : std_logic;
  SIGNAL Logical_Operator_out839_out1            : std_logic;
  SIGNAL Logical_Operator_out840_out1            : std_logic;
  SIGNAL Logical_Operator_out841_out1            : std_logic;
  SIGNAL Logical_Operator_out842_out1            : std_logic;
  SIGNAL Logical_Operator_out843_out1            : std_logic;
  SIGNAL Logical_Operator_out844_out1            : std_logic;
  SIGNAL Logical_Operator_out845_out1            : std_logic;
  SIGNAL Logical_Operator_out846_out1            : std_logic;
  SIGNAL Logical_Operator_out847_out1            : std_logic;
  SIGNAL Logical_Operator_out848_out1            : std_logic;
  SIGNAL Logical_Operator_out849_out1            : std_logic;
  SIGNAL Logical_Operator_out850_out1            : std_logic;
  SIGNAL Logical_Operator_out851_out1            : std_logic;
  SIGNAL Logical_Operator_out852_out1            : std_logic;
  SIGNAL Logical_Operator_out853_out1            : std_logic;
  SIGNAL Logical_Operator_out854_out1            : std_logic;
  SIGNAL Logical_Operator_out855_out1            : std_logic;
  SIGNAL Logical_Operator_out856_out1            : std_logic;
  SIGNAL Logical_Operator_out857_out1            : std_logic;
  SIGNAL Logical_Operator_out858_out1            : std_logic;
  SIGNAL Logical_Operator_out859_out1            : std_logic;
  SIGNAL Logical_Operator_out860_out1            : std_logic;
  SIGNAL Logical_Operator_out861_out1            : std_logic;
  SIGNAL Logical_Operator_out862_out1            : std_logic;
  SIGNAL Logical_Operator_out863_out1            : std_logic;
  SIGNAL Logical_Operator_out864_out1            : std_logic;
  SIGNAL Logical_Operator_out865_out1            : std_logic;
  SIGNAL Logical_Operator_out866_out1            : std_logic;
  SIGNAL Logical_Operator_out867_out1            : std_logic;
  SIGNAL Logical_Operator_out868_out1            : std_logic;
  SIGNAL Logical_Operator_out869_out1            : std_logic;
  SIGNAL Logical_Operator_out870_out1            : std_logic;
  SIGNAL Logical_Operator_out871_out1            : std_logic;
  SIGNAL Logical_Operator_out872_out1            : std_logic;
  SIGNAL Logical_Operator_out873_out1            : std_logic;
  SIGNAL Logical_Operator_out874_out1            : std_logic;
  SIGNAL Logical_Operator_out875_out1            : std_logic;
  SIGNAL Logical_Operator_out876_out1            : std_logic;
  SIGNAL Logical_Operator_out877_out1            : std_logic;
  SIGNAL Logical_Operator_out878_out1            : std_logic;
  SIGNAL Logical_Operator_out879_out1            : std_logic;
  SIGNAL Logical_Operator_out880_out1            : std_logic;
  SIGNAL Logical_Operator_out881_out1            : std_logic;
  SIGNAL Logical_Operator_out882_out1            : std_logic;
  SIGNAL Logical_Operator_out883_out1            : std_logic;
  SIGNAL Logical_Operator_out884_out1            : std_logic;
  SIGNAL Logical_Operator_out885_out1            : std_logic;
  SIGNAL Logical_Operator_out886_out1            : std_logic;
  SIGNAL Logical_Operator_out887_out1            : std_logic;
  SIGNAL Logical_Operator_out888_out1            : std_logic;
  SIGNAL Logical_Operator_out889_out1            : std_logic;
  SIGNAL Logical_Operator_out890_out1            : std_logic;
  SIGNAL Logical_Operator_out891_out1            : std_logic;
  SIGNAL Logical_Operator_out892_out1            : std_logic;
  SIGNAL Logical_Operator_out893_out1            : std_logic;
  SIGNAL Logical_Operator_out894_out1            : std_logic;
  SIGNAL Logical_Operator_out895_out1            : std_logic;
  SIGNAL Logical_Operator_out896_out1            : std_logic;
  SIGNAL Logical_Operator_out897_out1            : std_logic;
  SIGNAL Logical_Operator_out898_out1            : std_logic;
  SIGNAL Logical_Operator_out899_out1            : std_logic;
  SIGNAL Logical_Operator_out900_out1            : std_logic;
  SIGNAL Logical_Operator_out901_out1            : std_logic;
  SIGNAL Logical_Operator_out902_out1            : std_logic;
  SIGNAL Logical_Operator_out903_out1            : std_logic;
  SIGNAL Logical_Operator_out904_out1            : std_logic;
  SIGNAL Logical_Operator_out905_out1            : std_logic;
  SIGNAL Logical_Operator_out906_out1            : std_logic;
  SIGNAL Logical_Operator_out907_out1            : std_logic;
  SIGNAL Logical_Operator_out908_out1            : std_logic;
  SIGNAL Logical_Operator_out909_out1            : std_logic;
  SIGNAL Logical_Operator_out910_out1            : std_logic;
  SIGNAL Logical_Operator_out911_out1            : std_logic;
  SIGNAL Logical_Operator_out912_out1            : std_logic;
  SIGNAL Logical_Operator_out913_out1            : std_logic;
  SIGNAL Logical_Operator_out914_out1            : std_logic;
  SIGNAL Logical_Operator_out915_out1            : std_logic;
  SIGNAL Logical_Operator_out916_out1            : std_logic;
  SIGNAL Logical_Operator_out917_out1            : std_logic;
  SIGNAL Logical_Operator_out918_out1            : std_logic;
  SIGNAL Logical_Operator_out919_out1            : std_logic;
  SIGNAL Logical_Operator_out920_out1            : std_logic;
  SIGNAL Logical_Operator_out921_out1            : std_logic;
  SIGNAL Logical_Operator_out922_out1            : std_logic;
  SIGNAL Logical_Operator_out923_out1            : std_logic;
  SIGNAL Logical_Operator_out924_out1            : std_logic;
  SIGNAL Logical_Operator_out925_out1            : std_logic;
  SIGNAL Logical_Operator_out926_out1            : std_logic;
  SIGNAL Logical_Operator_out927_out1            : std_logic;
  SIGNAL Logical_Operator_out928_out1            : std_logic;
  SIGNAL Logical_Operator_out929_out1            : std_logic;
  SIGNAL Logical_Operator_out930_out1            : std_logic;
  SIGNAL Logical_Operator_out931_out1            : std_logic;
  SIGNAL Logical_Operator_out932_out1            : std_logic;
  SIGNAL Logical_Operator_out933_out1            : std_logic;
  SIGNAL Logical_Operator_out934_out1            : std_logic;
  SIGNAL Logical_Operator_out935_out1            : std_logic;
  SIGNAL Logical_Operator_out936_out1            : std_logic;
  SIGNAL Logical_Operator_out937_out1            : std_logic;
  SIGNAL Logical_Operator_out938_out1            : std_logic;
  SIGNAL Logical_Operator_out939_out1            : std_logic;
  SIGNAL Logical_Operator_out940_out1            : std_logic;
  SIGNAL Logical_Operator_out941_out1            : std_logic;
  SIGNAL Logical_Operator_out942_out1            : std_logic;
  SIGNAL Logical_Operator_out943_out1            : std_logic;
  SIGNAL Logical_Operator_out944_out1            : std_logic;
  SIGNAL Logical_Operator_out945_out1            : std_logic;
  SIGNAL Logical_Operator_out946_out1            : std_logic;
  SIGNAL Logical_Operator_out947_out1            : std_logic;
  SIGNAL Logical_Operator_out948_out1            : std_logic;
  SIGNAL Logical_Operator_out949_out1            : std_logic;
  SIGNAL Logical_Operator_out950_out1            : std_logic;
  SIGNAL Logical_Operator_out951_out1            : std_logic;
  SIGNAL Logical_Operator_out952_out1            : std_logic;
  SIGNAL Logical_Operator_out953_out1            : std_logic;
  SIGNAL Logical_Operator_out954_out1            : std_logic;
  SIGNAL Logical_Operator_out955_out1            : std_logic;
  SIGNAL Logical_Operator_out956_out1            : std_logic;
  SIGNAL Logical_Operator_out957_out1            : std_logic;
  SIGNAL Logical_Operator_out958_out1            : std_logic;
  SIGNAL Logical_Operator_out959_out1            : std_logic;
  SIGNAL Logical_Operator_out960_out1            : std_logic;
  SIGNAL Logical_Operator_out961_out1            : std_logic;
  SIGNAL Logical_Operator_out962_out1            : std_logic;
  SIGNAL Logical_Operator_out963_out1            : std_logic;
  SIGNAL Logical_Operator_out964_out1            : std_logic;
  SIGNAL Logical_Operator_out965_out1            : std_logic;
  SIGNAL Logical_Operator_out966_out1            : std_logic;
  SIGNAL Logical_Operator_out967_out1            : std_logic;
  SIGNAL Logical_Operator_out968_out1            : std_logic;
  SIGNAL Logical_Operator_out969_out1            : std_logic;
  SIGNAL Logical_Operator_out970_out1            : std_logic;
  SIGNAL Logical_Operator_out971_out1            : std_logic;
  SIGNAL Logical_Operator_out972_out1            : std_logic;
  SIGNAL Logical_Operator_out973_out1            : std_logic;
  SIGNAL Logical_Operator_out974_out1            : std_logic;
  SIGNAL Logical_Operator_out975_out1            : std_logic;
  SIGNAL Logical_Operator_out976_out1            : std_logic;
  SIGNAL Logical_Operator_out977_out1            : std_logic;
  SIGNAL Logical_Operator_out978_out1            : std_logic;
  SIGNAL Logical_Operator_out979_out1            : std_logic;
  SIGNAL Logical_Operator_out980_out1            : std_logic;
  SIGNAL Logical_Operator_out981_out1            : std_logic;
  SIGNAL Logical_Operator_out982_out1            : std_logic;
  SIGNAL Logical_Operator_out983_out1            : std_logic;
  SIGNAL Logical_Operator_out984_out1            : std_logic;
  SIGNAL Logical_Operator_out985_out1            : std_logic;
  SIGNAL Logical_Operator_out986_out1            : std_logic;
  SIGNAL Logical_Operator_out987_out1            : std_logic;
  SIGNAL Logical_Operator_out988_out1            : std_logic;
  SIGNAL Logical_Operator_out989_out1            : std_logic;
  SIGNAL Logical_Operator_out990_out1            : std_logic;
  SIGNAL Logical_Operator_out991_out1            : std_logic;
  SIGNAL Logical_Operator_out992_out1            : std_logic;
  SIGNAL Logical_Operator_out993_out1            : std_logic;
  SIGNAL Logical_Operator_out994_out1            : std_logic;
  SIGNAL Logical_Operator_out995_out1            : std_logic;
  SIGNAL Logical_Operator_out996_out1            : std_logic;
  SIGNAL Logical_Operator_out997_out1            : std_logic;
  SIGNAL Logical_Operator_out998_out1            : std_logic;
  SIGNAL Logical_Operator_out999_out1            : std_logic;
  SIGNAL Logical_Operator_out1000_out1            : std_logic;
  SIGNAL Logical_Operator_out1001_out1            : std_logic;
  SIGNAL Logical_Operator_out1002_out1            : std_logic;
  SIGNAL Logical_Operator_out1003_out1            : std_logic;
  SIGNAL Logical_Operator_out1004_out1            : std_logic;
  SIGNAL Logical_Operator_out1005_out1            : std_logic;
  SIGNAL Logical_Operator_out1006_out1            : std_logic;
  SIGNAL Logical_Operator_out1007_out1            : std_logic;
  SIGNAL Logical_Operator_out1008_out1            : std_logic;
  SIGNAL Logical_Operator_out1009_out1            : std_logic;
  SIGNAL Logical_Operator_out1010_out1            : std_logic;
  SIGNAL Logical_Operator_out1011_out1            : std_logic;
  SIGNAL Logical_Operator_out1012_out1            : std_logic;
  SIGNAL Logical_Operator_out1013_out1            : std_logic;
  SIGNAL Logical_Operator_out1014_out1            : std_logic;
  SIGNAL Logical_Operator_out1015_out1            : std_logic;
  SIGNAL Logical_Operator_out1016_out1            : std_logic;
  SIGNAL Logical_Operator_out1017_out1            : std_logic;
  SIGNAL Logical_Operator_out1018_out1            : std_logic;
  SIGNAL Logical_Operator_out1019_out1            : std_logic;
  SIGNAL Logical_Operator_out1020_out1            : std_logic;
  SIGNAL Logical_Operator_out1021_out1            : std_logic;
  SIGNAL Logical_Operator_out1022_out1            : std_logic;
  SIGNAL Logical_Operator_out1023_out1            : std_logic;
  SIGNAL Logical_Operator_out1024_out1            : std_logic;
  SIGNAL Logical_Operator_out1025_out1            : std_logic;
  SIGNAL Logical_Operator_out1026_out1            : std_logic;
  SIGNAL Logical_Operator_out1027_out1            : std_logic;
  SIGNAL Logical_Operator_out1028_out1            : std_logic;
  SIGNAL Logical_Operator_out1029_out1            : std_logic;
  SIGNAL Logical_Operator_out1030_out1            : std_logic;
  SIGNAL Logical_Operator_out1031_out1            : std_logic;
  SIGNAL Logical_Operator_out1032_out1            : std_logic;
  SIGNAL Logical_Operator_out1033_out1            : std_logic;
  SIGNAL Logical_Operator_out1034_out1            : std_logic;
  SIGNAL Logical_Operator_out1035_out1            : std_logic;
  SIGNAL Logical_Operator_out1036_out1            : std_logic;
  SIGNAL Logical_Operator_out1037_out1            : std_logic;
  SIGNAL Logical_Operator_out1038_out1            : std_logic;
  SIGNAL Logical_Operator_out1039_out1            : std_logic;
  SIGNAL Logical_Operator_out1040_out1            : std_logic;
  SIGNAL Logical_Operator_out1041_out1            : std_logic;
  SIGNAL Logical_Operator_out1042_out1            : std_logic;
  SIGNAL Logical_Operator_out1043_out1            : std_logic;
  SIGNAL Logical_Operator_out1044_out1            : std_logic;
  SIGNAL Logical_Operator_out1045_out1            : std_logic;
  SIGNAL Logical_Operator_out1046_out1            : std_logic;
  SIGNAL Logical_Operator_out1047_out1            : std_logic;
  SIGNAL Logical_Operator_out1048_out1            : std_logic;
  SIGNAL Logical_Operator_out1049_out1            : std_logic;
  SIGNAL Logical_Operator_out1050_out1            : std_logic;
  SIGNAL Logical_Operator_out1051_out1            : std_logic;
  SIGNAL Logical_Operator_out1052_out1            : std_logic;
  SIGNAL Logical_Operator_out1053_out1            : std_logic;
  SIGNAL Logical_Operator_out1054_out1            : std_logic;
  SIGNAL Logical_Operator_out1055_out1            : std_logic;
  SIGNAL Logical_Operator_out1056_out1            : std_logic;
  SIGNAL Logical_Operator_out1057_out1            : std_logic;
  SIGNAL Logical_Operator_out1058_out1            : std_logic;
  SIGNAL Logical_Operator_out1059_out1            : std_logic;
  SIGNAL Logical_Operator_out1060_out1            : std_logic;
  SIGNAL Logical_Operator_out1061_out1            : std_logic;
  SIGNAL Logical_Operator_out1062_out1            : std_logic;
  SIGNAL Logical_Operator_out1063_out1            : std_logic;
  SIGNAL Logical_Operator_out1064_out1            : std_logic;
  SIGNAL Logical_Operator_out1065_out1            : std_logic;
  SIGNAL Logical_Operator_out1066_out1            : std_logic;
  SIGNAL Logical_Operator_out1067_out1            : std_logic;
  SIGNAL Logical_Operator_out1068_out1            : std_logic;
  SIGNAL Logical_Operator_out1069_out1            : std_logic;
  SIGNAL Logical_Operator_out1070_out1            : std_logic;
  SIGNAL Logical_Operator_out1071_out1            : std_logic;
  SIGNAL Logical_Operator_out1072_out1            : std_logic;
  SIGNAL Logical_Operator_out1073_out1            : std_logic;
  SIGNAL Logical_Operator_out1074_out1            : std_logic;
  SIGNAL Logical_Operator_out1075_out1            : std_logic;
  SIGNAL Logical_Operator_out1076_out1            : std_logic;
  SIGNAL Logical_Operator_out1077_out1            : std_logic;
  SIGNAL Logical_Operator_out1078_out1            : std_logic;
  SIGNAL Logical_Operator_out1079_out1            : std_logic;
  SIGNAL Logical_Operator_out1080_out1            : std_logic;
  SIGNAL Logical_Operator_out1081_out1            : std_logic;
  SIGNAL Logical_Operator_out1082_out1            : std_logic;
  SIGNAL Logical_Operator_out1083_out1            : std_logic;
  SIGNAL Logical_Operator_out1084_out1            : std_logic;
  SIGNAL Logical_Operator_out1085_out1            : std_logic;
  SIGNAL Logical_Operator_out1086_out1            : std_logic;
  SIGNAL Logical_Operator_out1087_out1            : std_logic;
  SIGNAL Logical_Operator_out1088_out1            : std_logic;
  SIGNAL Logical_Operator_out1089_out1            : std_logic;
  SIGNAL Logical_Operator_out1090_out1            : std_logic;
  SIGNAL Logical_Operator_out1091_out1            : std_logic;
  SIGNAL Logical_Operator_out1092_out1            : std_logic;
  SIGNAL Logical_Operator_out1093_out1            : std_logic;
  SIGNAL Logical_Operator_out1094_out1            : std_logic;
  SIGNAL Logical_Operator_out1095_out1            : std_logic;
  SIGNAL Logical_Operator_out1096_out1            : std_logic;
  SIGNAL Logical_Operator_out1097_out1            : std_logic;
  SIGNAL Logical_Operator_out1098_out1            : std_logic;
  SIGNAL Logical_Operator_out1099_out1            : std_logic;
  SIGNAL Logical_Operator_out1100_out1            : std_logic;
  SIGNAL Logical_Operator_out1101_out1            : std_logic;
  SIGNAL Logical_Operator_out1102_out1            : std_logic;
  SIGNAL Logical_Operator_out1103_out1            : std_logic;
  SIGNAL Logical_Operator_out1104_out1            : std_logic;
  SIGNAL Logical_Operator_out1105_out1            : std_logic;
  SIGNAL Logical_Operator_out1106_out1            : std_logic;
  SIGNAL Logical_Operator_out1107_out1            : std_logic;
  SIGNAL Logical_Operator_out1108_out1            : std_logic;
  SIGNAL Logical_Operator_out1109_out1            : std_logic;
  SIGNAL Logical_Operator_out1110_out1            : std_logic;
  SIGNAL Logical_Operator_out1111_out1            : std_logic;
  SIGNAL Logical_Operator_out1112_out1            : std_logic;
  SIGNAL Logical_Operator_out1113_out1            : std_logic;
  SIGNAL Logical_Operator_out1114_out1            : std_logic;
  SIGNAL Logical_Operator_out1115_out1            : std_logic;
  SIGNAL Logical_Operator_out1116_out1            : std_logic;
  SIGNAL Logical_Operator_out1117_out1            : std_logic;
  SIGNAL Logical_Operator_out1118_out1            : std_logic;
  SIGNAL Logical_Operator_out1119_out1            : std_logic;
  SIGNAL Logical_Operator_out1120_out1            : std_logic;
  SIGNAL Logical_Operator_out1121_out1            : std_logic;
  SIGNAL Logical_Operator_out1122_out1            : std_logic;
  SIGNAL Logical_Operator_out1123_out1            : std_logic;
  SIGNAL Logical_Operator_out1124_out1            : std_logic;
  SIGNAL Logical_Operator_out1125_out1            : std_logic;
  SIGNAL Logical_Operator_out1126_out1            : std_logic;
  SIGNAL Logical_Operator_out1127_out1            : std_logic;
  SIGNAL Logical_Operator_out1128_out1            : std_logic;
  SIGNAL Logical_Operator_out1129_out1            : std_logic;
  SIGNAL Logical_Operator_out1130_out1            : std_logic;
  SIGNAL Logical_Operator_out1131_out1            : std_logic;
  SIGNAL Logical_Operator_out1132_out1            : std_logic;
  SIGNAL Logical_Operator_out1133_out1            : std_logic;
  SIGNAL Logical_Operator_out1134_out1            : std_logic;
  SIGNAL Logical_Operator_out1135_out1            : std_logic;
  SIGNAL Logical_Operator_out1136_out1            : std_logic;
  SIGNAL Logical_Operator_out1137_out1            : std_logic;
  SIGNAL Logical_Operator_out1138_out1            : std_logic;
  SIGNAL Logical_Operator_out1139_out1            : std_logic;
  SIGNAL Logical_Operator_out1140_out1            : std_logic;
  SIGNAL Logical_Operator_out1141_out1            : std_logic;
  SIGNAL Logical_Operator_out1142_out1            : std_logic;
  SIGNAL Logical_Operator_out1143_out1            : std_logic;
  SIGNAL Logical_Operator_out1144_out1            : std_logic;
  SIGNAL Logical_Operator_out1145_out1            : std_logic;
  SIGNAL Logical_Operator_out1146_out1            : std_logic;
  SIGNAL Logical_Operator_out1147_out1            : std_logic;
  SIGNAL Logical_Operator_out1148_out1            : std_logic;
  SIGNAL Logical_Operator_out1149_out1            : std_logic;
  SIGNAL Logical_Operator_out1150_out1            : std_logic;
  SIGNAL Logical_Operator_out1151_out1            : std_logic;
  SIGNAL Logical_Operator_out1152_out1            : std_logic;
  SIGNAL Logical_Operator_out1153_out1            : std_logic;
  SIGNAL Logical_Operator_out1154_out1            : std_logic;
  SIGNAL Logical_Operator_out1155_out1            : std_logic;
  SIGNAL Logical_Operator_out1156_out1            : std_logic;
  SIGNAL Logical_Operator_out1157_out1            : std_logic;
  SIGNAL Logical_Operator_out1158_out1            : std_logic;
  SIGNAL Logical_Operator_out1159_out1            : std_logic;
  SIGNAL Logical_Operator_out1160_out1            : std_logic;
  SIGNAL Logical_Operator_out1161_out1            : std_logic;
  SIGNAL Logical_Operator_out1162_out1            : std_logic;
  SIGNAL Logical_Operator_out1163_out1            : std_logic;
  SIGNAL Logical_Operator_out1164_out1            : std_logic;
  SIGNAL Logical_Operator_out1165_out1            : std_logic;
  SIGNAL Logical_Operator_out1166_out1            : std_logic;
  SIGNAL Logical_Operator_out1167_out1            : std_logic;
  SIGNAL Logical_Operator_out1168_out1            : std_logic;
  SIGNAL Logical_Operator_out1169_out1            : std_logic;
  SIGNAL Logical_Operator_out1170_out1            : std_logic;
  SIGNAL Logical_Operator_out1171_out1            : std_logic;
  SIGNAL Logical_Operator_out1172_out1            : std_logic;
  SIGNAL Logical_Operator_out1173_out1            : std_logic;
  SIGNAL Logical_Operator_out1174_out1            : std_logic;
  SIGNAL Logical_Operator_out1175_out1            : std_logic;
  SIGNAL Logical_Operator_out1176_out1            : std_logic;
  SIGNAL Logical_Operator_out1177_out1            : std_logic;
  SIGNAL Logical_Operator_out1178_out1            : std_logic;
  SIGNAL Logical_Operator_out1179_out1            : std_logic;
  SIGNAL Logical_Operator_out1180_out1            : std_logic;
  SIGNAL Logical_Operator_out1181_out1            : std_logic;
  SIGNAL Logical_Operator_out1182_out1            : std_logic;
  SIGNAL Logical_Operator_out1183_out1            : std_logic;
  SIGNAL Logical_Operator_out1184_out1            : std_logic;
  SIGNAL Logical_Operator_out1185_out1            : std_logic;
  SIGNAL Logical_Operator_out1186_out1            : std_logic;
  SIGNAL Logical_Operator_out1187_out1            : std_logic;
  SIGNAL Logical_Operator_out1188_out1            : std_logic;
  SIGNAL Logical_Operator_out1189_out1            : std_logic;
  SIGNAL Logical_Operator_out1190_out1            : std_logic;
  SIGNAL Logical_Operator_out1191_out1            : std_logic;
  SIGNAL Logical_Operator_out1192_out1            : std_logic;
  SIGNAL Logical_Operator_out1193_out1            : std_logic;
  SIGNAL Logical_Operator_out1194_out1            : std_logic;
  SIGNAL Logical_Operator_out1195_out1            : std_logic;
  SIGNAL Logical_Operator_out1196_out1            : std_logic;
  SIGNAL Logical_Operator_out1197_out1            : std_logic;
  SIGNAL Logical_Operator_out1198_out1            : std_logic;
  SIGNAL Logical_Operator_out1199_out1            : std_logic;
  SIGNAL Logical_Operator_out1200_out1            : std_logic;
  SIGNAL Logical_Operator_out1201_out1            : std_logic;
  SIGNAL Logical_Operator_out1202_out1            : std_logic;
  SIGNAL Logical_Operator_out1203_out1            : std_logic;
  SIGNAL Logical_Operator_out1204_out1            : std_logic;
  SIGNAL Logical_Operator_out1205_out1            : std_logic;
  SIGNAL Logical_Operator_out1206_out1            : std_logic;
  SIGNAL Logical_Operator_out1207_out1            : std_logic;
  SIGNAL Logical_Operator_out1208_out1            : std_logic;
  SIGNAL Logical_Operator_out1209_out1            : std_logic;
  SIGNAL Logical_Operator_out1210_out1            : std_logic;
  SIGNAL Logical_Operator_out1211_out1            : std_logic;
  SIGNAL Logical_Operator_out1212_out1            : std_logic;
  SIGNAL Logical_Operator_out1213_out1            : std_logic;
  SIGNAL Logical_Operator_out1214_out1            : std_logic;
  SIGNAL Logical_Operator_out1215_out1            : std_logic;
  SIGNAL Logical_Operator_out1216_out1            : std_logic;
  SIGNAL Logical_Operator_out1217_out1            : std_logic;
  SIGNAL Logical_Operator_out1218_out1            : std_logic;
  SIGNAL Logical_Operator_out1219_out1            : std_logic;
  SIGNAL Logical_Operator_out1220_out1            : std_logic;
  SIGNAL Logical_Operator_out1221_out1            : std_logic;
  SIGNAL Logical_Operator_out1222_out1            : std_logic;
  SIGNAL Logical_Operator_out1223_out1            : std_logic;
  SIGNAL Logical_Operator_out1224_out1            : std_logic;
  SIGNAL Logical_Operator_out1225_out1            : std_logic;
  SIGNAL Logical_Operator_out1226_out1            : std_logic;
  SIGNAL Logical_Operator_out1227_out1            : std_logic;
  SIGNAL Logical_Operator_out1228_out1            : std_logic;
  SIGNAL Logical_Operator_out1229_out1            : std_logic;
  SIGNAL Logical_Operator_out1230_out1            : std_logic;
  SIGNAL Logical_Operator_out1231_out1            : std_logic;
  SIGNAL Logical_Operator_out1232_out1            : std_logic;
  SIGNAL Logical_Operator_out1233_out1            : std_logic;
  SIGNAL Logical_Operator_out1234_out1            : std_logic;
  SIGNAL Logical_Operator_out1235_out1            : std_logic;
  SIGNAL Logical_Operator_out1236_out1            : std_logic;
  SIGNAL Logical_Operator_out1237_out1            : std_logic;
  SIGNAL Logical_Operator_out1238_out1            : std_logic;
  SIGNAL Logical_Operator_out1239_out1            : std_logic;
  SIGNAL Logical_Operator_out1240_out1            : std_logic;
  SIGNAL Logical_Operator_out1241_out1            : std_logic;
  SIGNAL Logical_Operator_out1242_out1            : std_logic;
  SIGNAL Logical_Operator_out1243_out1            : std_logic;
  SIGNAL Logical_Operator_out1244_out1            : std_logic;
  SIGNAL Logical_Operator_out1245_out1            : std_logic;
  SIGNAL Logical_Operator_out1246_out1            : std_logic;
  SIGNAL Logical_Operator_out1247_out1            : std_logic;
  SIGNAL Logical_Operator_out1248_out1            : std_logic;
  SIGNAL Logical_Operator_out1249_out1            : std_logic;
  SIGNAL Logical_Operator_out1250_out1            : std_logic;
  SIGNAL Logical_Operator_out1251_out1            : std_logic;
  SIGNAL Logical_Operator_out1252_out1            : std_logic;
  SIGNAL Logical_Operator_out1253_out1            : std_logic;
  SIGNAL Logical_Operator_out1254_out1            : std_logic;
  SIGNAL Logical_Operator_out1255_out1            : std_logic;
  SIGNAL Logical_Operator_out1256_out1            : std_logic;
  SIGNAL Logical_Operator_out1257_out1            : std_logic;
  SIGNAL Logical_Operator_out1258_out1            : std_logic;
  SIGNAL Logical_Operator_out1259_out1            : std_logic;
  SIGNAL Logical_Operator_out1260_out1            : std_logic;
  SIGNAL Logical_Operator_out1261_out1            : std_logic;
  SIGNAL Logical_Operator_out1262_out1            : std_logic;
  SIGNAL Logical_Operator_out1263_out1            : std_logic;
  SIGNAL Logical_Operator_out1264_out1            : std_logic;
  SIGNAL Logical_Operator_out1265_out1            : std_logic;
  SIGNAL Logical_Operator_out1266_out1            : std_logic;
  SIGNAL Logical_Operator_out1267_out1            : std_logic;
  SIGNAL Logical_Operator_out1268_out1            : std_logic;
  SIGNAL Logical_Operator_out1269_out1            : std_logic;
  SIGNAL Logical_Operator_out1270_out1            : std_logic;
  SIGNAL Logical_Operator_out1271_out1            : std_logic;
  SIGNAL Logical_Operator_out1272_out1            : std_logic;
  SIGNAL Logical_Operator_out1273_out1            : std_logic;
  SIGNAL Logical_Operator_out1274_out1            : std_logic;
  SIGNAL Logical_Operator_out1275_out1            : std_logic;
  SIGNAL Logical_Operator_out1276_out1            : std_logic;
  SIGNAL Logical_Operator_out1277_out1            : std_logic;
  SIGNAL Logical_Operator_out1278_out1            : std_logic;
  SIGNAL Logical_Operator_out1279_out1            : std_logic;
  SIGNAL Logical_Operator_out1280_out1            : std_logic;
  SIGNAL Logical_Operator_out1281_out1            : std_logic;
  SIGNAL Logical_Operator_out1282_out1            : std_logic;
  SIGNAL Logical_Operator_out1283_out1            : std_logic;
  SIGNAL Logical_Operator_out1284_out1            : std_logic;
  SIGNAL Logical_Operator_out1285_out1            : std_logic;
  SIGNAL Logical_Operator_out1286_out1            : std_logic;
  SIGNAL Logical_Operator_out1287_out1            : std_logic;
  SIGNAL Logical_Operator_out1288_out1            : std_logic;
  SIGNAL Logical_Operator_out1289_out1            : std_logic;
  SIGNAL Logical_Operator_out1290_out1            : std_logic;
  SIGNAL Logical_Operator_out1291_out1            : std_logic;
  SIGNAL Logical_Operator_out1292_out1            : std_logic;
  SIGNAL Logical_Operator_out1293_out1            : std_logic;
  SIGNAL Logical_Operator_out1294_out1            : std_logic;
  SIGNAL Logical_Operator_out1295_out1            : std_logic;
  SIGNAL Logical_Operator_out1296_out1            : std_logic;
  SIGNAL Logical_Operator_out1297_out1            : std_logic;
  SIGNAL Logical_Operator_out1298_out1            : std_logic;
  SIGNAL Logical_Operator_out1299_out1            : std_logic;
  SIGNAL Logical_Operator_out1300_out1            : std_logic;
  SIGNAL Logical_Operator_out1301_out1            : std_logic;
  SIGNAL Logical_Operator_out1302_out1            : std_logic;
  SIGNAL Logical_Operator_out1303_out1            : std_logic;
  SIGNAL Logical_Operator_out1304_out1            : std_logic;
  SIGNAL Logical_Operator_out1305_out1            : std_logic;
  SIGNAL Logical_Operator_out1306_out1            : std_logic;
  SIGNAL Logical_Operator_out1307_out1            : std_logic;
  SIGNAL Logical_Operator_out1308_out1            : std_logic;
  SIGNAL Logical_Operator_out1309_out1            : std_logic;
  SIGNAL Logical_Operator_out1310_out1            : std_logic;
  SIGNAL Logical_Operator_out1311_out1            : std_logic;
  SIGNAL Logical_Operator_out1312_out1            : std_logic;
  SIGNAL Logical_Operator_out1313_out1            : std_logic;
  SIGNAL Logical_Operator_out1314_out1            : std_logic;
  SIGNAL Logical_Operator_out1315_out1            : std_logic;
  SIGNAL Logical_Operator_out1316_out1            : std_logic;
  SIGNAL Logical_Operator_out1317_out1            : std_logic;
  SIGNAL Logical_Operator_out1318_out1            : std_logic;
  SIGNAL Logical_Operator_out1319_out1            : std_logic;
  SIGNAL Logical_Operator_out1320_out1            : std_logic;
  SIGNAL Logical_Operator_out1321_out1            : std_logic;
  SIGNAL Logical_Operator_out1322_out1            : std_logic;
  SIGNAL Logical_Operator_out1323_out1            : std_logic;
  SIGNAL Logical_Operator_out1324_out1            : std_logic;
  SIGNAL Logical_Operator_out1325_out1            : std_logic;
  SIGNAL Logical_Operator_out1326_out1            : std_logic;
  SIGNAL Logical_Operator_out1327_out1            : std_logic;
  SIGNAL Logical_Operator_out1328_out1            : std_logic;
  SIGNAL Logical_Operator_out1329_out1            : std_logic;
  SIGNAL Logical_Operator_out1330_out1            : std_logic;
  SIGNAL Logical_Operator_out1331_out1            : std_logic;
  SIGNAL Logical_Operator_out1332_out1            : std_logic;
  SIGNAL Logical_Operator_out1333_out1            : std_logic;
  SIGNAL Logical_Operator_out1334_out1            : std_logic;
  SIGNAL Logical_Operator_out1335_out1            : std_logic;
  SIGNAL Logical_Operator_out1336_out1            : std_logic;
  SIGNAL Logical_Operator_out1337_out1            : std_logic;
  SIGNAL Logical_Operator_out1338_out1            : std_logic;
  SIGNAL Logical_Operator_out1339_out1            : std_logic;
  SIGNAL Logical_Operator_out1340_out1            : std_logic;
  SIGNAL Logical_Operator_out1341_out1            : std_logic;
  SIGNAL Logical_Operator_out1342_out1            : std_logic;
  SIGNAL Logical_Operator_out1343_out1            : std_logic;
  SIGNAL Logical_Operator_out1344_out1            : std_logic;
  SIGNAL Logical_Operator_out1345_out1            : std_logic;
  SIGNAL Logical_Operator_out1346_out1            : std_logic;
  SIGNAL Logical_Operator_out1347_out1            : std_logic;
  SIGNAL Logical_Operator_out1348_out1            : std_logic;
  SIGNAL Logical_Operator_out1349_out1            : std_logic;
  SIGNAL Logical_Operator_out1350_out1            : std_logic;
  SIGNAL Logical_Operator_out1351_out1            : std_logic;
  SIGNAL Logical_Operator_out1352_out1            : std_logic;
  SIGNAL Logical_Operator_out1353_out1            : std_logic;
  SIGNAL Logical_Operator_out1354_out1            : std_logic;
  SIGNAL Logical_Operator_out1355_out1            : std_logic;
  SIGNAL Logical_Operator_out1356_out1            : std_logic;
  SIGNAL Logical_Operator_out1357_out1            : std_logic;
  SIGNAL Logical_Operator_out1358_out1            : std_logic;
  SIGNAL Logical_Operator_out1359_out1            : std_logic;
  SIGNAL Logical_Operator_out1360_out1            : std_logic;
  SIGNAL Logical_Operator_out1361_out1            : std_logic;
  SIGNAL Logical_Operator_out1362_out1            : std_logic;
  SIGNAL Logical_Operator_out1363_out1            : std_logic;
  SIGNAL Logical_Operator_out1364_out1            : std_logic;
  SIGNAL Logical_Operator_out1365_out1            : std_logic;
  SIGNAL Logical_Operator_out1366_out1            : std_logic;
  SIGNAL Logical_Operator_out1367_out1            : std_logic;
  SIGNAL Logical_Operator_out1368_out1            : std_logic;
  SIGNAL Logical_Operator_out1369_out1            : std_logic;
  SIGNAL Logical_Operator_out1370_out1            : std_logic;
  SIGNAL Logical_Operator_out1371_out1            : std_logic;
  SIGNAL Logical_Operator_out1372_out1            : std_logic;
  SIGNAL Logical_Operator_out1373_out1            : std_logic;
  SIGNAL Logical_Operator_out1374_out1            : std_logic;
  SIGNAL Logical_Operator_out1375_out1            : std_logic;
  SIGNAL Logical_Operator_out1376_out1            : std_logic;
  SIGNAL Logical_Operator_out1377_out1            : std_logic;
  SIGNAL Logical_Operator_out1378_out1            : std_logic;
  SIGNAL Logical_Operator_out1379_out1            : std_logic;
  SIGNAL Logical_Operator_out1380_out1            : std_logic;
  SIGNAL Logical_Operator_out1381_out1            : std_logic;
  SIGNAL Logical_Operator_out1382_out1            : std_logic;
  SIGNAL Logical_Operator_out1383_out1            : std_logic;
  SIGNAL Logical_Operator_out1384_out1            : std_logic;
  SIGNAL Logical_Operator_out1385_out1            : std_logic;
  SIGNAL Logical_Operator_out1386_out1            : std_logic;
  SIGNAL Logical_Operator_out1387_out1            : std_logic;
  SIGNAL Logical_Operator_out1388_out1            : std_logic;
  SIGNAL Logical_Operator_out1389_out1            : std_logic;
  SIGNAL Logical_Operator_out1390_out1            : std_logic;
  SIGNAL Logical_Operator_out1391_out1            : std_logic;
  SIGNAL Logical_Operator_out1392_out1            : std_logic;
  SIGNAL Logical_Operator_out1393_out1            : std_logic;
  SIGNAL Logical_Operator_out1394_out1            : std_logic;
  SIGNAL Logical_Operator_out1395_out1            : std_logic;
  SIGNAL Logical_Operator_out1396_out1            : std_logic;
  SIGNAL Logical_Operator_out1397_out1            : std_logic;
  SIGNAL Logical_Operator_out1398_out1            : std_logic;
  SIGNAL Logical_Operator_out1399_out1            : std_logic;
  SIGNAL Logical_Operator_out1400_out1            : std_logic;
  SIGNAL Logical_Operator_out1401_out1            : std_logic;
  SIGNAL Logical_Operator_out1402_out1            : std_logic;
  SIGNAL Logical_Operator_out1403_out1            : std_logic;
  SIGNAL Logical_Operator_out1404_out1            : std_logic;
  SIGNAL Logical_Operator_out1405_out1            : std_logic;
  SIGNAL Logical_Operator_out1406_out1            : std_logic;
  SIGNAL Logical_Operator_out1407_out1            : std_logic;
  SIGNAL Logical_Operator_out1408_out1            : std_logic;
  SIGNAL Logical_Operator_out1409_out1            : std_logic;
  SIGNAL Logical_Operator_out1410_out1            : std_logic;
  SIGNAL Logical_Operator_out1411_out1            : std_logic;
  SIGNAL Logical_Operator_out1412_out1            : std_logic;
  SIGNAL Logical_Operator_out1413_out1            : std_logic;
  SIGNAL Logical_Operator_out1414_out1            : std_logic;
  SIGNAL Logical_Operator_out1415_out1            : std_logic;
  SIGNAL Logical_Operator_out1416_out1            : std_logic;
  SIGNAL Logical_Operator_out1417_out1            : std_logic;
  SIGNAL Logical_Operator_out1418_out1            : std_logic;
  SIGNAL Logical_Operator_out1419_out1            : std_logic;
  SIGNAL Logical_Operator_out1420_out1            : std_logic;
  SIGNAL Logical_Operator_out1421_out1            : std_logic;
  SIGNAL Logical_Operator_out1422_out1            : std_logic;
  SIGNAL Logical_Operator_out1423_out1            : std_logic;
  SIGNAL Logical_Operator_out1424_out1            : std_logic;
  SIGNAL Logical_Operator_out1425_out1            : std_logic;
  SIGNAL Logical_Operator_out1426_out1            : std_logic;
  SIGNAL Logical_Operator_out1427_out1            : std_logic;
  SIGNAL Logical_Operator_out1428_out1            : std_logic;
  SIGNAL Logical_Operator_out1429_out1            : std_logic;
  SIGNAL Logical_Operator_out1430_out1            : std_logic;
  SIGNAL Logical_Operator_out1431_out1            : std_logic;
  SIGNAL Logical_Operator_out1432_out1            : std_logic;
  SIGNAL Logical_Operator_out1433_out1            : std_logic;
  SIGNAL Logical_Operator_out1434_out1            : std_logic;
  SIGNAL Logical_Operator_out1435_out1            : std_logic;
  SIGNAL Logical_Operator_out1436_out1            : std_logic;
  SIGNAL Logical_Operator_out1437_out1            : std_logic;
  SIGNAL Logical_Operator_out1438_out1            : std_logic;
  SIGNAL Logical_Operator_out1439_out1            : std_logic;
  SIGNAL Logical_Operator_out1440_out1            : std_logic;
  SIGNAL Logical_Operator_out1441_out1            : std_logic;
  SIGNAL Logical_Operator_out1442_out1            : std_logic;
  SIGNAL Logical_Operator_out1443_out1            : std_logic;
  SIGNAL Logical_Operator_out1444_out1            : std_logic;
  SIGNAL Logical_Operator_out1445_out1            : std_logic;
  SIGNAL Logical_Operator_out1446_out1            : std_logic;
  SIGNAL Logical_Operator_out1447_out1            : std_logic;
  SIGNAL Logical_Operator_out1448_out1            : std_logic;
  SIGNAL Logical_Operator_out1449_out1            : std_logic;
  SIGNAL Logical_Operator_out1450_out1            : std_logic;
  SIGNAL Logical_Operator_out1451_out1            : std_logic;
  SIGNAL Logical_Operator_out1452_out1            : std_logic;
  SIGNAL Logical_Operator_out1453_out1            : std_logic;
  SIGNAL Logical_Operator_out1454_out1            : std_logic;
  SIGNAL Logical_Operator_out1455_out1            : std_logic;
  SIGNAL Logical_Operator_out1456_out1            : std_logic;
  SIGNAL Logical_Operator_out1457_out1            : std_logic;
  SIGNAL Logical_Operator_out1458_out1            : std_logic;
  SIGNAL Logical_Operator_out1459_out1            : std_logic;
  SIGNAL Logical_Operator_out1460_out1            : std_logic;
  SIGNAL Logical_Operator_out1461_out1            : std_logic;
  SIGNAL Logical_Operator_out1462_out1            : std_logic;
  SIGNAL Logical_Operator_out1463_out1            : std_logic;
  SIGNAL Logical_Operator_out1464_out1            : std_logic;
  SIGNAL Logical_Operator_out1465_out1            : std_logic;
  SIGNAL Logical_Operator_out1466_out1            : std_logic;
  SIGNAL Logical_Operator_out1467_out1            : std_logic;
  SIGNAL Logical_Operator_out1468_out1            : std_logic;
  SIGNAL Logical_Operator_out1469_out1            : std_logic;
  SIGNAL Logical_Operator_out1470_out1            : std_logic;
  SIGNAL Logical_Operator_out1471_out1            : std_logic;
  SIGNAL Logical_Operator_out1472_out1            : std_logic;
  SIGNAL Logical_Operator_out1473_out1            : std_logic;
  SIGNAL Logical_Operator_out1474_out1            : std_logic;
  SIGNAL Logical_Operator_out1475_out1            : std_logic;
  SIGNAL Logical_Operator_out1476_out1            : std_logic;
  SIGNAL Logical_Operator_out1477_out1            : std_logic;
  SIGNAL Logical_Operator_out1478_out1            : std_logic;
  SIGNAL Logical_Operator_out1479_out1            : std_logic;
  SIGNAL Logical_Operator_out1480_out1            : std_logic;
  SIGNAL Logical_Operator_out1481_out1            : std_logic;
  SIGNAL Logical_Operator_out1482_out1            : std_logic;
  SIGNAL Logical_Operator_out1483_out1            : std_logic;
  SIGNAL Logical_Operator_out1484_out1            : std_logic;
  SIGNAL Logical_Operator_out1485_out1            : std_logic;
  SIGNAL Logical_Operator_out1486_out1            : std_logic;
  SIGNAL Logical_Operator_out1487_out1            : std_logic;
  SIGNAL Logical_Operator_out1488_out1            : std_logic;
  SIGNAL Logical_Operator_out1489_out1            : std_logic;
  SIGNAL Logical_Operator_out1490_out1            : std_logic;
  SIGNAL Logical_Operator_out1491_out1            : std_logic;
  SIGNAL Logical_Operator_out1492_out1            : std_logic;
  SIGNAL Logical_Operator_out1493_out1            : std_logic;
  SIGNAL Logical_Operator_out1494_out1            : std_logic;
  SIGNAL Logical_Operator_out1495_out1            : std_logic;
  SIGNAL Logical_Operator_out1496_out1            : std_logic;
  SIGNAL Logical_Operator_out1497_out1            : std_logic;
  SIGNAL Logical_Operator_out1498_out1            : std_logic;
  SIGNAL Logical_Operator_out1499_out1            : std_logic;
  SIGNAL Logical_Operator_out1500_out1            : std_logic;
  SIGNAL Logical_Operator_out1501_out1            : std_logic;
  SIGNAL Logical_Operator_out1502_out1            : std_logic;
  SIGNAL Logical_Operator_out1503_out1            : std_logic;
  SIGNAL Logical_Operator_out1504_out1            : std_logic;
  SIGNAL Logical_Operator_out1505_out1            : std_logic;
  SIGNAL Logical_Operator_out1506_out1            : std_logic;
  SIGNAL Logical_Operator_out1507_out1            : std_logic;
  SIGNAL Logical_Operator_out1508_out1            : std_logic;
  SIGNAL Logical_Operator_out1509_out1            : std_logic;
  SIGNAL Logical_Operator_out1510_out1            : std_logic;
  SIGNAL Logical_Operator_out1511_out1            : std_logic;
  SIGNAL Logical_Operator_out1512_out1            : std_logic;
  SIGNAL Logical_Operator_out1513_out1            : std_logic;
  SIGNAL Logical_Operator_out1514_out1            : std_logic;
  SIGNAL Logical_Operator_out1515_out1            : std_logic;
  SIGNAL Logical_Operator_out1516_out1            : std_logic;
  SIGNAL Logical_Operator_out1517_out1            : std_logic;
  SIGNAL Logical_Operator_out1518_out1            : std_logic;
  SIGNAL Logical_Operator_out1519_out1            : std_logic;
  SIGNAL Logical_Operator_out1520_out1            : std_logic;
  SIGNAL Logical_Operator_out1521_out1            : std_logic;
  SIGNAL Logical_Operator_out1522_out1            : std_logic;
  SIGNAL Logical_Operator_out1523_out1            : std_logic;
  SIGNAL Logical_Operator_out1524_out1            : std_logic;
  SIGNAL Logical_Operator_out1525_out1            : std_logic;
  SIGNAL Logical_Operator_out1526_out1            : std_logic;
  SIGNAL Logical_Operator_out1527_out1            : std_logic;
  SIGNAL Logical_Operator_out1528_out1            : std_logic;
  SIGNAL Logical_Operator_out1529_out1            : std_logic;
  SIGNAL Logical_Operator_out1530_out1            : std_logic;
  SIGNAL Logical_Operator_out1531_out1            : std_logic;
  SIGNAL Logical_Operator_out1532_out1            : std_logic;
  SIGNAL Logical_Operator_out1533_out1            : std_logic;
  SIGNAL Logical_Operator_out1534_out1            : std_logic;
  SIGNAL Logical_Operator_out1535_out1            : std_logic;
  SIGNAL Logical_Operator_out1536_out1            : std_logic;
  SIGNAL Logical_Operator_out1537_out1            : std_logic;
  SIGNAL Logical_Operator_out1538_out1            : std_logic;
  SIGNAL Logical_Operator_out1539_out1            : std_logic;
  SIGNAL Logical_Operator_out1540_out1            : std_logic;
  SIGNAL Logical_Operator_out1541_out1            : std_logic;
  SIGNAL Logical_Operator_out1542_out1            : std_logic;
  SIGNAL Logical_Operator_out1543_out1            : std_logic;
  SIGNAL Logical_Operator_out1544_out1            : std_logic;
  SIGNAL Logical_Operator_out1545_out1            : std_logic;
  SIGNAL Logical_Operator_out1546_out1            : std_logic;
  SIGNAL Logical_Operator_out1547_out1            : std_logic;
  SIGNAL Logical_Operator_out1548_out1            : std_logic;
  SIGNAL Logical_Operator_out1549_out1            : std_logic;
  SIGNAL Logical_Operator_out1550_out1            : std_logic;
  SIGNAL Logical_Operator_out1551_out1            : std_logic;
  SIGNAL Logical_Operator_out1552_out1            : std_logic;
  SIGNAL Logical_Operator_out1553_out1            : std_logic;
  SIGNAL Logical_Operator_out1554_out1            : std_logic;
  SIGNAL Logical_Operator_out1555_out1            : std_logic;
  SIGNAL Logical_Operator_out1556_out1            : std_logic;
  SIGNAL Logical_Operator_out1557_out1            : std_logic;
  SIGNAL Logical_Operator_out1558_out1            : std_logic;
  SIGNAL Logical_Operator_out1559_out1            : std_logic;
  SIGNAL Logical_Operator_out1560_out1            : std_logic;
  SIGNAL Logical_Operator_out1561_out1            : std_logic;
  SIGNAL Logical_Operator_out1562_out1            : std_logic;
  SIGNAL Logical_Operator_out1563_out1            : std_logic;
  SIGNAL Logical_Operator_out1564_out1            : std_logic;
  SIGNAL Logical_Operator_out1565_out1            : std_logic;
  SIGNAL Logical_Operator_out1566_out1            : std_logic;
  SIGNAL Logical_Operator_out1567_out1            : std_logic;
  SIGNAL Logical_Operator_out1568_out1            : std_logic;
  SIGNAL Logical_Operator_out1569_out1            : std_logic;
  SIGNAL Logical_Operator_out1570_out1            : std_logic;
  SIGNAL Logical_Operator_out1571_out1            : std_logic;
  SIGNAL Logical_Operator_out1572_out1            : std_logic;
  SIGNAL Logical_Operator_out1573_out1            : std_logic;
  SIGNAL Logical_Operator_out1574_out1            : std_logic;
  SIGNAL Logical_Operator_out1575_out1            : std_logic;
  SIGNAL Logical_Operator_out1576_out1            : std_logic;
  SIGNAL Logical_Operator_out1577_out1            : std_logic;
  SIGNAL Logical_Operator_out1578_out1            : std_logic;
  SIGNAL Logical_Operator_out1579_out1            : std_logic;
  SIGNAL Logical_Operator_out1580_out1            : std_logic;
  SIGNAL Logical_Operator_out1581_out1            : std_logic;
  SIGNAL Logical_Operator_out1582_out1            : std_logic;
  SIGNAL Logical_Operator_out1583_out1            : std_logic;
  SIGNAL Logical_Operator_out1584_out1            : std_logic;
  SIGNAL Logical_Operator_out1585_out1            : std_logic;
  SIGNAL Logical_Operator_out1586_out1            : std_logic;
  SIGNAL Logical_Operator_out1587_out1            : std_logic;
  SIGNAL Logical_Operator_out1588_out1            : std_logic;
  SIGNAL Logical_Operator_out1589_out1            : std_logic;
  SIGNAL Logical_Operator_out1590_out1            : std_logic;
  SIGNAL Logical_Operator_out1591_out1            : std_logic;
  SIGNAL Logical_Operator_out1592_out1            : std_logic;
  SIGNAL Logical_Operator_out1593_out1            : std_logic;
  SIGNAL Logical_Operator_out1594_out1            : std_logic;
  SIGNAL Logical_Operator_out1595_out1            : std_logic;
  SIGNAL Logical_Operator_out1596_out1            : std_logic;
  SIGNAL Logical_Operator_out1597_out1            : std_logic;
  SIGNAL Logical_Operator_out1598_out1            : std_logic;
  SIGNAL Logical_Operator_out1599_out1            : std_logic;
  SIGNAL Logical_Operator_out1600_out1            : std_logic;
  SIGNAL Logical_Operator_out1601_out1            : std_logic;
  SIGNAL Logical_Operator_out1602_out1            : std_logic;
  SIGNAL Logical_Operator_out1603_out1            : std_logic;
  SIGNAL Logical_Operator_out1604_out1            : std_logic;
  SIGNAL Logical_Operator_out1605_out1            : std_logic;
  SIGNAL Logical_Operator_out1606_out1            : std_logic;
  SIGNAL Logical_Operator_out1607_out1            : std_logic;
  SIGNAL Logical_Operator_out1608_out1            : std_logic;
  SIGNAL Logical_Operator_out1609_out1            : std_logic;
  SIGNAL Logical_Operator_out1610_out1            : std_logic;
  SIGNAL Logical_Operator_out1611_out1            : std_logic;
  SIGNAL Logical_Operator_out1612_out1            : std_logic;
  SIGNAL Logical_Operator_out1613_out1            : std_logic;
  SIGNAL Logical_Operator_out1614_out1            : std_logic;
  SIGNAL Logical_Operator_out1615_out1            : std_logic;
  SIGNAL Logical_Operator_out1616_out1            : std_logic;
  SIGNAL Logical_Operator_out1617_out1            : std_logic;
  SIGNAL Logical_Operator_out1618_out1            : std_logic;
  SIGNAL Logical_Operator_out1619_out1            : std_logic;
  SIGNAL Logical_Operator_out1620_out1            : std_logic;
  SIGNAL Logical_Operator_out1621_out1            : std_logic;
  SIGNAL Logical_Operator_out1622_out1            : std_logic;
  SIGNAL Logical_Operator_out1623_out1            : std_logic;
  SIGNAL Logical_Operator_out1624_out1            : std_logic;
  SIGNAL Logical_Operator_out1625_out1            : std_logic;
  SIGNAL Logical_Operator_out1626_out1            : std_logic;
  SIGNAL Logical_Operator_out1627_out1            : std_logic;
  SIGNAL Logical_Operator_out1628_out1            : std_logic;
  SIGNAL Logical_Operator_out1629_out1            : std_logic;
  SIGNAL Logical_Operator_out1630_out1            : std_logic;
  SIGNAL Logical_Operator_out1631_out1            : std_logic;
  SIGNAL Logical_Operator_out1632_out1            : std_logic;
  SIGNAL Logical_Operator_out1633_out1            : std_logic;
  SIGNAL Logical_Operator_out1634_out1            : std_logic;
  SIGNAL Logical_Operator_out1635_out1            : std_logic;
  SIGNAL Logical_Operator_out1636_out1            : std_logic;
  SIGNAL Logical_Operator_out1637_out1            : std_logic;
  SIGNAL Logical_Operator_out1638_out1            : std_logic;
  SIGNAL Logical_Operator_out1639_out1            : std_logic;
  SIGNAL Logical_Operator_out1640_out1            : std_logic;
  SIGNAL Logical_Operator_out1641_out1            : std_logic;
  SIGNAL Logical_Operator_out1642_out1            : std_logic;
  SIGNAL Logical_Operator_out1643_out1            : std_logic;
  SIGNAL Logical_Operator_out1644_out1            : std_logic;
  SIGNAL Logical_Operator_out1645_out1            : std_logic;
  SIGNAL Logical_Operator_out1646_out1            : std_logic;
  SIGNAL Logical_Operator_out1647_out1            : std_logic;
  SIGNAL Logical_Operator_out1648_out1            : std_logic;
  SIGNAL Logical_Operator_out1649_out1            : std_logic;
  SIGNAL Logical_Operator_out1650_out1            : std_logic;
  SIGNAL Logical_Operator_out1651_out1            : std_logic;
  SIGNAL Logical_Operator_out1652_out1            : std_logic;
  SIGNAL Logical_Operator_out1653_out1            : std_logic;
  SIGNAL Logical_Operator_out1654_out1            : std_logic;
  SIGNAL Logical_Operator_out1655_out1            : std_logic;
  SIGNAL Logical_Operator_out1656_out1            : std_logic;
  SIGNAL Logical_Operator_out1657_out1            : std_logic;
  SIGNAL Logical_Operator_out1658_out1            : std_logic;
  SIGNAL Logical_Operator_out1659_out1            : std_logic;
  SIGNAL Logical_Operator_out1660_out1            : std_logic;
  SIGNAL Logical_Operator_out1661_out1            : std_logic;
  SIGNAL Logical_Operator_out1662_out1            : std_logic;
  SIGNAL Logical_Operator_out1663_out1            : std_logic;
  SIGNAL Logical_Operator_out1664_out1            : std_logic;
  SIGNAL Logical_Operator_out1665_out1            : std_logic;
  SIGNAL Logical_Operator_out1666_out1            : std_logic;
  SIGNAL Logical_Operator_out1667_out1            : std_logic;
  SIGNAL Logical_Operator_out1668_out1            : std_logic;
  SIGNAL Logical_Operator_out1669_out1            : std_logic;
  SIGNAL Logical_Operator_out1670_out1            : std_logic;
  SIGNAL Logical_Operator_out1671_out1            : std_logic;
  SIGNAL Logical_Operator_out1672_out1            : std_logic;
  SIGNAL Logical_Operator_out1673_out1            : std_logic;
  SIGNAL Logical_Operator_out1674_out1            : std_logic;
  SIGNAL Logical_Operator_out1675_out1            : std_logic;
  SIGNAL Logical_Operator_out1676_out1            : std_logic;
  SIGNAL Logical_Operator_out1677_out1            : std_logic;
  SIGNAL Logical_Operator_out1678_out1            : std_logic;
  SIGNAL Logical_Operator_out1679_out1            : std_logic;
  SIGNAL Logical_Operator_out1680_out1            : std_logic;
  SIGNAL Logical_Operator_out1681_out1            : std_logic;
  SIGNAL Logical_Operator_out1682_out1            : std_logic;
  SIGNAL Logical_Operator_out1683_out1            : std_logic;
  SIGNAL Logical_Operator_out1684_out1            : std_logic;
  SIGNAL Logical_Operator_out1685_out1            : std_logic;
  SIGNAL Logical_Operator_out1686_out1            : std_logic;
  SIGNAL Logical_Operator_out1687_out1            : std_logic;
  SIGNAL Logical_Operator_out1688_out1            : std_logic;
  SIGNAL Logical_Operator_out1689_out1            : std_logic;
  SIGNAL Logical_Operator_out1690_out1            : std_logic;
  SIGNAL Logical_Operator_out1691_out1            : std_logic;
  SIGNAL Logical_Operator_out1692_out1            : std_logic;
  SIGNAL Logical_Operator_out1693_out1            : std_logic;
  SIGNAL Logical_Operator_out1694_out1            : std_logic;
  SIGNAL Logical_Operator_out1695_out1            : std_logic;
  SIGNAL Logical_Operator_out1696_out1            : std_logic;
  SIGNAL Logical_Operator_out1697_out1            : std_logic;
  SIGNAL Logical_Operator_out1698_out1            : std_logic;
  SIGNAL Logical_Operator_out1699_out1            : std_logic;
  SIGNAL Logical_Operator_out1700_out1            : std_logic;
  SIGNAL Logical_Operator_out1701_out1            : std_logic;
  SIGNAL Logical_Operator_out1702_out1            : std_logic;
  SIGNAL Logical_Operator_out1703_out1            : std_logic;
  SIGNAL Logical_Operator_out1704_out1            : std_logic;
  SIGNAL Logical_Operator_out1705_out1            : std_logic;
  SIGNAL Logical_Operator_out1706_out1            : std_logic;
  SIGNAL Logical_Operator_out1707_out1            : std_logic;
  SIGNAL Logical_Operator_out1708_out1            : std_logic;
  SIGNAL Logical_Operator_out1709_out1            : std_logic;
  SIGNAL Logical_Operator_out1710_out1            : std_logic;
  SIGNAL Logical_Operator_out1711_out1            : std_logic;
  SIGNAL Logical_Operator_out1712_out1            : std_logic;
  SIGNAL Logical_Operator_out1713_out1            : std_logic;
  SIGNAL Logical_Operator_out1714_out1            : std_logic;
  SIGNAL Logical_Operator_out1715_out1            : std_logic;
  SIGNAL Logical_Operator_out1716_out1            : std_logic;
  SIGNAL Logical_Operator_out1717_out1            : std_logic;
  SIGNAL Logical_Operator_out1718_out1            : std_logic;
  SIGNAL Logical_Operator_out1719_out1            : std_logic;
  SIGNAL Logical_Operator_out1720_out1            : std_logic;
  SIGNAL Logical_Operator_out1721_out1            : std_logic;
  SIGNAL Logical_Operator_out1722_out1            : std_logic;
  SIGNAL Logical_Operator_out1723_out1            : std_logic;
  SIGNAL Logical_Operator_out1724_out1            : std_logic;
  SIGNAL Logical_Operator_out1725_out1            : std_logic;
  SIGNAL Logical_Operator_out1726_out1            : std_logic;
  SIGNAL Logical_Operator_out1727_out1            : std_logic;
  SIGNAL Logical_Operator_out1728_out1            : std_logic;
  SIGNAL Logical_Operator_out1729_out1            : std_logic;
  SIGNAL Logical_Operator_out1730_out1            : std_logic;
  SIGNAL Logical_Operator_out1731_out1            : std_logic;
  SIGNAL Logical_Operator_out1732_out1            : std_logic;
  SIGNAL Logical_Operator_out1733_out1            : std_logic;
  SIGNAL Logical_Operator_out1734_out1            : std_logic;
  SIGNAL Logical_Operator_out1735_out1            : std_logic;
  SIGNAL Logical_Operator_out1736_out1            : std_logic;
  SIGNAL Logical_Operator_out1737_out1            : std_logic;
  SIGNAL Logical_Operator_out1738_out1            : std_logic;
  SIGNAL Logical_Operator_out1739_out1            : std_logic;
  SIGNAL Logical_Operator_out1740_out1            : std_logic;
  SIGNAL Logical_Operator_out1741_out1            : std_logic;
  SIGNAL Logical_Operator_out1742_out1            : std_logic;
  SIGNAL Logical_Operator_out1743_out1            : std_logic;
  SIGNAL Logical_Operator_out1744_out1            : std_logic;
  SIGNAL Logical_Operator_out1745_out1            : std_logic;
  SIGNAL Logical_Operator_out1746_out1            : std_logic;
  SIGNAL Logical_Operator_out1747_out1            : std_logic;
  SIGNAL Logical_Operator_out1748_out1            : std_logic;
  SIGNAL Logical_Operator_out1749_out1            : std_logic;
  SIGNAL Logical_Operator_out1750_out1            : std_logic;
  SIGNAL Logical_Operator_out1751_out1            : std_logic;
  SIGNAL Logical_Operator_out1752_out1            : std_logic;
  SIGNAL Logical_Operator_out1753_out1            : std_logic;
  SIGNAL Logical_Operator_out1754_out1            : std_logic;
  SIGNAL Logical_Operator_out1755_out1            : std_logic;
  SIGNAL Logical_Operator_out1756_out1            : std_logic;
  SIGNAL Logical_Operator_out1757_out1            : std_logic;
  SIGNAL Logical_Operator_out1758_out1            : std_logic;
  SIGNAL Logical_Operator_out1759_out1            : std_logic;
  SIGNAL Logical_Operator_out1760_out1            : std_logic;
  SIGNAL Logical_Operator_out1761_out1            : std_logic;
  SIGNAL Logical_Operator_out1762_out1            : std_logic;
  SIGNAL Logical_Operator_out1763_out1            : std_logic;
  SIGNAL Logical_Operator_out1764_out1            : std_logic;
  SIGNAL Logical_Operator_out1765_out1            : std_logic;
  SIGNAL Logical_Operator_out1766_out1            : std_logic;
  SIGNAL Logical_Operator_out1767_out1            : std_logic;
  SIGNAL Logical_Operator_out1768_out1            : std_logic;
  SIGNAL Logical_Operator_out1769_out1            : std_logic;
  SIGNAL Logical_Operator_out1770_out1            : std_logic;
  SIGNAL Logical_Operator_out1771_out1            : std_logic;
  SIGNAL Logical_Operator_out1772_out1            : std_logic;
  SIGNAL Logical_Operator_out1773_out1            : std_logic;
  SIGNAL Logical_Operator_out1774_out1            : std_logic;
  SIGNAL Logical_Operator_out1775_out1            : std_logic;
  SIGNAL Logical_Operator_out1776_out1            : std_logic;
  SIGNAL Logical_Operator_out1777_out1            : std_logic;
  SIGNAL Logical_Operator_out1778_out1            : std_logic;
  SIGNAL Logical_Operator_out1779_out1            : std_logic;
  SIGNAL Logical_Operator_out1780_out1            : std_logic;
  SIGNAL Logical_Operator_out1781_out1            : std_logic;
  SIGNAL Logical_Operator_out1782_out1            : std_logic;
  SIGNAL Logical_Operator_out1783_out1            : std_logic;
  SIGNAL Logical_Operator_out1784_out1            : std_logic;
  SIGNAL Logical_Operator_out1785_out1            : std_logic;
  SIGNAL Logical_Operator_out1786_out1            : std_logic;
  SIGNAL Logical_Operator_out1787_out1            : std_logic;
  SIGNAL Logical_Operator_out1788_out1            : std_logic;
  SIGNAL Logical_Operator_out1789_out1            : std_logic;
  SIGNAL Logical_Operator_out1790_out1            : std_logic;
  SIGNAL Logical_Operator_out1791_out1            : std_logic;
  SIGNAL Logical_Operator_out1792_out1            : std_logic;
  SIGNAL Logical_Operator_out1793_out1            : std_logic;
  SIGNAL Logical_Operator_out1794_out1            : std_logic;
  SIGNAL Logical_Operator_out1795_out1            : std_logic;
  SIGNAL Logical_Operator_out1796_out1            : std_logic;
  SIGNAL Logical_Operator_out1797_out1            : std_logic;
  SIGNAL Logical_Operator_out1798_out1            : std_logic;
  SIGNAL Logical_Operator_out1799_out1            : std_logic;
  SIGNAL Logical_Operator_out1800_out1            : std_logic;
  SIGNAL Logical_Operator_out1801_out1            : std_logic;
  SIGNAL Logical_Operator_out1802_out1            : std_logic;
  SIGNAL Logical_Operator_out1803_out1            : std_logic;
  SIGNAL Logical_Operator_out1804_out1            : std_logic;
  SIGNAL Logical_Operator_out1805_out1            : std_logic;
  SIGNAL Logical_Operator_out1806_out1            : std_logic;
  SIGNAL Logical_Operator_out1807_out1            : std_logic;
  SIGNAL Logical_Operator_out1808_out1            : std_logic;
  SIGNAL Logical_Operator_out1809_out1            : std_logic;
  SIGNAL Logical_Operator_out1810_out1            : std_logic;
  SIGNAL Logical_Operator_out1811_out1            : std_logic;
  SIGNAL Logical_Operator_out1812_out1            : std_logic;
  SIGNAL Logical_Operator_out1813_out1            : std_logic;
  SIGNAL Logical_Operator_out1814_out1            : std_logic;
  SIGNAL Logical_Operator_out1815_out1            : std_logic;
  SIGNAL Logical_Operator_out1816_out1            : std_logic;
  SIGNAL Logical_Operator_out1817_out1            : std_logic;
  SIGNAL Logical_Operator_out1818_out1            : std_logic;
  SIGNAL Logical_Operator_out1819_out1            : std_logic;
  SIGNAL Logical_Operator_out1820_out1            : std_logic;
  SIGNAL Logical_Operator_out1821_out1            : std_logic;
  SIGNAL Logical_Operator_out1822_out1            : std_logic;
  SIGNAL Logical_Operator_out1823_out1            : std_logic;
  SIGNAL Logical_Operator_out1824_out1            : std_logic;
  SIGNAL Logical_Operator_out1825_out1            : std_logic;
  SIGNAL Logical_Operator_out1826_out1            : std_logic;
  SIGNAL Logical_Operator_out1827_out1            : std_logic;
  SIGNAL Logical_Operator_out1828_out1            : std_logic;
  SIGNAL Logical_Operator_out1829_out1            : std_logic;
  SIGNAL Logical_Operator_out1830_out1            : std_logic;
  SIGNAL Logical_Operator_out1831_out1            : std_logic;
  SIGNAL Logical_Operator_out1832_out1            : std_logic;
  SIGNAL Logical_Operator_out1833_out1            : std_logic;
  SIGNAL Logical_Operator_out1834_out1            : std_logic;
  SIGNAL Logical_Operator_out1835_out1            : std_logic;
  SIGNAL Logical_Operator_out1836_out1            : std_logic;
  SIGNAL Logical_Operator_out1837_out1            : std_logic;
  SIGNAL Logical_Operator_out1838_out1            : std_logic;
  SIGNAL Logical_Operator_out1839_out1            : std_logic;
  SIGNAL Logical_Operator_out1840_out1            : std_logic;
  SIGNAL Logical_Operator_out1841_out1            : std_logic;
  SIGNAL Logical_Operator_out1842_out1            : std_logic;
  SIGNAL Logical_Operator_out1843_out1            : std_logic;
  SIGNAL Logical_Operator_out1844_out1            : std_logic;
  SIGNAL Logical_Operator_out1845_out1            : std_logic;
  SIGNAL Logical_Operator_out1846_out1            : std_logic;
  SIGNAL Logical_Operator_out1847_out1            : std_logic;
  SIGNAL Logical_Operator_out1848_out1            : std_logic;
  SIGNAL Logical_Operator_out1849_out1            : std_logic;
  SIGNAL Logical_Operator_out1850_out1            : std_logic;
  SIGNAL Logical_Operator_out1851_out1            : std_logic;
  SIGNAL Logical_Operator_out1852_out1            : std_logic;
  SIGNAL Logical_Operator_out1853_out1            : std_logic;
  SIGNAL Logical_Operator_out1854_out1            : std_logic;
  SIGNAL Logical_Operator_out1855_out1            : std_logic;
  SIGNAL Logical_Operator_out1856_out1            : std_logic;
  SIGNAL Logical_Operator_out1857_out1            : std_logic;
  SIGNAL Logical_Operator_out1858_out1            : std_logic;
  SIGNAL Logical_Operator_out1859_out1            : std_logic;
  SIGNAL Logical_Operator_out1860_out1            : std_logic;
  SIGNAL Logical_Operator_out1861_out1            : std_logic;
  SIGNAL Logical_Operator_out1862_out1            : std_logic;
  SIGNAL Logical_Operator_out1863_out1            : std_logic;
  SIGNAL Logical_Operator_out1864_out1            : std_logic;
  SIGNAL Logical_Operator_out1865_out1            : std_logic;
  SIGNAL Logical_Operator_out1866_out1            : std_logic;
  SIGNAL Logical_Operator_out1867_out1            : std_logic;
  SIGNAL Logical_Operator_out1868_out1            : std_logic;
  SIGNAL Logical_Operator_out1869_out1            : std_logic;
  SIGNAL Logical_Operator_out1870_out1            : std_logic;
  SIGNAL Logical_Operator_out1871_out1            : std_logic;
  SIGNAL Logical_Operator_out1872_out1            : std_logic;
  SIGNAL Logical_Operator_out1873_out1            : std_logic;
  SIGNAL Logical_Operator_out1874_out1            : std_logic;
  SIGNAL Logical_Operator_out1875_out1            : std_logic;
  SIGNAL Logical_Operator_out1876_out1            : std_logic;
  SIGNAL Logical_Operator_out1877_out1            : std_logic;
  SIGNAL Logical_Operator_out1878_out1            : std_logic;
  SIGNAL Logical_Operator_out1879_out1            : std_logic;
  SIGNAL Logical_Operator_out1880_out1            : std_logic;
  SIGNAL Logical_Operator_out1881_out1            : std_logic;
  SIGNAL Logical_Operator_out1882_out1            : std_logic;
  SIGNAL Logical_Operator_out1883_out1            : std_logic;
  SIGNAL Logical_Operator_out1884_out1            : std_logic;
  SIGNAL Logical_Operator_out1885_out1            : std_logic;
  SIGNAL Logical_Operator_out1886_out1            : std_logic;
  SIGNAL Logical_Operator_out1887_out1            : std_logic;
  SIGNAL Logical_Operator_out1888_out1            : std_logic;
  SIGNAL Logical_Operator_out1889_out1            : std_logic;
  SIGNAL Logical_Operator_out1890_out1            : std_logic;
  SIGNAL Logical_Operator_out1891_out1            : std_logic;
  SIGNAL Logical_Operator_out1892_out1            : std_logic;
  SIGNAL Logical_Operator_out1893_out1            : std_logic;
  SIGNAL Logical_Operator_out1894_out1            : std_logic;
  SIGNAL Logical_Operator_out1895_out1            : std_logic;
  SIGNAL Logical_Operator_out1896_out1            : std_logic;
  SIGNAL Logical_Operator_out1897_out1            : std_logic;
  SIGNAL Logical_Operator_out1898_out1            : std_logic;
  SIGNAL Logical_Operator_out1899_out1            : std_logic;
  SIGNAL Logical_Operator_out1900_out1            : std_logic;
  SIGNAL Logical_Operator_out1901_out1            : std_logic;
  SIGNAL Logical_Operator_out1902_out1            : std_logic;
  SIGNAL Logical_Operator_out1903_out1            : std_logic;
  SIGNAL Logical_Operator_out1904_out1            : std_logic;
  SIGNAL Logical_Operator_out1905_out1            : std_logic;
  SIGNAL Logical_Operator_out1906_out1            : std_logic;
  SIGNAL Logical_Operator_out1907_out1            : std_logic;
  SIGNAL Logical_Operator_out1908_out1            : std_logic;
  SIGNAL Logical_Operator_out1909_out1            : std_logic;
  SIGNAL Logical_Operator_out1910_out1            : std_logic;
  SIGNAL Logical_Operator_out1911_out1            : std_logic;
  SIGNAL Logical_Operator_out1912_out1            : std_logic;
  SIGNAL Logical_Operator_out1913_out1            : std_logic;
  SIGNAL Logical_Operator_out1914_out1            : std_logic;
  SIGNAL Logical_Operator_out1915_out1            : std_logic;
  SIGNAL Logical_Operator_out1916_out1            : std_logic;
  SIGNAL Logical_Operator_out1917_out1            : std_logic;
  SIGNAL Logical_Operator_out1918_out1            : std_logic;
  SIGNAL Logical_Operator_out1919_out1            : std_logic;
  SIGNAL Logical_Operator_out1920_out1            : std_logic;
  SIGNAL Logical_Operator_out1921_out1            : std_logic;
  SIGNAL Logical_Operator_out1922_out1            : std_logic;
  SIGNAL Logical_Operator_out1923_out1            : std_logic;
  SIGNAL Logical_Operator_out1924_out1            : std_logic;
  SIGNAL Logical_Operator_out1925_out1            : std_logic;
  SIGNAL Logical_Operator_out1926_out1            : std_logic;
  SIGNAL Logical_Operator_out1927_out1            : std_logic;
  SIGNAL Logical_Operator_out1928_out1            : std_logic;
  SIGNAL Logical_Operator_out1929_out1            : std_logic;
  SIGNAL Logical_Operator_out1930_out1            : std_logic;
  SIGNAL Logical_Operator_out1931_out1            : std_logic;
  SIGNAL Logical_Operator_out1932_out1            : std_logic;
  SIGNAL Logical_Operator_out1933_out1            : std_logic;
  SIGNAL Logical_Operator_out1934_out1            : std_logic;
  SIGNAL Logical_Operator_out1935_out1            : std_logic;
  SIGNAL Logical_Operator_out1936_out1            : std_logic;
  SIGNAL Logical_Operator_out1937_out1            : std_logic;
  SIGNAL Logical_Operator_out1938_out1            : std_logic;
  SIGNAL Logical_Operator_out1939_out1            : std_logic;
  SIGNAL Logical_Operator_out1940_out1            : std_logic;
  SIGNAL Logical_Operator_out1941_out1            : std_logic;
  SIGNAL Logical_Operator_out1942_out1            : std_logic;
  SIGNAL Logical_Operator_out1943_out1            : std_logic;
  SIGNAL Logical_Operator_out1944_out1            : std_logic;
  SIGNAL Logical_Operator_out1945_out1            : std_logic;
  SIGNAL Logical_Operator_out1946_out1            : std_logic;
  SIGNAL Logical_Operator_out1947_out1            : std_logic;
  SIGNAL Logical_Operator_out1948_out1            : std_logic;
  SIGNAL Logical_Operator_out1949_out1            : std_logic;
  SIGNAL Logical_Operator_out1950_out1            : std_logic;
  SIGNAL Logical_Operator_out1951_out1            : std_logic;
  SIGNAL Logical_Operator_out1952_out1            : std_logic;
  SIGNAL Logical_Operator_out1953_out1            : std_logic;
  SIGNAL Logical_Operator_out1954_out1            : std_logic;
  SIGNAL Logical_Operator_out1955_out1            : std_logic;
  SIGNAL Logical_Operator_out1956_out1            : std_logic;
  SIGNAL Logical_Operator_out1957_out1            : std_logic;
  SIGNAL Logical_Operator_out1958_out1            : std_logic;
  SIGNAL Logical_Operator_out1959_out1            : std_logic;
  SIGNAL Logical_Operator_out1960_out1            : std_logic;
  SIGNAL Logical_Operator_out1961_out1            : std_logic;
  SIGNAL Logical_Operator_out1962_out1            : std_logic;
  SIGNAL Logical_Operator_out1963_out1            : std_logic;
  SIGNAL Logical_Operator_out1964_out1            : std_logic;
  SIGNAL Logical_Operator_out1965_out1            : std_logic;
  SIGNAL Logical_Operator_out1966_out1            : std_logic;
  SIGNAL Logical_Operator_out1967_out1            : std_logic;
  SIGNAL Logical_Operator_out1968_out1            : std_logic;
  SIGNAL Logical_Operator_out1969_out1            : std_logic;
  SIGNAL Logical_Operator_out1970_out1            : std_logic;
  SIGNAL Logical_Operator_out1971_out1            : std_logic;
  SIGNAL Logical_Operator_out1972_out1            : std_logic;
  SIGNAL Logical_Operator_out1973_out1            : std_logic;
  SIGNAL Logical_Operator_out1974_out1            : std_logic;
  SIGNAL Logical_Operator_out1975_out1            : std_logic;
  SIGNAL Logical_Operator_out1976_out1            : std_logic;
  SIGNAL Logical_Operator_out1977_out1            : std_logic;
  SIGNAL Logical_Operator_out1978_out1            : std_logic;
  SIGNAL Logical_Operator_out1979_out1            : std_logic;
  SIGNAL Logical_Operator_out1980_out1            : std_logic;
  SIGNAL Logical_Operator_out1981_out1            : std_logic;
  SIGNAL Logical_Operator_out1982_out1            : std_logic;
  SIGNAL Logical_Operator_out1983_out1            : std_logic;
  SIGNAL Logical_Operator_out1984_out1            : std_logic;
  SIGNAL Logical_Operator_out1985_out1            : std_logic;
  SIGNAL Logical_Operator_out1986_out1            : std_logic;
  SIGNAL Logical_Operator_out1987_out1            : std_logic;
  SIGNAL Logical_Operator_out1988_out1            : std_logic;
  SIGNAL Logical_Operator_out1989_out1            : std_logic;
  SIGNAL Logical_Operator_out1990_out1            : std_logic;
  SIGNAL Logical_Operator_out1991_out1            : std_logic;
  SIGNAL Logical_Operator_out1992_out1            : std_logic;
  SIGNAL Logical_Operator_out1993_out1            : std_logic;
  SIGNAL Logical_Operator_out1994_out1            : std_logic;
  SIGNAL Logical_Operator_out1995_out1            : std_logic;
  SIGNAL Logical_Operator_out1996_out1            : std_logic;
  SIGNAL Logical_Operator_out1997_out1            : std_logic;
  SIGNAL Logical_Operator_out1998_out1            : std_logic;
  SIGNAL Logical_Operator_out1999_out1            : std_logic;
  SIGNAL Logical_Operator_out2000_out1            : std_logic;
  SIGNAL Logical_Operator_out2001_out1            : std_logic;
  SIGNAL Logical_Operator_out2002_out1            : std_logic;
  SIGNAL Logical_Operator_out2003_out1            : std_logic;
  SIGNAL Logical_Operator_out2004_out1            : std_logic;
  SIGNAL Logical_Operator_out2005_out1            : std_logic;
  SIGNAL Logical_Operator_out2006_out1            : std_logic;
  SIGNAL Logical_Operator_out2007_out1            : std_logic;
  SIGNAL Logical_Operator_out2008_out1            : std_logic;
  SIGNAL Logical_Operator_out2009_out1            : std_logic;
  SIGNAL Logical_Operator_out2010_out1            : std_logic;
  SIGNAL Logical_Operator_out2011_out1            : std_logic;
  SIGNAL Logical_Operator_out2012_out1            : std_logic;
  SIGNAL Logical_Operator_out2013_out1            : std_logic;
  SIGNAL Logical_Operator_out2014_out1            : std_logic;
  SIGNAL Logical_Operator_out2015_out1            : std_logic;
  SIGNAL Logical_Operator_out2016_out1            : std_logic;
  SIGNAL Logical_Operator_out2017_out1            : std_logic;
  SIGNAL Logical_Operator_out2018_out1            : std_logic;
  SIGNAL Logical_Operator_out2019_out1            : std_logic;
  SIGNAL Logical_Operator_out2020_out1            : std_logic;
  SIGNAL Logical_Operator_out2021_out1            : std_logic;
  SIGNAL Logical_Operator_out2022_out1            : std_logic;
  SIGNAL Logical_Operator_out2023_out1            : std_logic;
  SIGNAL Logical_Operator_out2024_out1            : std_logic;
  SIGNAL Logical_Operator_out2025_out1            : std_logic;
  SIGNAL Logical_Operator_out2026_out1            : std_logic;
  SIGNAL Logical_Operator_out2027_out1            : std_logic;
  SIGNAL Logical_Operator_out2028_out1            : std_logic;
  SIGNAL Logical_Operator_out2029_out1            : std_logic;
  SIGNAL Logical_Operator_out2030_out1            : std_logic;
  SIGNAL Logical_Operator_out2031_out1            : std_logic;
  SIGNAL Logical_Operator_out2032_out1            : std_logic;
  SIGNAL Logical_Operator_out2033_out1            : std_logic;
  SIGNAL Logical_Operator_out2034_out1            : std_logic;
  SIGNAL Logical_Operator_out2035_out1            : std_logic;
  SIGNAL Logical_Operator_out2036_out1            : std_logic;
  SIGNAL Logical_Operator_out2037_out1            : std_logic;
  SIGNAL Logical_Operator_out2038_out1            : std_logic;
  SIGNAL Logical_Operator_out2039_out1            : std_logic;
  SIGNAL Logical_Operator_out2040_out1            : std_logic;
  SIGNAL Logical_Operator_out2041_out1            : std_logic;
  SIGNAL Logical_Operator_out2042_out1            : std_logic;
  SIGNAL Logical_Operator_out2043_out1            : std_logic;
  SIGNAL Logical_Operator_out2044_out1            : std_logic;
  SIGNAL Logical_Operator_out2045_out1            : std_logic;
  SIGNAL Logical_Operator_out2046_out1            : std_logic;
  SIGNAL Logical_Operator_out2047_out1            : std_logic;
  SIGNAL Logical_Operator_out2048_out1            : std_logic;
  SIGNAL Logical_Operator_out2049_out1            : std_logic;
  SIGNAL Logical_Operator_out2050_out1            : std_logic;
  SIGNAL Logical_Operator_out2051_out1            : std_logic;
  SIGNAL Logical_Operator_out2052_out1            : std_logic;
  SIGNAL Logical_Operator_out2053_out1            : std_logic;
  SIGNAL Logical_Operator_out2054_out1            : std_logic;
  SIGNAL Logical_Operator_out2055_out1            : std_logic;
  SIGNAL Logical_Operator_out2056_out1            : std_logic;
  SIGNAL Logical_Operator_out2057_out1            : std_logic;
  SIGNAL Logical_Operator_out2058_out1            : std_logic;
  SIGNAL Logical_Operator_out2059_out1            : std_logic;
  SIGNAL Logical_Operator_out2060_out1            : std_logic;
  SIGNAL Logical_Operator_out2061_out1            : std_logic;
  SIGNAL Logical_Operator_out2062_out1            : std_logic;
  SIGNAL Logical_Operator_out2063_out1            : std_logic;
  SIGNAL Logical_Operator_out2064_out1            : std_logic;
  SIGNAL Logical_Operator_out2065_out1            : std_logic;
  SIGNAL Logical_Operator_out2066_out1            : std_logic;
  SIGNAL Logical_Operator_out2067_out1            : std_logic;
  SIGNAL Logical_Operator_out2068_out1            : std_logic;
  SIGNAL Logical_Operator_out2069_out1            : std_logic;
  SIGNAL Logical_Operator_out2070_out1            : std_logic;
  SIGNAL Logical_Operator_out2071_out1            : std_logic;
  SIGNAL Logical_Operator_out2072_out1            : std_logic;
  SIGNAL Logical_Operator_out2073_out1            : std_logic;
  SIGNAL Logical_Operator_out2074_out1            : std_logic;
  SIGNAL Logical_Operator_out2075_out1            : std_logic;
  SIGNAL Logical_Operator_out2076_out1            : std_logic;
  SIGNAL Logical_Operator_out2077_out1            : std_logic;
  SIGNAL Logical_Operator_out2078_out1            : std_logic;
  SIGNAL Logical_Operator_out2079_out1            : std_logic;
  SIGNAL Logical_Operator_out2080_out1            : std_logic;
  SIGNAL Logical_Operator_out2081_out1            : std_logic;
  SIGNAL Logical_Operator_out2082_out1            : std_logic;
  SIGNAL Logical_Operator_out2083_out1            : std_logic;
  SIGNAL Logical_Operator_out2084_out1            : std_logic;
  SIGNAL Logical_Operator_out2085_out1            : std_logic;
  SIGNAL Logical_Operator_out2086_out1            : std_logic;
  SIGNAL Logical_Operator_out2087_out1            : std_logic;
  SIGNAL Logical_Operator_out2088_out1            : std_logic;
  SIGNAL Logical_Operator_out2089_out1            : std_logic;
  SIGNAL Logical_Operator_out2090_out1            : std_logic;
  SIGNAL Logical_Operator_out2091_out1            : std_logic;
  SIGNAL Logical_Operator_out2092_out1            : std_logic;
  SIGNAL Logical_Operator_out2093_out1            : std_logic;
  SIGNAL Logical_Operator_out2094_out1            : std_logic;
  SIGNAL Logical_Operator_out2095_out1            : std_logic;
  SIGNAL Logical_Operator_out2096_out1            : std_logic;
  SIGNAL Logical_Operator_out2097_out1            : std_logic;
  SIGNAL Logical_Operator_out2098_out1            : std_logic;
  SIGNAL Logical_Operator_out2099_out1            : std_logic;
  SIGNAL Logical_Operator_out2100_out1            : std_logic;
  SIGNAL Logical_Operator_out2101_out1            : std_logic;
  SIGNAL Logical_Operator_out2102_out1            : std_logic;
  SIGNAL Logical_Operator_out2103_out1            : std_logic;
  SIGNAL Logical_Operator_out2104_out1            : std_logic;
  SIGNAL Logical_Operator_out2105_out1            : std_logic;
  SIGNAL Logical_Operator_out2106_out1            : std_logic;
  SIGNAL Logical_Operator_out2107_out1            : std_logic;
  SIGNAL Logical_Operator_out2108_out1            : std_logic;
  SIGNAL Logical_Operator_out2109_out1            : std_logic;
  SIGNAL Logical_Operator_out2110_out1            : std_logic;
  SIGNAL Logical_Operator_out2111_out1            : std_logic;
  SIGNAL Logical_Operator_out2112_out1            : std_logic;
  SIGNAL Logical_Operator_out2113_out1            : std_logic;
  SIGNAL Logical_Operator_out2114_out1            : std_logic;
  SIGNAL Logical_Operator_out2115_out1            : std_logic;
  SIGNAL Logical_Operator_out2116_out1            : std_logic;
  SIGNAL Logical_Operator_out2117_out1            : std_logic;
  SIGNAL Logical_Operator_out2118_out1            : std_logic;
  SIGNAL Logical_Operator_out2119_out1            : std_logic;
  SIGNAL Logical_Operator_out2120_out1            : std_logic;
  SIGNAL Logical_Operator_out2121_out1            : std_logic;
  SIGNAL Logical_Operator_out2122_out1            : std_logic;
  SIGNAL Logical_Operator_out2123_out1            : std_logic;
  SIGNAL Logical_Operator_out2124_out1            : std_logic;
  SIGNAL Logical_Operator_out2125_out1            : std_logic;
  SIGNAL Logical_Operator_out2126_out1            : std_logic;
  SIGNAL Logical_Operator_out2127_out1            : std_logic;
  SIGNAL Logical_Operator_out2128_out1            : std_logic;
  SIGNAL Logical_Operator_out2129_out1            : std_logic;
  SIGNAL Logical_Operator_out2130_out1            : std_logic;
  SIGNAL Logical_Operator_out2131_out1            : std_logic;
  SIGNAL Logical_Operator_out2132_out1            : std_logic;
  SIGNAL Logical_Operator_out2133_out1            : std_logic;
  SIGNAL Logical_Operator_out2134_out1            : std_logic;
  SIGNAL Logical_Operator_out2135_out1            : std_logic;
  SIGNAL Logical_Operator_out2136_out1            : std_logic;
  SIGNAL Logical_Operator_out2137_out1            : std_logic;
  SIGNAL Logical_Operator_out2138_out1            : std_logic;
  SIGNAL Logical_Operator_out2139_out1            : std_logic;
  SIGNAL Logical_Operator_out2140_out1            : std_logic;
  SIGNAL Logical_Operator_out2141_out1            : std_logic;
  SIGNAL Logical_Operator_out2142_out1            : std_logic;
  SIGNAL Logical_Operator_out2143_out1            : std_logic;
  SIGNAL Logical_Operator_out2144_out1            : std_logic;
  SIGNAL Logical_Operator_out2145_out1            : std_logic;
  SIGNAL Logical_Operator_out2146_out1            : std_logic;
  SIGNAL Logical_Operator_out2147_out1            : std_logic;
  SIGNAL Logical_Operator_out2148_out1            : std_logic;
  SIGNAL Logical_Operator_out2149_out1            : std_logic;
  SIGNAL Logical_Operator_out2150_out1            : std_logic;
  SIGNAL Logical_Operator_out2151_out1            : std_logic;
  SIGNAL Logical_Operator_out2152_out1            : std_logic;
  SIGNAL Logical_Operator_out2153_out1            : std_logic;
  SIGNAL Logical_Operator_out2154_out1            : std_logic;
  SIGNAL Logical_Operator_out2155_out1            : std_logic;
  SIGNAL Logical_Operator_out2156_out1            : std_logic;
  SIGNAL Logical_Operator_out2157_out1            : std_logic;
  SIGNAL Logical_Operator_out2158_out1            : std_logic;
  SIGNAL Logical_Operator_out2159_out1            : std_logic;
  SIGNAL Logical_Operator_out2160_out1            : std_logic;
  SIGNAL Logical_Operator_out2161_out1            : std_logic;
  SIGNAL Logical_Operator_out2162_out1            : std_logic;
  SIGNAL Logical_Operator_out2163_out1            : std_logic;
  SIGNAL Logical_Operator_out2164_out1            : std_logic;
  SIGNAL Logical_Operator_out2165_out1            : std_logic;
  SIGNAL Logical_Operator_out2166_out1            : std_logic;
  SIGNAL Logical_Operator_out2167_out1            : std_logic;
  SIGNAL Logical_Operator_out2168_out1            : std_logic;
  SIGNAL Logical_Operator_out2169_out1            : std_logic;
  SIGNAL Logical_Operator_out2170_out1            : std_logic;
  SIGNAL Logical_Operator_out2171_out1            : std_logic;
  SIGNAL Logical_Operator_out2172_out1            : std_logic;
  SIGNAL Logical_Operator_out2173_out1            : std_logic;
  SIGNAL Logical_Operator_out2174_out1            : std_logic;
  SIGNAL Logical_Operator_out2175_out1            : std_logic;
  SIGNAL Logical_Operator_out2176_out1            : std_logic;
  SIGNAL Logical_Operator_out2177_out1            : std_logic;
  SIGNAL Logical_Operator_out2178_out1            : std_logic;
  SIGNAL Logical_Operator_out2179_out1            : std_logic;
  SIGNAL Logical_Operator_out2180_out1            : std_logic;
  SIGNAL Logical_Operator_out2181_out1            : std_logic;
  SIGNAL Logical_Operator_out2182_out1            : std_logic;
  SIGNAL Logical_Operator_out2183_out1            : std_logic;
  SIGNAL Logical_Operator_out2184_out1            : std_logic;
  SIGNAL Logical_Operator_out2185_out1            : std_logic;
  SIGNAL Logical_Operator_out2186_out1            : std_logic;
  SIGNAL Logical_Operator_out2187_out1            : std_logic;
  SIGNAL Logical_Operator_out2188_out1            : std_logic;
  SIGNAL Logical_Operator_out2189_out1            : std_logic;
  SIGNAL Logical_Operator_out2190_out1            : std_logic;
  SIGNAL Logical_Operator_out2191_out1            : std_logic;
  SIGNAL Logical_Operator_out2192_out1            : std_logic;
  SIGNAL Logical_Operator_out2193_out1            : std_logic;
  SIGNAL Logical_Operator_out2194_out1            : std_logic;
  SIGNAL Logical_Operator_out2195_out1            : std_logic;
  SIGNAL Logical_Operator_out2196_out1            : std_logic;
  SIGNAL Logical_Operator_out2197_out1            : std_logic;
  SIGNAL Logical_Operator_out2198_out1            : std_logic;
  SIGNAL Logical_Operator_out2199_out1            : std_logic;
  SIGNAL Logical_Operator_out2200_out1            : std_logic;
  SIGNAL Logical_Operator_out2201_out1            : std_logic;
  SIGNAL Logical_Operator_out2202_out1            : std_logic;
  SIGNAL Logical_Operator_out2203_out1            : std_logic;
  SIGNAL Logical_Operator_out2204_out1            : std_logic;
  SIGNAL Logical_Operator_out2205_out1            : std_logic;
  SIGNAL Logical_Operator_out2206_out1            : std_logic;
  SIGNAL Logical_Operator_out2207_out1            : std_logic;
  SIGNAL Logical_Operator_out2208_out1            : std_logic;
  SIGNAL Logical_Operator_out2209_out1            : std_logic;
  SIGNAL Logical_Operator_out2210_out1            : std_logic;
  SIGNAL Logical_Operator_out2211_out1            : std_logic;
  SIGNAL Logical_Operator_out2212_out1            : std_logic;
  SIGNAL Logical_Operator_out2213_out1            : std_logic;
  SIGNAL Logical_Operator_out2214_out1            : std_logic;
  SIGNAL Logical_Operator_out2215_out1            : std_logic;
  SIGNAL Logical_Operator_out2216_out1            : std_logic;
  SIGNAL Logical_Operator_out2217_out1            : std_logic;
  SIGNAL Logical_Operator_out2218_out1            : std_logic;
  SIGNAL Logical_Operator_out2219_out1            : std_logic;
  SIGNAL Logical_Operator_out2220_out1            : std_logic;
  SIGNAL Logical_Operator_out2221_out1            : std_logic;
  SIGNAL Logical_Operator_out2222_out1            : std_logic;
  SIGNAL Logical_Operator_out2223_out1            : std_logic;
  SIGNAL Logical_Operator_out2224_out1            : std_logic;
  SIGNAL Logical_Operator_out2225_out1            : std_logic;
  SIGNAL Logical_Operator_out2226_out1            : std_logic;
  SIGNAL Logical_Operator_out2227_out1            : std_logic;
  SIGNAL Logical_Operator_out2228_out1            : std_logic;
  SIGNAL Logical_Operator_out2229_out1            : std_logic;
  SIGNAL Logical_Operator_out2230_out1            : std_logic;
  SIGNAL Logical_Operator_out2231_out1            : std_logic;
  SIGNAL Logical_Operator_out2232_out1            : std_logic;
  SIGNAL Logical_Operator_out2233_out1            : std_logic;
  SIGNAL Logical_Operator_out2234_out1            : std_logic;
  SIGNAL Logical_Operator_out2235_out1            : std_logic;
  SIGNAL Logical_Operator_out2236_out1            : std_logic;
  SIGNAL Logical_Operator_out2237_out1            : std_logic;
  SIGNAL Logical_Operator_out2238_out1            : std_logic;
  SIGNAL Logical_Operator_out2239_out1            : std_logic;
  SIGNAL Logical_Operator_out2240_out1            : std_logic;
  SIGNAL Logical_Operator_out2241_out1            : std_logic;
  SIGNAL Logical_Operator_out2242_out1            : std_logic;
  SIGNAL Logical_Operator_out2243_out1            : std_logic;
  SIGNAL Logical_Operator_out2244_out1            : std_logic;
  SIGNAL Logical_Operator_out2245_out1            : std_logic;
  SIGNAL Logical_Operator_out2246_out1            : std_logic;
  SIGNAL Logical_Operator_out2247_out1            : std_logic;
  SIGNAL Logical_Operator_out2248_out1            : std_logic;
  SIGNAL Logical_Operator_out2249_out1            : std_logic;
  SIGNAL Logical_Operator_out2250_out1            : std_logic;
  SIGNAL Logical_Operator_out2251_out1            : std_logic;
  SIGNAL Logical_Operator_out2252_out1            : std_logic;
  SIGNAL Logical_Operator_out2253_out1            : std_logic;
  SIGNAL Logical_Operator_out2254_out1            : std_logic;
  SIGNAL Logical_Operator_out2255_out1            : std_logic;
  SIGNAL Logical_Operator_out2256_out1            : std_logic;
  SIGNAL Logical_Operator_out2257_out1            : std_logic;
  SIGNAL Logical_Operator_out2258_out1            : std_logic;
  SIGNAL Logical_Operator_out2259_out1            : std_logic;
  SIGNAL Logical_Operator_out2260_out1            : std_logic;
  SIGNAL Logical_Operator_out2261_out1            : std_logic;
  SIGNAL Logical_Operator_out2262_out1            : std_logic;
  SIGNAL Logical_Operator_out2263_out1            : std_logic;
  SIGNAL Logical_Operator_out2264_out1            : std_logic;
  SIGNAL Logical_Operator_out2265_out1            : std_logic;
  SIGNAL Logical_Operator_out2266_out1            : std_logic;
  SIGNAL Logical_Operator_out2267_out1            : std_logic;
  SIGNAL Logical_Operator_out2268_out1            : std_logic;
  SIGNAL Logical_Operator_out2269_out1            : std_logic;
  SIGNAL Logical_Operator_out2270_out1            : std_logic;
  SIGNAL Logical_Operator_out2271_out1            : std_logic;
  SIGNAL Logical_Operator_out2272_out1            : std_logic;
  SIGNAL Logical_Operator_out2273_out1            : std_logic;
  SIGNAL Logical_Operator_out2274_out1            : std_logic;
  SIGNAL Logical_Operator_out2275_out1            : std_logic;
  SIGNAL Logical_Operator_out2276_out1            : std_logic;
  SIGNAL Logical_Operator_out2277_out1            : std_logic;
  SIGNAL Logical_Operator_out2278_out1            : std_logic;
  SIGNAL Logical_Operator_out2279_out1            : std_logic;
  SIGNAL Logical_Operator_out2280_out1            : std_logic;
  SIGNAL Logical_Operator_out2281_out1            : std_logic;
  SIGNAL Logical_Operator_out2282_out1            : std_logic;
  SIGNAL Logical_Operator_out2283_out1            : std_logic;
  SIGNAL Logical_Operator_out2284_out1            : std_logic;
  SIGNAL Logical_Operator_out2285_out1            : std_logic;
  SIGNAL Logical_Operator_out2286_out1            : std_logic;
  SIGNAL Logical_Operator_out2287_out1            : std_logic;
  SIGNAL Logical_Operator_out2288_out1            : std_logic;
  SIGNAL Logical_Operator_out2289_out1            : std_logic;
  SIGNAL Logical_Operator_out2290_out1            : std_logic;
  SIGNAL Logical_Operator_out2291_out1            : std_logic;
  SIGNAL Logical_Operator_out2292_out1            : std_logic;
  SIGNAL Logical_Operator_out2293_out1            : std_logic;
  SIGNAL Logical_Operator_out2294_out1            : std_logic;
  SIGNAL Logical_Operator_out2295_out1            : std_logic;
  SIGNAL Logical_Operator_out2296_out1            : std_logic;
  SIGNAL Logical_Operator_out2297_out1            : std_logic;
  SIGNAL Logical_Operator_out2298_out1            : std_logic;
  SIGNAL Logical_Operator_out2299_out1            : std_logic;
  SIGNAL Logical_Operator_out2300_out1            : std_logic;
  SIGNAL Logical_Operator_out2301_out1            : std_logic;
  SIGNAL Logical_Operator_out2302_out1            : std_logic;
  SIGNAL Logical_Operator_out2303_out1            : std_logic;
  SIGNAL Logical_Operator_out2304_out1            : std_logic;
  SIGNAL Logical_Operator_out2305_out1            : std_logic;
  SIGNAL Logical_Operator_out2306_out1            : std_logic;
  SIGNAL Logical_Operator_out2307_out1            : std_logic;
  SIGNAL Logical_Operator_out2308_out1            : std_logic;
  SIGNAL Logical_Operator_out2309_out1            : std_logic;
  SIGNAL Logical_Operator_out2310_out1            : std_logic;
  SIGNAL Logical_Operator_out2311_out1            : std_logic;
  SIGNAL Logical_Operator_out2312_out1            : std_logic;
  SIGNAL Logical_Operator_out2313_out1            : std_logic;
  SIGNAL Logical_Operator_out2314_out1            : std_logic;
  SIGNAL Logical_Operator_out2315_out1            : std_logic;
  SIGNAL Logical_Operator_out2316_out1            : std_logic;
  SIGNAL Logical_Operator_out2317_out1            : std_logic;
  SIGNAL Logical_Operator_out2318_out1            : std_logic;
  SIGNAL Logical_Operator_out2319_out1            : std_logic;
  SIGNAL Logical_Operator_out2320_out1            : std_logic;
  SIGNAL Logical_Operator_out2321_out1            : std_logic;
  SIGNAL Logical_Operator_out2322_out1            : std_logic;
  SIGNAL Logical_Operator_out2323_out1            : std_logic;
  SIGNAL Logical_Operator_out2324_out1            : std_logic;
  SIGNAL Logical_Operator_out2325_out1            : std_logic;
  SIGNAL Logical_Operator_out2326_out1            : std_logic;
  SIGNAL Logical_Operator_out2327_out1            : std_logic;
  SIGNAL Logical_Operator_out2328_out1            : std_logic;
  SIGNAL Logical_Operator_out2329_out1            : std_logic;
  SIGNAL Logical_Operator_out2330_out1            : std_logic;
  SIGNAL Logical_Operator_out2331_out1            : std_logic;
  SIGNAL Logical_Operator_out2332_out1            : std_logic;
  SIGNAL Logical_Operator_out2333_out1            : std_logic;
  SIGNAL Logical_Operator_out2334_out1            : std_logic;
  SIGNAL Logical_Operator_out2335_out1            : std_logic;
  SIGNAL Logical_Operator_out2336_out1            : std_logic;
  SIGNAL Logical_Operator_out2337_out1            : std_logic;
  SIGNAL Logical_Operator_out2338_out1            : std_logic;
  SIGNAL Logical_Operator_out2339_out1            : std_logic;
  SIGNAL Logical_Operator_out2340_out1            : std_logic;
  SIGNAL Logical_Operator_out2341_out1            : std_logic;
  SIGNAL Logical_Operator_out2342_out1            : std_logic;
  SIGNAL Logical_Operator_out2343_out1            : std_logic;
  SIGNAL Logical_Operator_out2344_out1            : std_logic;
  SIGNAL Logical_Operator_out2345_out1            : std_logic;
  SIGNAL Logical_Operator_out2346_out1            : std_logic;
  SIGNAL Logical_Operator_out2347_out1            : std_logic;
  SIGNAL Logical_Operator_out2348_out1            : std_logic;
  SIGNAL Logical_Operator_out2349_out1            : std_logic;
  SIGNAL Logical_Operator_out2350_out1            : std_logic;
  SIGNAL Logical_Operator_out2351_out1            : std_logic;
  SIGNAL Logical_Operator_out2352_out1            : std_logic;
  SIGNAL Logical_Operator_out2353_out1            : std_logic;
  SIGNAL Logical_Operator_out2354_out1            : std_logic;
  SIGNAL Logical_Operator_out2355_out1            : std_logic;
  SIGNAL Logical_Operator_out2356_out1            : std_logic;
  SIGNAL Logical_Operator_out2357_out1            : std_logic;
  SIGNAL Logical_Operator_out2358_out1            : std_logic;
  SIGNAL Logical_Operator_out2359_out1            : std_logic;
  SIGNAL Logical_Operator_out2360_out1            : std_logic;
  SIGNAL Logical_Operator_out2361_out1            : std_logic;
  SIGNAL Logical_Operator_out2362_out1            : std_logic;
  SIGNAL Logical_Operator_out2363_out1            : std_logic;
  SIGNAL Logical_Operator_out2364_out1            : std_logic;
  SIGNAL Logical_Operator_out2365_out1            : std_logic;
  SIGNAL Logical_Operator_out2366_out1            : std_logic;
  SIGNAL Logical_Operator_out2367_out1            : std_logic;
  SIGNAL Logical_Operator_out2368_out1            : std_logic;
  SIGNAL Logical_Operator_out2369_out1            : std_logic;
  SIGNAL Logical_Operator_out2370_out1            : std_logic;
  SIGNAL Logical_Operator_out2371_out1            : std_logic;
  SIGNAL Logical_Operator_out2372_out1            : std_logic;
  SIGNAL Logical_Operator_out2373_out1            : std_logic;
  SIGNAL Logical_Operator_out2374_out1            : std_logic;
  SIGNAL Logical_Operator_out2375_out1            : std_logic;
  SIGNAL Logical_Operator_out2376_out1            : std_logic;
  SIGNAL Logical_Operator_out2377_out1            : std_logic;
  SIGNAL Logical_Operator_out2378_out1            : std_logic;
  SIGNAL Logical_Operator_out2379_out1            : std_logic;
  SIGNAL Logical_Operator_out2380_out1            : std_logic;
  SIGNAL Logical_Operator_out2381_out1            : std_logic;
  SIGNAL Logical_Operator_out2382_out1            : std_logic;
  SIGNAL Logical_Operator_out2383_out1            : std_logic;
  SIGNAL Logical_Operator_out2384_out1            : std_logic;
  SIGNAL Logical_Operator_out2385_out1            : std_logic;
  SIGNAL Logical_Operator_out2386_out1            : std_logic;
  SIGNAL Logical_Operator_out2387_out1            : std_logic;
  SIGNAL Logical_Operator_out2388_out1            : std_logic;
  SIGNAL Logical_Operator_out2389_out1            : std_logic;
  SIGNAL Logical_Operator_out2390_out1            : std_logic;
  SIGNAL Logical_Operator_out2391_out1            : std_logic;
  SIGNAL Logical_Operator_out2392_out1            : std_logic;
  SIGNAL Logical_Operator_out2393_out1            : std_logic;
  SIGNAL Logical_Operator_out2394_out1            : std_logic;
  SIGNAL Logical_Operator_out2395_out1            : std_logic;
  SIGNAL Logical_Operator_out2396_out1            : std_logic;
  SIGNAL Logical_Operator_out2397_out1            : std_logic;
  SIGNAL Logical_Operator_out2398_out1            : std_logic;
  SIGNAL Logical_Operator_out2399_out1            : std_logic;
  SIGNAL Logical_Operator_out2400_out1            : std_logic;
  SIGNAL Logical_Operator_out2401_out1            : std_logic;
  SIGNAL Logical_Operator_out2402_out1            : std_logic;
  SIGNAL Logical_Operator_out2403_out1            : std_logic;
  SIGNAL Logical_Operator_out2404_out1            : std_logic;
  SIGNAL Logical_Operator_out2405_out1            : std_logic;
  SIGNAL Logical_Operator_out2406_out1            : std_logic;
  SIGNAL Logical_Operator_out2407_out1            : std_logic;
  SIGNAL Logical_Operator_out2408_out1            : std_logic;
  SIGNAL Logical_Operator_out2409_out1            : std_logic;
  SIGNAL Logical_Operator_out2410_out1            : std_logic;
  SIGNAL Logical_Operator_out2411_out1            : std_logic;
  SIGNAL Logical_Operator_out2412_out1            : std_logic;
  SIGNAL Logical_Operator_out2413_out1            : std_logic;
  SIGNAL Logical_Operator_out2414_out1            : std_logic;
  SIGNAL Logical_Operator_out2415_out1            : std_logic;
  SIGNAL Logical_Operator_out2416_out1            : std_logic;
  SIGNAL Logical_Operator_out2417_out1            : std_logic;
  SIGNAL Logical_Operator_out2418_out1            : std_logic;
  SIGNAL Logical_Operator_out2419_out1            : std_logic;
  SIGNAL Logical_Operator_out2420_out1            : std_logic;
  SIGNAL Logical_Operator_out2421_out1            : std_logic;
  SIGNAL Logical_Operator_out2422_out1            : std_logic;
  SIGNAL Logical_Operator_out2423_out1            : std_logic;
  SIGNAL Logical_Operator_out2424_out1            : std_logic;
  SIGNAL Logical_Operator_out2425_out1            : std_logic;
  SIGNAL Logical_Operator_out2426_out1            : std_logic;
  SIGNAL Logical_Operator_out2427_out1            : std_logic;
  SIGNAL Logical_Operator_out2428_out1            : std_logic;
  SIGNAL Logical_Operator_out2429_out1            : std_logic;
  SIGNAL Logical_Operator_out2430_out1            : std_logic;
  SIGNAL Logical_Operator_out2431_out1            : std_logic;
  SIGNAL Logical_Operator_out2432_out1            : std_logic;
  SIGNAL Logical_Operator_out2433_out1            : std_logic;
  SIGNAL Logical_Operator_out2434_out1            : std_logic;
  SIGNAL Logical_Operator_out2435_out1            : std_logic;
  SIGNAL Logical_Operator_out2436_out1            : std_logic;
  SIGNAL Logical_Operator_out2437_out1            : std_logic;
  SIGNAL Logical_Operator_out2438_out1            : std_logic;
  SIGNAL Logical_Operator_out2439_out1            : std_logic;
  SIGNAL Logical_Operator_out2440_out1            : std_logic;
  SIGNAL Logical_Operator_out2441_out1            : std_logic;
  SIGNAL Logical_Operator_out2442_out1            : std_logic;
  SIGNAL Logical_Operator_out2443_out1            : std_logic;
  SIGNAL Logical_Operator_out2444_out1            : std_logic;
  SIGNAL Logical_Operator_out2445_out1            : std_logic;
  SIGNAL Logical_Operator_out2446_out1            : std_logic;
  SIGNAL Logical_Operator_out2447_out1            : std_logic;
  SIGNAL Logical_Operator_out2448_out1            : std_logic;
  SIGNAL Logical_Operator_out2449_out1            : std_logic;
  SIGNAL Logical_Operator_out2450_out1            : std_logic;
  SIGNAL Logical_Operator_out2451_out1            : std_logic;
  SIGNAL Logical_Operator_out2452_out1            : std_logic;
  SIGNAL Logical_Operator_out2453_out1            : std_logic;
  SIGNAL Logical_Operator_out2454_out1            : std_logic;
  SIGNAL Logical_Operator_out2455_out1            : std_logic;
  SIGNAL Logical_Operator_out2456_out1            : std_logic;
  SIGNAL Logical_Operator_out2457_out1            : std_logic;
  SIGNAL Logical_Operator_out2458_out1            : std_logic;
  SIGNAL Logical_Operator_out2459_out1            : std_logic;
  SIGNAL Logical_Operator_out2460_out1            : std_logic;
  SIGNAL Logical_Operator_out2461_out1            : std_logic;
  SIGNAL Logical_Operator_out2462_out1            : std_logic;
  SIGNAL Logical_Operator_out2463_out1            : std_logic;
  SIGNAL Logical_Operator_out2464_out1            : std_logic;
  SIGNAL Logical_Operator_out2465_out1            : std_logic;
  SIGNAL Logical_Operator_out2466_out1            : std_logic;
  SIGNAL Logical_Operator_out2467_out1            : std_logic;
  SIGNAL Logical_Operator_out2468_out1            : std_logic;
  SIGNAL Logical_Operator_out2469_out1            : std_logic;
  SIGNAL Logical_Operator_out2470_out1            : std_logic;
  SIGNAL Logical_Operator_out2471_out1            : std_logic;
  SIGNAL Logical_Operator_out2472_out1            : std_logic;
  SIGNAL Logical_Operator_out2473_out1            : std_logic;
  SIGNAL Logical_Operator_out2474_out1            : std_logic;
  SIGNAL Logical_Operator_out2475_out1            : std_logic;
  SIGNAL Logical_Operator_out2476_out1            : std_logic;
  SIGNAL Logical_Operator_out2477_out1            : std_logic;
  SIGNAL Logical_Operator_out2478_out1            : std_logic;
  SIGNAL Logical_Operator_out2479_out1            : std_logic;
  SIGNAL Logical_Operator_out2480_out1            : std_logic;
  SIGNAL Logical_Operator_out2481_out1            : std_logic;
  SIGNAL Logical_Operator_out2482_out1            : std_logic;
  SIGNAL Logical_Operator_out2483_out1            : std_logic;
  SIGNAL Logical_Operator_out2484_out1            : std_logic;
  SIGNAL Logical_Operator_out2485_out1            : std_logic;
  SIGNAL Logical_Operator_out2486_out1            : std_logic;
  SIGNAL Logical_Operator_out2487_out1            : std_logic;
  SIGNAL Logical_Operator_out2488_out1            : std_logic;
  SIGNAL Logical_Operator_out2489_out1            : std_logic;
  SIGNAL Logical_Operator_out2490_out1            : std_logic;
  SIGNAL Logical_Operator_out2491_out1            : std_logic;
  SIGNAL Logical_Operator_out2492_out1            : std_logic;
  SIGNAL Logical_Operator_out2493_out1            : std_logic;
  SIGNAL Logical_Operator_out2494_out1            : std_logic;
  SIGNAL Logical_Operator_out2495_out1            : std_logic;
  SIGNAL Logical_Operator_out2496_out1            : std_logic;
  SIGNAL Logical_Operator_out2497_out1            : std_logic;
  SIGNAL Logical_Operator_out2498_out1            : std_logic;
  SIGNAL Logical_Operator_out2499_out1            : std_logic;
  SIGNAL Logical_Operator_out2500_out1            : std_logic;
  SIGNAL Logical_Operator_out2501_out1            : std_logic;
  SIGNAL Logical_Operator_out2502_out1            : std_logic;
  SIGNAL Logical_Operator_out2503_out1            : std_logic;
  SIGNAL Logical_Operator_out2504_out1            : std_logic;
  SIGNAL Logical_Operator_out2505_out1            : std_logic;
  SIGNAL Logical_Operator_out2506_out1            : std_logic;
  SIGNAL Logical_Operator_out2507_out1            : std_logic;
  SIGNAL Logical_Operator_out2508_out1            : std_logic;
  SIGNAL Logical_Operator_out2509_out1            : std_logic;
  SIGNAL Logical_Operator_out2510_out1            : std_logic;
  SIGNAL Logical_Operator_out2511_out1            : std_logic;
  SIGNAL Logical_Operator_out2512_out1            : std_logic;
  SIGNAL Logical_Operator_out2513_out1            : std_logic;
  SIGNAL Logical_Operator_out2514_out1            : std_logic;
  SIGNAL Logical_Operator_out2515_out1            : std_logic;
  SIGNAL Logical_Operator_out2516_out1            : std_logic;
  SIGNAL Logical_Operator_out2517_out1            : std_logic;
  SIGNAL Logical_Operator_out2518_out1            : std_logic;
  SIGNAL Logical_Operator_out2519_out1            : std_logic;
  SIGNAL Logical_Operator_out2520_out1            : std_logic;
  SIGNAL Logical_Operator_out2521_out1            : std_logic;
  SIGNAL Logical_Operator_out2522_out1            : std_logic;
  SIGNAL Logical_Operator_out2523_out1            : std_logic;
  SIGNAL Logical_Operator_out2524_out1            : std_logic;
  SIGNAL Logical_Operator_out2525_out1            : std_logic;
  SIGNAL Logical_Operator_out2526_out1            : std_logic;
  SIGNAL Logical_Operator_out2527_out1            : std_logic;
  SIGNAL Logical_Operator_out2528_out1            : std_logic;
  SIGNAL Logical_Operator_out2529_out1            : std_logic;
  SIGNAL Logical_Operator_out2530_out1            : std_logic;
  SIGNAL Logical_Operator_out2531_out1            : std_logic;
  SIGNAL Logical_Operator_out2532_out1            : std_logic;
  SIGNAL Logical_Operator_out2533_out1            : std_logic;
  SIGNAL Logical_Operator_out2534_out1            : std_logic;
  SIGNAL Logical_Operator_out2535_out1            : std_logic;
  SIGNAL Logical_Operator_out2536_out1            : std_logic;
  SIGNAL Logical_Operator_out2537_out1            : std_logic;
  SIGNAL Logical_Operator_out2538_out1            : std_logic;
  SIGNAL Logical_Operator_out2539_out1            : std_logic;
  SIGNAL Logical_Operator_out2540_out1            : std_logic;
  SIGNAL Logical_Operator_out2541_out1            : std_logic;
  SIGNAL Logical_Operator_out2542_out1            : std_logic;
  SIGNAL Logical_Operator_out2543_out1            : std_logic;
  SIGNAL Logical_Operator_out2544_out1            : std_logic;
  SIGNAL Logical_Operator_out2545_out1            : std_logic;
  SIGNAL Logical_Operator_out2546_out1            : std_logic;
  SIGNAL Logical_Operator_out2547_out1            : std_logic;
  SIGNAL Logical_Operator_out2548_out1            : std_logic;
  SIGNAL Logical_Operator_out2549_out1            : std_logic;
  SIGNAL Logical_Operator_out2550_out1            : std_logic;
  SIGNAL Logical_Operator_out2551_out1            : std_logic;
  SIGNAL Logical_Operator_out2552_out1            : std_logic;
  SIGNAL Logical_Operator_out2553_out1            : std_logic;
  SIGNAL Logical_Operator_out2554_out1            : std_logic;
  SIGNAL Logical_Operator_out2555_out1            : std_logic;
  SIGNAL Logical_Operator_out2556_out1            : std_logic;
  SIGNAL Logical_Operator_out2557_out1            : std_logic;
  SIGNAL Logical_Operator_out2558_out1            : std_logic;
  SIGNAL Logical_Operator_out2559_out1            : std_logic;
  SIGNAL Logical_Operator_out2560_out1            : std_logic;
  SIGNAL Logical_Operator_out2561_out1            : std_logic;
  SIGNAL Logical_Operator_out2562_out1            : std_logic;
  SIGNAL Logical_Operator_out2563_out1            : std_logic;
  SIGNAL Logical_Operator_out2564_out1            : std_logic;
  SIGNAL Logical_Operator_out2565_out1            : std_logic;
  SIGNAL Logical_Operator_out2566_out1            : std_logic;
  SIGNAL Logical_Operator_out2567_out1            : std_logic;
  SIGNAL Logical_Operator_out2568_out1            : std_logic;
  SIGNAL Logical_Operator_out2569_out1            : std_logic;
  SIGNAL Logical_Operator_out2570_out1            : std_logic;
  SIGNAL Logical_Operator_out2571_out1            : std_logic;
  SIGNAL Logical_Operator_out2572_out1            : std_logic;
  SIGNAL Logical_Operator_out2573_out1            : std_logic;
  SIGNAL Logical_Operator_out2574_out1            : std_logic;
  SIGNAL Logical_Operator_out2575_out1            : std_logic;
  SIGNAL Logical_Operator_out2576_out1            : std_logic;
  SIGNAL Logical_Operator_out2577_out1            : std_logic;
  SIGNAL Logical_Operator_out2578_out1            : std_logic;
  SIGNAL Logical_Operator_out2579_out1            : std_logic;
  SIGNAL Logical_Operator_out2580_out1            : std_logic;
  SIGNAL Logical_Operator_out2581_out1            : std_logic;
  SIGNAL Logical_Operator_out2582_out1            : std_logic;
  SIGNAL Logical_Operator_out2583_out1            : std_logic;
  SIGNAL Logical_Operator_out2584_out1            : std_logic;
  SIGNAL Logical_Operator_out2585_out1            : std_logic;
  SIGNAL Logical_Operator_out2586_out1            : std_logic;
  SIGNAL Logical_Operator_out2587_out1            : std_logic;
  SIGNAL Logical_Operator_out2588_out1            : std_logic;
  SIGNAL Logical_Operator_out2589_out1            : std_logic;
  SIGNAL Logical_Operator_out2590_out1            : std_logic;
  SIGNAL Logical_Operator_out2591_out1            : std_logic;
  SIGNAL Logical_Operator_out2592_out1            : std_logic;
  SIGNAL Logical_Operator_out2593_out1            : std_logic;
  SIGNAL Logical_Operator_out2594_out1            : std_logic;
  SIGNAL Logical_Operator_out2595_out1            : std_logic;
  SIGNAL Logical_Operator_out2596_out1            : std_logic;
  SIGNAL Logical_Operator_out2597_out1            : std_logic;
  SIGNAL Logical_Operator_out2598_out1            : std_logic;
  SIGNAL Logical_Operator_out2599_out1            : std_logic;
  SIGNAL Logical_Operator_out2600_out1            : std_logic;
  SIGNAL Logical_Operator_out2601_out1            : std_logic;
  SIGNAL Logical_Operator_out2602_out1            : std_logic;
  SIGNAL Logical_Operator_out2603_out1            : std_logic;
  SIGNAL Logical_Operator_out2604_out1            : std_logic;
  SIGNAL Logical_Operator_out2605_out1            : std_logic;
  SIGNAL Logical_Operator_out2606_out1            : std_logic;
  SIGNAL Logical_Operator_out2607_out1            : std_logic;
  SIGNAL Logical_Operator_out2608_out1            : std_logic;
  SIGNAL Logical_Operator_out2609_out1            : std_logic;
  SIGNAL Logical_Operator_out2610_out1            : std_logic;
  SIGNAL Logical_Operator_out2611_out1            : std_logic;
  SIGNAL Logical_Operator_out2612_out1            : std_logic;
  SIGNAL Logical_Operator_out2613_out1            : std_logic;
  SIGNAL Logical_Operator_out2614_out1            : std_logic;
  SIGNAL Logical_Operator_out2615_out1            : std_logic;
  SIGNAL Logical_Operator_out2616_out1            : std_logic;
  SIGNAL Logical_Operator_out2617_out1            : std_logic;
  SIGNAL Logical_Operator_out2618_out1            : std_logic;
  SIGNAL Logical_Operator_out2619_out1            : std_logic;
  SIGNAL Logical_Operator_out2620_out1            : std_logic;
  SIGNAL Logical_Operator_out2621_out1            : std_logic;
  SIGNAL Logical_Operator_out2622_out1            : std_logic;
  SIGNAL Logical_Operator_out2623_out1            : std_logic;
  SIGNAL Logical_Operator_out2624_out1            : std_logic;
  SIGNAL Logical_Operator_out2625_out1            : std_logic;
  SIGNAL Logical_Operator_out2626_out1            : std_logic;
  SIGNAL Logical_Operator_out2627_out1            : std_logic;
  SIGNAL Logical_Operator_out2628_out1            : std_logic;
  SIGNAL Logical_Operator_out2629_out1            : std_logic;
  SIGNAL Logical_Operator_out2630_out1            : std_logic;
  SIGNAL Logical_Operator_out2631_out1            : std_logic;
  SIGNAL Logical_Operator_out2632_out1            : std_logic;
  SIGNAL Logical_Operator_out2633_out1            : std_logic;
  SIGNAL Logical_Operator_out2634_out1            : std_logic;
  SIGNAL Logical_Operator_out2635_out1            : std_logic;
  SIGNAL Logical_Operator_out2636_out1            : std_logic;
  SIGNAL Logical_Operator_out2637_out1            : std_logic;
  SIGNAL Logical_Operator_out2638_out1            : std_logic;
  SIGNAL Logical_Operator_out2639_out1            : std_logic;
  SIGNAL Logical_Operator_out2640_out1            : std_logic;
  SIGNAL Logical_Operator_out2641_out1            : std_logic;
  SIGNAL Logical_Operator_out2642_out1            : std_logic;
  SIGNAL Logical_Operator_out2643_out1            : std_logic;
  SIGNAL Logical_Operator_out2644_out1            : std_logic;
  SIGNAL Logical_Operator_out2645_out1            : std_logic;
  SIGNAL Logical_Operator_out2646_out1            : std_logic;
  SIGNAL Logical_Operator_out2647_out1            : std_logic;
  SIGNAL Logical_Operator_out2648_out1            : std_logic;
  SIGNAL Logical_Operator_out2649_out1            : std_logic;
  SIGNAL Logical_Operator_out2650_out1            : std_logic;
  SIGNAL Logical_Operator_out2651_out1            : std_logic;
  SIGNAL Logical_Operator_out2652_out1            : std_logic;
  SIGNAL Logical_Operator_out2653_out1            : std_logic;
  SIGNAL Logical_Operator_out2654_out1            : std_logic;
  SIGNAL Logical_Operator_out2655_out1            : std_logic;
  SIGNAL Logical_Operator_out2656_out1            : std_logic;
  SIGNAL Logical_Operator_out2657_out1            : std_logic;
  SIGNAL Logical_Operator_out2658_out1            : std_logic;
  SIGNAL Logical_Operator_out2659_out1            : std_logic;
  SIGNAL Logical_Operator_out2660_out1            : std_logic;
  SIGNAL Logical_Operator_out2661_out1            : std_logic;
  SIGNAL Logical_Operator_out2662_out1            : std_logic;
  SIGNAL Logical_Operator_out2663_out1            : std_logic;
  SIGNAL Logical_Operator_out2664_out1            : std_logic;
  SIGNAL Logical_Operator_out2665_out1            : std_logic;
  SIGNAL Logical_Operator_out2666_out1            : std_logic;
  SIGNAL Logical_Operator_out2667_out1            : std_logic;
  SIGNAL Logical_Operator_out2668_out1            : std_logic;
  SIGNAL Logical_Operator_out2669_out1            : std_logic;
  SIGNAL Logical_Operator_out2670_out1            : std_logic;
  SIGNAL Logical_Operator_out2671_out1            : std_logic;
  SIGNAL Logical_Operator_out2672_out1            : std_logic;
  SIGNAL Logical_Operator_out2673_out1            : std_logic;
  SIGNAL Logical_Operator_out2674_out1            : std_logic;
  SIGNAL Logical_Operator_out2675_out1            : std_logic;
  SIGNAL Logical_Operator_out2676_out1            : std_logic;
  SIGNAL Logical_Operator_out2677_out1            : std_logic;
  SIGNAL Logical_Operator_out2678_out1            : std_logic;
  SIGNAL Logical_Operator_out2679_out1            : std_logic;
  SIGNAL Logical_Operator_out2680_out1            : std_logic;
  SIGNAL Logical_Operator_out2681_out1            : std_logic;
  SIGNAL Logical_Operator_out2682_out1            : std_logic;
  SIGNAL Logical_Operator_out2683_out1            : std_logic;
  SIGNAL Logical_Operator_out2684_out1            : std_logic;
  SIGNAL Logical_Operator_out2685_out1            : std_logic;
  SIGNAL Logical_Operator_out2686_out1            : std_logic;
  SIGNAL Logical_Operator_out2687_out1            : std_logic;
  SIGNAL Logical_Operator_out2688_out1            : std_logic;
  SIGNAL Logical_Operator_out2689_out1            : std_logic;
  SIGNAL Logical_Operator_out2690_out1            : std_logic;
  SIGNAL Logical_Operator_out2691_out1            : std_logic;
  SIGNAL Logical_Operator_out2692_out1            : std_logic;
  SIGNAL Logical_Operator_out2693_out1            : std_logic;
  SIGNAL Logical_Operator_out2694_out1            : std_logic;
  SIGNAL Logical_Operator_out2695_out1            : std_logic;
  SIGNAL Logical_Operator_out2696_out1            : std_logic;
  SIGNAL Logical_Operator_out2697_out1            : std_logic;
  SIGNAL Logical_Operator_out2698_out1            : std_logic;
  SIGNAL Logical_Operator_out2699_out1            : std_logic;
  SIGNAL Logical_Operator_out2700_out1            : std_logic;
  SIGNAL Logical_Operator_out2701_out1            : std_logic;
  SIGNAL Logical_Operator_out2702_out1            : std_logic;
  SIGNAL Logical_Operator_out2703_out1            : std_logic;
  SIGNAL Logical_Operator_out2704_out1            : std_logic;
  SIGNAL Logical_Operator_out2705_out1            : std_logic;
  SIGNAL Logical_Operator_out2706_out1            : std_logic;
  SIGNAL Logical_Operator_out2707_out1            : std_logic;
  SIGNAL Logical_Operator_out2708_out1            : std_logic;
  SIGNAL Logical_Operator_out2709_out1            : std_logic;
  SIGNAL Logical_Operator_out2710_out1            : std_logic;
  SIGNAL Logical_Operator_out2711_out1            : std_logic;
  SIGNAL Logical_Operator_out2712_out1            : std_logic;
  SIGNAL Logical_Operator_out2713_out1            : std_logic;
  SIGNAL Logical_Operator_out2714_out1            : std_logic;
  SIGNAL Logical_Operator_out2715_out1            : std_logic;
  SIGNAL Logical_Operator_out2716_out1            : std_logic;
  SIGNAL Logical_Operator_out2717_out1            : std_logic;
  SIGNAL Logical_Operator_out2718_out1            : std_logic;
  SIGNAL Logical_Operator_out2719_out1            : std_logic;
  SIGNAL Logical_Operator_out2720_out1            : std_logic;
  SIGNAL Logical_Operator_out2721_out1            : std_logic;
  SIGNAL Logical_Operator_out2722_out1            : std_logic;
  SIGNAL Logical_Operator_out2723_out1            : std_logic;
  SIGNAL Logical_Operator_out2724_out1            : std_logic;
  SIGNAL Logical_Operator_out2725_out1            : std_logic;
  SIGNAL Logical_Operator_out2726_out1            : std_logic;
  SIGNAL Logical_Operator_out2727_out1            : std_logic;
  SIGNAL Logical_Operator_out2728_out1            : std_logic;
  SIGNAL Logical_Operator_out2729_out1            : std_logic;
  SIGNAL Logical_Operator_out2730_out1            : std_logic;
  SIGNAL Logical_Operator_out2731_out1            : std_logic;
  SIGNAL Logical_Operator_out2732_out1            : std_logic;
  SIGNAL Logical_Operator_out2733_out1            : std_logic;
  SIGNAL Logical_Operator_out2734_out1            : std_logic;
  SIGNAL Logical_Operator_out2735_out1            : std_logic;
  SIGNAL Logical_Operator_out2736_out1            : std_logic;
  SIGNAL Logical_Operator_out2737_out1            : std_logic;
  SIGNAL Logical_Operator_out2738_out1            : std_logic;
  SIGNAL Logical_Operator_out2739_out1            : std_logic;
  SIGNAL Logical_Operator_out2740_out1            : std_logic;
  SIGNAL Logical_Operator_out2741_out1            : std_logic;
  SIGNAL Logical_Operator_out2742_out1            : std_logic;
  SIGNAL Logical_Operator_out2743_out1            : std_logic;
  SIGNAL Logical_Operator_out2744_out1            : std_logic;
  SIGNAL Logical_Operator_out2745_out1            : std_logic;
  SIGNAL Logical_Operator_out2746_out1            : std_logic;
  SIGNAL Logical_Operator_out2747_out1            : std_logic;
  SIGNAL Logical_Operator_out2748_out1            : std_logic;
  SIGNAL Logical_Operator_out2749_out1            : std_logic;
  SIGNAL Logical_Operator_out2750_out1            : std_logic;
  SIGNAL Logical_Operator_out2751_out1            : std_logic;
  SIGNAL Logical_Operator_out2752_out1            : std_logic;
  SIGNAL Logical_Operator_out2753_out1            : std_logic;
  SIGNAL Logical_Operator_out2754_out1            : std_logic;
  SIGNAL Logical_Operator_out2755_out1            : std_logic;
  SIGNAL Logical_Operator_out2756_out1            : std_logic;
  SIGNAL Logical_Operator_out2757_out1            : std_logic;
  SIGNAL Logical_Operator_out2758_out1            : std_logic;
  SIGNAL Logical_Operator_out2759_out1            : std_logic;
  SIGNAL Logical_Operator_out2760_out1            : std_logic;
  SIGNAL Logical_Operator_out2761_out1            : std_logic;
  SIGNAL Logical_Operator_out2762_out1            : std_logic;
  SIGNAL Logical_Operator_out2763_out1            : std_logic;
  SIGNAL Logical_Operator_out2764_out1            : std_logic;
  SIGNAL Logical_Operator_out2765_out1            : std_logic;
  SIGNAL Logical_Operator_out2766_out1            : std_logic;
  SIGNAL Logical_Operator_out2767_out1            : std_logic;
  SIGNAL Logical_Operator_out2768_out1            : std_logic;
  SIGNAL Logical_Operator_out2769_out1            : std_logic;
  SIGNAL Logical_Operator_out2770_out1            : std_logic;
  SIGNAL Logical_Operator_out2771_out1            : std_logic;
  SIGNAL Logical_Operator_out2772_out1            : std_logic;
  SIGNAL Logical_Operator_out2773_out1            : std_logic;
  SIGNAL Logical_Operator_out2774_out1            : std_logic;
  SIGNAL Logical_Operator_out2775_out1            : std_logic;
  SIGNAL Logical_Operator_out2776_out1            : std_logic;
  SIGNAL Logical_Operator_out2777_out1            : std_logic;
  SIGNAL Logical_Operator_out2778_out1            : std_logic;
  SIGNAL Logical_Operator_out2779_out1            : std_logic;
  SIGNAL Logical_Operator_out2780_out1            : std_logic;
  SIGNAL Logical_Operator_out2781_out1            : std_logic;
  SIGNAL Logical_Operator_out2782_out1            : std_logic;
  SIGNAL Logical_Operator_out2783_out1            : std_logic;
  SIGNAL Logical_Operator_out2784_out1            : std_logic;
  SIGNAL Logical_Operator_out2785_out1            : std_logic;
  SIGNAL Logical_Operator_out2786_out1            : std_logic;
  SIGNAL Logical_Operator_out2787_out1            : std_logic;
  SIGNAL Logical_Operator_out2788_out1            : std_logic;
  SIGNAL Logical_Operator_out2789_out1            : std_logic;
  SIGNAL Logical_Operator_out2790_out1            : std_logic;
  SIGNAL Logical_Operator_out2791_out1            : std_logic;
  SIGNAL Logical_Operator_out2792_out1            : std_logic;
  SIGNAL Logical_Operator_out2793_out1            : std_logic;
  SIGNAL Logical_Operator_out2794_out1            : std_logic;
  SIGNAL Logical_Operator_out2795_out1            : std_logic;
  SIGNAL Logical_Operator_out2796_out1            : std_logic;
  SIGNAL Logical_Operator_out2797_out1            : std_logic;
  SIGNAL Logical_Operator_out2798_out1            : std_logic;
  SIGNAL Logical_Operator_out2799_out1            : std_logic;
  SIGNAL Logical_Operator_out2800_out1            : std_logic;
  SIGNAL Logical_Operator_out2801_out1            : std_logic;
  SIGNAL Logical_Operator_out2802_out1            : std_logic;
  SIGNAL Logical_Operator_out2803_out1            : std_logic;
  SIGNAL Logical_Operator_out2804_out1            : std_logic;
  SIGNAL Logical_Operator_out2805_out1            : std_logic;
  SIGNAL Logical_Operator_out2806_out1            : std_logic;
  SIGNAL Logical_Operator_out2807_out1            : std_logic;
  SIGNAL Logical_Operator_out2808_out1            : std_logic;
  SIGNAL Logical_Operator_out2809_out1            : std_logic;
  SIGNAL Logical_Operator_out2810_out1            : std_logic;
  SIGNAL Logical_Operator_out2811_out1            : std_logic;
  SIGNAL Logical_Operator_out2812_out1            : std_logic;
  SIGNAL Logical_Operator_out2813_out1            : std_logic;
  SIGNAL Logical_Operator_out2814_out1            : std_logic;
  SIGNAL Logical_Operator_out2815_out1            : std_logic;
  SIGNAL Logical_Operator_out2816_out1            : std_logic;
  SIGNAL Logical_Operator_out2817_out1            : std_logic;
  SIGNAL Logical_Operator_out2818_out1            : std_logic;
  SIGNAL Logical_Operator_out2819_out1            : std_logic;
  SIGNAL Logical_Operator_out2820_out1            : std_logic;
  SIGNAL Logical_Operator_out2821_out1            : std_logic;
  SIGNAL Logical_Operator_out2822_out1            : std_logic;
  SIGNAL Logical_Operator_out2823_out1            : std_logic;
  SIGNAL Logical_Operator_out2824_out1            : std_logic;
  SIGNAL Logical_Operator_out2825_out1            : std_logic;
  SIGNAL Logical_Operator_out2826_out1            : std_logic;
  SIGNAL Logical_Operator_out2827_out1            : std_logic;
  SIGNAL Logical_Operator_out2828_out1            : std_logic;
  SIGNAL Logical_Operator_out2829_out1            : std_logic;
  SIGNAL Logical_Operator_out2830_out1            : std_logic;
  SIGNAL Logical_Operator_out2831_out1            : std_logic;
  SIGNAL Logical_Operator_out2832_out1            : std_logic;
  SIGNAL Logical_Operator_out2833_out1            : std_logic;
  SIGNAL Logical_Operator_out2834_out1            : std_logic;
  SIGNAL Logical_Operator_out2835_out1            : std_logic;
  SIGNAL Logical_Operator_out2836_out1            : std_logic;
  SIGNAL Logical_Operator_out2837_out1            : std_logic;
  SIGNAL Logical_Operator_out2838_out1            : std_logic;
  SIGNAL Logical_Operator_out2839_out1            : std_logic;
  SIGNAL Logical_Operator_out2840_out1            : std_logic;
  SIGNAL Logical_Operator_out2841_out1            : std_logic;
  SIGNAL Logical_Operator_out2842_out1            : std_logic;
  SIGNAL Logical_Operator_out2843_out1            : std_logic;
  SIGNAL Logical_Operator_out2844_out1            : std_logic;
  SIGNAL Logical_Operator_out2845_out1            : std_logic;
  SIGNAL Logical_Operator_out2846_out1            : std_logic;
  SIGNAL Logical_Operator_out2847_out1            : std_logic;
  SIGNAL Logical_Operator_out2848_out1            : std_logic;
  SIGNAL Logical_Operator_out2849_out1            : std_logic;
  SIGNAL Logical_Operator_out2850_out1            : std_logic;
  SIGNAL Logical_Operator_out2851_out1            : std_logic;
  SIGNAL Logical_Operator_out2852_out1            : std_logic;
  SIGNAL Logical_Operator_out2853_out1            : std_logic;
  SIGNAL Logical_Operator_out2854_out1            : std_logic;
  SIGNAL Logical_Operator_out2855_out1            : std_logic;
  SIGNAL Logical_Operator_out2856_out1            : std_logic;
  SIGNAL Logical_Operator_out2857_out1            : std_logic;
  SIGNAL Logical_Operator_out2858_out1            : std_logic;
  SIGNAL Logical_Operator_out2859_out1            : std_logic;
  SIGNAL Logical_Operator_out2860_out1            : std_logic;
  SIGNAL Logical_Operator_out2861_out1            : std_logic;
  SIGNAL Logical_Operator_out2862_out1            : std_logic;
  SIGNAL Logical_Operator_out2863_out1            : std_logic;
  SIGNAL Logical_Operator_out2864_out1            : std_logic;
  SIGNAL Logical_Operator_out2865_out1            : std_logic;
  SIGNAL Logical_Operator_out2866_out1            : std_logic;
  SIGNAL Logical_Operator_out2867_out1            : std_logic;
  SIGNAL Logical_Operator_out2868_out1            : std_logic;
  SIGNAL Logical_Operator_out2869_out1            : std_logic;
  SIGNAL Logical_Operator_out2870_out1            : std_logic;
  SIGNAL Logical_Operator_out2871_out1            : std_logic;
  SIGNAL Logical_Operator_out2872_out1            : std_logic;
  SIGNAL Logical_Operator_out2873_out1            : std_logic;
  SIGNAL Logical_Operator_out2874_out1            : std_logic;
  SIGNAL Logical_Operator_out2875_out1            : std_logic;
  SIGNAL Logical_Operator_out2876_out1            : std_logic;
  SIGNAL Logical_Operator_out2877_out1            : std_logic;
  SIGNAL Logical_Operator_out2878_out1            : std_logic;
  SIGNAL Logical_Operator_out2879_out1            : std_logic;
  SIGNAL Logical_Operator_out2880_out1            : std_logic;
  SIGNAL Logical_Operator_out2881_out1            : std_logic;
  SIGNAL Logical_Operator_out2882_out1            : std_logic;
  SIGNAL Logical_Operator_out2883_out1            : std_logic;
  SIGNAL Logical_Operator_out2884_out1            : std_logic;
  SIGNAL Logical_Operator_out2885_out1            : std_logic;
  SIGNAL Logical_Operator_out2886_out1            : std_logic;
  SIGNAL Logical_Operator_out2887_out1            : std_logic;
  SIGNAL Logical_Operator_out2888_out1            : std_logic;
  SIGNAL Logical_Operator_out2889_out1            : std_logic;
  SIGNAL Logical_Operator_out2890_out1            : std_logic;
  SIGNAL Logical_Operator_out2891_out1            : std_logic;
  SIGNAL Logical_Operator_out2892_out1            : std_logic;
  SIGNAL Logical_Operator_out2893_out1            : std_logic;
  SIGNAL Logical_Operator_out2894_out1            : std_logic;
  SIGNAL Logical_Operator_out2895_out1            : std_logic;
  SIGNAL Logical_Operator_out2896_out1            : std_logic;
  SIGNAL Logical_Operator_out2897_out1            : std_logic;
  SIGNAL Logical_Operator_out2898_out1            : std_logic;
  SIGNAL Logical_Operator_out2899_out1            : std_logic;
  SIGNAL Logical_Operator_out2900_out1            : std_logic;
  SIGNAL Logical_Operator_out2901_out1            : std_logic;
  SIGNAL Logical_Operator_out2902_out1            : std_logic;
  SIGNAL Logical_Operator_out2903_out1            : std_logic;
  SIGNAL Logical_Operator_out2904_out1            : std_logic;
  SIGNAL Logical_Operator_out2905_out1            : std_logic;
  SIGNAL Logical_Operator_out2906_out1            : std_logic;
  SIGNAL Logical_Operator_out2907_out1            : std_logic;
  SIGNAL Logical_Operator_out2908_out1            : std_logic;
  SIGNAL Logical_Operator_out2909_out1            : std_logic;
  SIGNAL Logical_Operator_out2910_out1            : std_logic;
  SIGNAL Logical_Operator_out2911_out1            : std_logic;
  SIGNAL Logical_Operator_out2912_out1            : std_logic;
  SIGNAL Logical_Operator_out2913_out1            : std_logic;
  SIGNAL Logical_Operator_out2914_out1            : std_logic;
  SIGNAL Logical_Operator_out2915_out1            : std_logic;
  SIGNAL Logical_Operator_out2916_out1            : std_logic;
  SIGNAL Logical_Operator_out2917_out1            : std_logic;
  SIGNAL Logical_Operator_out2918_out1            : std_logic;
  SIGNAL Logical_Operator_out2919_out1            : std_logic;
  SIGNAL Logical_Operator_out2920_out1            : std_logic;
  SIGNAL Logical_Operator_out2921_out1            : std_logic;
  SIGNAL Logical_Operator_out2922_out1            : std_logic;
  SIGNAL Logical_Operator_out2923_out1            : std_logic;
  SIGNAL Logical_Operator_out2924_out1            : std_logic;
  SIGNAL Logical_Operator_out2925_out1            : std_logic;
  SIGNAL Logical_Operator_out2926_out1            : std_logic;
  SIGNAL Logical_Operator_out2927_out1            : std_logic;
  SIGNAL Logical_Operator_out2928_out1            : std_logic;
  SIGNAL Logical_Operator_out2929_out1            : std_logic;
  SIGNAL Logical_Operator_out2930_out1            : std_logic;
  SIGNAL Logical_Operator_out2931_out1            : std_logic;
  SIGNAL Logical_Operator_out2932_out1            : std_logic;
  SIGNAL Logical_Operator_out2933_out1            : std_logic;
  SIGNAL Logical_Operator_out2934_out1            : std_logic;
  SIGNAL Logical_Operator_out2935_out1            : std_logic;
  SIGNAL Logical_Operator_out2936_out1            : std_logic;
  SIGNAL Logical_Operator_out2937_out1            : std_logic;
  SIGNAL Logical_Operator_out2938_out1            : std_logic;
  SIGNAL Logical_Operator_out2939_out1            : std_logic;
  SIGNAL Logical_Operator_out2940_out1            : std_logic;
  SIGNAL Logical_Operator_out2941_out1            : std_logic;
  SIGNAL Logical_Operator_out2942_out1            : std_logic;
  SIGNAL Logical_Operator_out2943_out1            : std_logic;
  SIGNAL Logical_Operator_out2944_out1            : std_logic;
  SIGNAL Logical_Operator_out2945_out1            : std_logic;
  SIGNAL Logical_Operator_out2946_out1            : std_logic;
  SIGNAL Logical_Operator_out2947_out1            : std_logic;
  SIGNAL Logical_Operator_out2948_out1            : std_logic;
  SIGNAL Logical_Operator_out2949_out1            : std_logic;
  SIGNAL Logical_Operator_out2950_out1            : std_logic;
  SIGNAL Logical_Operator_out2951_out1            : std_logic;
  SIGNAL Logical_Operator_out2952_out1            : std_logic;
  SIGNAL Logical_Operator_out2953_out1            : std_logic;
  SIGNAL Logical_Operator_out2954_out1            : std_logic;
  SIGNAL Logical_Operator_out2955_out1            : std_logic;
  SIGNAL Logical_Operator_out2956_out1            : std_logic;
  SIGNAL Logical_Operator_out2957_out1            : std_logic;
  SIGNAL Logical_Operator_out2958_out1            : std_logic;
  SIGNAL Logical_Operator_out2959_out1            : std_logic;
  SIGNAL Logical_Operator_out2960_out1            : std_logic;
  SIGNAL Logical_Operator_out2961_out1            : std_logic;
  SIGNAL Logical_Operator_out2962_out1            : std_logic;
  SIGNAL Logical_Operator_out2963_out1            : std_logic;
  SIGNAL Logical_Operator_out2964_out1            : std_logic;
  SIGNAL Logical_Operator_out2965_out1            : std_logic;
  SIGNAL Logical_Operator_out2966_out1            : std_logic;
  SIGNAL Logical_Operator_out2967_out1            : std_logic;
  SIGNAL Logical_Operator_out2968_out1            : std_logic;
  SIGNAL Logical_Operator_out2969_out1            : std_logic;
  SIGNAL Logical_Operator_out2970_out1            : std_logic;
  SIGNAL Logical_Operator_out2971_out1            : std_logic;
  SIGNAL Logical_Operator_out2972_out1            : std_logic;
  SIGNAL Logical_Operator_out2973_out1            : std_logic;
  SIGNAL Logical_Operator_out2974_out1            : std_logic;
  SIGNAL Logical_Operator_out2975_out1            : std_logic;
  SIGNAL Logical_Operator_out2976_out1            : std_logic;
  SIGNAL Logical_Operator_out2977_out1            : std_logic;
  SIGNAL Logical_Operator_out2978_out1            : std_logic;
  SIGNAL Logical_Operator_out2979_out1            : std_logic;
  SIGNAL Logical_Operator_out2980_out1            : std_logic;
  SIGNAL Logical_Operator_out2981_out1            : std_logic;
  SIGNAL Logical_Operator_out2982_out1            : std_logic;
  SIGNAL Logical_Operator_out2983_out1            : std_logic;
  SIGNAL Logical_Operator_out2984_out1            : std_logic;
  SIGNAL Logical_Operator_out2985_out1            : std_logic;
  SIGNAL Logical_Operator_out2986_out1            : std_logic;
  SIGNAL Logical_Operator_out2987_out1            : std_logic;
  SIGNAL Logical_Operator_out2988_out1            : std_logic;
  SIGNAL Logical_Operator_out2989_out1            : std_logic;
  SIGNAL Logical_Operator_out2990_out1            : std_logic;
  SIGNAL Logical_Operator_out2991_out1            : std_logic;
  SIGNAL Logical_Operator_out2992_out1            : std_logic;
  SIGNAL Logical_Operator_out2993_out1            : std_logic;
  SIGNAL Logical_Operator_out2994_out1            : std_logic;
  SIGNAL Logical_Operator_out2995_out1            : std_logic;
  SIGNAL Logical_Operator_out2996_out1            : std_logic;
  SIGNAL Logical_Operator_out2997_out1            : std_logic;
  SIGNAL Logical_Operator_out2998_out1            : std_logic;
  SIGNAL Logical_Operator_out2999_out1            : std_logic;
  SIGNAL Logical_Operator_out3000_out1            : std_logic;
  SIGNAL Logical_Operator_out3001_out1            : std_logic;
  SIGNAL Logical_Operator_out3002_out1            : std_logic;
  SIGNAL Logical_Operator_out3003_out1            : std_logic;
  SIGNAL Logical_Operator_out3004_out1            : std_logic;
  SIGNAL Logical_Operator_out3005_out1            : std_logic;
  SIGNAL Logical_Operator_out3006_out1            : std_logic;
  SIGNAL Logical_Operator_out3007_out1            : std_logic;
  SIGNAL Logical_Operator_out3008_out1            : std_logic;
  SIGNAL Logical_Operator_out3009_out1            : std_logic;
  SIGNAL Logical_Operator_out3010_out1            : std_logic;
  SIGNAL Logical_Operator_out3011_out1            : std_logic;
  SIGNAL Logical_Operator_out3012_out1            : std_logic;
  SIGNAL Logical_Operator_out3013_out1            : std_logic;
  SIGNAL Logical_Operator_out3014_out1            : std_logic;
  SIGNAL Logical_Operator_out3015_out1            : std_logic;
  SIGNAL Logical_Operator_out3016_out1            : std_logic;
  SIGNAL Logical_Operator_out3017_out1            : std_logic;
  SIGNAL Logical_Operator_out3018_out1            : std_logic;
  SIGNAL Logical_Operator_out3019_out1            : std_logic;
  SIGNAL Logical_Operator_out3020_out1            : std_logic;
  SIGNAL Logical_Operator_out3021_out1            : std_logic;
  SIGNAL Logical_Operator_out3022_out1            : std_logic;
  SIGNAL Logical_Operator_out3023_out1            : std_logic;
  SIGNAL Logical_Operator_out3024_out1            : std_logic;
  SIGNAL Logical_Operator_out3025_out1            : std_logic;
  SIGNAL Logical_Operator_out3026_out1            : std_logic;
  SIGNAL Logical_Operator_out3027_out1            : std_logic;
  SIGNAL Logical_Operator_out3028_out1            : std_logic;
  SIGNAL Logical_Operator_out3029_out1            : std_logic;
  SIGNAL Logical_Operator_out3030_out1            : std_logic;
  SIGNAL Logical_Operator_out3031_out1            : std_logic;
  SIGNAL Logical_Operator_out3032_out1            : std_logic;
  SIGNAL Logical_Operator_out3033_out1            : std_logic;
  SIGNAL Logical_Operator_out3034_out1            : std_logic;
  SIGNAL Logical_Operator_out3035_out1            : std_logic;
  SIGNAL Logical_Operator_out3036_out1            : std_logic;
  SIGNAL Logical_Operator_out3037_out1            : std_logic;
  SIGNAL Logical_Operator_out3038_out1            : std_logic;
  SIGNAL Logical_Operator_out3039_out1            : std_logic;
  SIGNAL Logical_Operator_out3040_out1            : std_logic;
  SIGNAL Logical_Operator_out3041_out1            : std_logic;
  SIGNAL Logical_Operator_out3042_out1            : std_logic;
  SIGNAL Logical_Operator_out3043_out1            : std_logic;
  SIGNAL Logical_Operator_out3044_out1            : std_logic;
  SIGNAL Logical_Operator_out3045_out1            : std_logic;
  SIGNAL Logical_Operator_out3046_out1            : std_logic;
  SIGNAL Logical_Operator_out3047_out1            : std_logic;
  SIGNAL Logical_Operator_out3048_out1            : std_logic;
  SIGNAL Logical_Operator_out3049_out1            : std_logic;
  SIGNAL Logical_Operator_out3050_out1            : std_logic;
  SIGNAL Logical_Operator_out3051_out1            : std_logic;
  SIGNAL Logical_Operator_out3052_out1            : std_logic;
  SIGNAL Logical_Operator_out3053_out1            : std_logic;
  SIGNAL Logical_Operator_out3054_out1            : std_logic;
  SIGNAL Logical_Operator_out3055_out1            : std_logic;
  SIGNAL Logical_Operator_out3056_out1            : std_logic;
  SIGNAL Logical_Operator_out3057_out1            : std_logic;
  SIGNAL Logical_Operator_out3058_out1            : std_logic;
  SIGNAL Logical_Operator_out3059_out1            : std_logic;
  SIGNAL Logical_Operator_out3060_out1            : std_logic;
  SIGNAL Logical_Operator_out3061_out1            : std_logic;
  SIGNAL Logical_Operator_out3062_out1            : std_logic;
  SIGNAL Logical_Operator_out3063_out1            : std_logic;
  SIGNAL Logical_Operator_out3064_out1            : std_logic;
  SIGNAL Logical_Operator_out3065_out1            : std_logic;
  SIGNAL Logical_Operator_out3066_out1            : std_logic;
  SIGNAL Logical_Operator_out3067_out1            : std_logic;
  SIGNAL Logical_Operator_out3068_out1            : std_logic;
  SIGNAL Logical_Operator_out3069_out1            : std_logic;
  SIGNAL Logical_Operator_out3070_out1            : std_logic;
  SIGNAL Logical_Operator_out3071_out1            : std_logic;
  SIGNAL Logical_Operator_out3072_out1            : std_logic;
  SIGNAL Logical_Operator_out3073_out1            : std_logic;
  SIGNAL Logical_Operator_out3074_out1            : std_logic;
  SIGNAL Logical_Operator_out3075_out1            : std_logic;
  SIGNAL Logical_Operator_out3076_out1            : std_logic;
  SIGNAL Logical_Operator_out3077_out1            : std_logic;
  SIGNAL Logical_Operator_out3078_out1            : std_logic;
  SIGNAL Logical_Operator_out3079_out1            : std_logic;
  SIGNAL Logical_Operator_out3080_out1            : std_logic;
  SIGNAL Logical_Operator_out3081_out1            : std_logic;
  SIGNAL Logical_Operator_out3082_out1            : std_logic;
  SIGNAL Logical_Operator_out3083_out1            : std_logic;
  SIGNAL Logical_Operator_out3084_out1            : std_logic;
  SIGNAL Logical_Operator_out3085_out1            : std_logic;
  SIGNAL Logical_Operator_out3086_out1            : std_logic;
  SIGNAL Logical_Operator_out3087_out1            : std_logic;
  SIGNAL Logical_Operator_out3088_out1            : std_logic;
  SIGNAL Logical_Operator_out3089_out1            : std_logic;
  SIGNAL Logical_Operator_out3090_out1            : std_logic;
  SIGNAL Logical_Operator_out3091_out1            : std_logic;
  SIGNAL Logical_Operator_out3092_out1            : std_logic;
  SIGNAL Logical_Operator_out3093_out1            : std_logic;
  SIGNAL Logical_Operator_out3094_out1            : std_logic;
  SIGNAL Logical_Operator_out3095_out1            : std_logic;
  SIGNAL Logical_Operator_out3096_out1            : std_logic;
  SIGNAL Logical_Operator_out3097_out1            : std_logic;
  SIGNAL Logical_Operator_out3098_out1            : std_logic;
  SIGNAL Logical_Operator_out3099_out1            : std_logic;
  SIGNAL Logical_Operator_out3100_out1            : std_logic;
  SIGNAL Logical_Operator_out3101_out1            : std_logic;
  SIGNAL Logical_Operator_out3102_out1            : std_logic;
  SIGNAL Logical_Operator_out3103_out1            : std_logic;
  SIGNAL Logical_Operator_out3104_out1            : std_logic;
  SIGNAL Logical_Operator_out3105_out1            : std_logic;
  SIGNAL Logical_Operator_out3106_out1            : std_logic;
  SIGNAL Logical_Operator_out3107_out1            : std_logic;
  SIGNAL Logical_Operator_out3108_out1            : std_logic;
  SIGNAL Logical_Operator_out3109_out1            : std_logic;
  SIGNAL Logical_Operator_out3110_out1            : std_logic;
  SIGNAL Logical_Operator_out3111_out1            : std_logic;
  SIGNAL Logical_Operator_out3112_out1            : std_logic;
  SIGNAL Logical_Operator_out3113_out1            : std_logic;
  SIGNAL Logical_Operator_out3114_out1            : std_logic;
  SIGNAL Logical_Operator_out3115_out1            : std_logic;
  SIGNAL Logical_Operator_out3116_out1            : std_logic;
  SIGNAL Logical_Operator_out3117_out1            : std_logic;
  SIGNAL Logical_Operator_out3118_out1            : std_logic;
  SIGNAL Logical_Operator_out3119_out1            : std_logic;
  SIGNAL Logical_Operator_out3120_out1            : std_logic;
  SIGNAL Logical_Operator_out3121_out1            : std_logic;
  SIGNAL Logical_Operator_out3122_out1            : std_logic;
  SIGNAL Logical_Operator_out3123_out1            : std_logic;
  SIGNAL Logical_Operator_out3124_out1            : std_logic;
  SIGNAL Logical_Operator_out3125_out1            : std_logic;
  SIGNAL Logical_Operator_out3126_out1            : std_logic;
  SIGNAL Logical_Operator_out3127_out1            : std_logic;
  SIGNAL Logical_Operator_out3128_out1            : std_logic;
  SIGNAL Logical_Operator_out3129_out1            : std_logic;
  SIGNAL Logical_Operator_out3130_out1            : std_logic;
  SIGNAL Logical_Operator_out3131_out1            : std_logic;
  SIGNAL Logical_Operator_out3132_out1            : std_logic;
  SIGNAL Logical_Operator_out3133_out1            : std_logic;
  SIGNAL Logical_Operator_out3134_out1            : std_logic;
  SIGNAL Logical_Operator_out3135_out1            : std_logic;
  SIGNAL Logical_Operator_out3136_out1            : std_logic;
  SIGNAL Logical_Operator_out3137_out1            : std_logic;
  SIGNAL Logical_Operator_out3138_out1            : std_logic;
  SIGNAL Logical_Operator_out3139_out1            : std_logic;
  SIGNAL Logical_Operator_out3140_out1            : std_logic;
  SIGNAL Logical_Operator_out3141_out1            : std_logic;
  SIGNAL Logical_Operator_out3142_out1            : std_logic;
  SIGNAL Logical_Operator_out3143_out1            : std_logic;
  SIGNAL Logical_Operator_out3144_out1            : std_logic;
  SIGNAL Logical_Operator_out3145_out1            : std_logic;
  SIGNAL Logical_Operator_out3146_out1            : std_logic;
  SIGNAL Logical_Operator_out3147_out1            : std_logic;
  SIGNAL Logical_Operator_out3148_out1            : std_logic;
  SIGNAL Logical_Operator_out3149_out1            : std_logic;
  SIGNAL Logical_Operator_out3150_out1            : std_logic;
  SIGNAL Logical_Operator_out3151_out1            : std_logic;
  SIGNAL Logical_Operator_out3152_out1            : std_logic;
  SIGNAL Logical_Operator_out3153_out1            : std_logic;
  SIGNAL Logical_Operator_out3154_out1            : std_logic;
  SIGNAL Logical_Operator_out3155_out1            : std_logic;
  SIGNAL Logical_Operator_out3156_out1            : std_logic;
  SIGNAL Logical_Operator_out3157_out1            : std_logic;
  SIGNAL Logical_Operator_out3158_out1            : std_logic;
  SIGNAL Logical_Operator_out3159_out1            : std_logic;
  SIGNAL Logical_Operator_out3160_out1            : std_logic;
  SIGNAL Logical_Operator_out3161_out1            : std_logic;
  SIGNAL Logical_Operator_out3162_out1            : std_logic;
  SIGNAL Logical_Operator_out3163_out1            : std_logic;
  SIGNAL Logical_Operator_out3164_out1            : std_logic;
  SIGNAL Logical_Operator_out3165_out1            : std_logic;
  SIGNAL Logical_Operator_out3166_out1            : std_logic;
  SIGNAL Logical_Operator_out3167_out1            : std_logic;
  SIGNAL Logical_Operator_out3168_out1            : std_logic;
  SIGNAL Logical_Operator_out3169_out1            : std_logic;
  SIGNAL Logical_Operator_out3170_out1            : std_logic;
  SIGNAL Logical_Operator_out3171_out1            : std_logic;
  SIGNAL Logical_Operator_out3172_out1            : std_logic;
  SIGNAL Logical_Operator_out3173_out1            : std_logic;
  SIGNAL Logical_Operator_out3174_out1            : std_logic;
  SIGNAL Logical_Operator_out3175_out1            : std_logic;
  SIGNAL Logical_Operator_out3176_out1            : std_logic;
  SIGNAL Logical_Operator_out3177_out1            : std_logic;
  SIGNAL Logical_Operator_out3178_out1            : std_logic;
  SIGNAL Logical_Operator_out3179_out1            : std_logic;
  SIGNAL Logical_Operator_out3180_out1            : std_logic;
  SIGNAL Logical_Operator_out3181_out1            : std_logic;
  SIGNAL Logical_Operator_out3182_out1            : std_logic;
  SIGNAL Logical_Operator_out3183_out1            : std_logic;
  SIGNAL Logical_Operator_out3184_out1            : std_logic;
  SIGNAL Logical_Operator_out3185_out1            : std_logic;
  SIGNAL Logical_Operator_out3186_out1            : std_logic;
  SIGNAL Logical_Operator_out3187_out1            : std_logic;
  SIGNAL Logical_Operator_out3188_out1            : std_logic;
  SIGNAL Logical_Operator_out3189_out1            : std_logic;
  SIGNAL Logical_Operator_out3190_out1            : std_logic;
  SIGNAL Logical_Operator_out3191_out1            : std_logic;
  SIGNAL Logical_Operator_out3192_out1            : std_logic;
  SIGNAL Logical_Operator_out3193_out1            : std_logic;
  SIGNAL Logical_Operator_out3194_out1            : std_logic;
  SIGNAL Logical_Operator_out3195_out1            : std_logic;
  SIGNAL Logical_Operator_out3196_out1            : std_logic;
  SIGNAL Logical_Operator_out3197_out1            : std_logic;
  SIGNAL Logical_Operator_out3198_out1            : std_logic;
  SIGNAL Logical_Operator_out3199_out1            : std_logic;
  SIGNAL Logical_Operator_out3200_out1            : std_logic;
  SIGNAL Logical_Operator_out3201_out1            : std_logic;
  SIGNAL Logical_Operator_out3202_out1            : std_logic;
  SIGNAL Logical_Operator_out3203_out1            : std_logic;
  SIGNAL Logical_Operator_out3204_out1            : std_logic;
  SIGNAL Logical_Operator_out3205_out1            : std_logic;
  SIGNAL Logical_Operator_out3206_out1            : std_logic;
  SIGNAL Logical_Operator_out3207_out1            : std_logic;
  SIGNAL Logical_Operator_out3208_out1            : std_logic;
  SIGNAL Logical_Operator_out3209_out1            : std_logic;
  SIGNAL Logical_Operator_out3210_out1            : std_logic;
  SIGNAL Logical_Operator_out3211_out1            : std_logic;
  SIGNAL Logical_Operator_out3212_out1            : std_logic;
  SIGNAL Logical_Operator_out3213_out1            : std_logic;
  SIGNAL Logical_Operator_out3214_out1            : std_logic;
  SIGNAL Logical_Operator_out3215_out1            : std_logic;
  SIGNAL Logical_Operator_out3216_out1            : std_logic;
  SIGNAL Logical_Operator_out3217_out1            : std_logic;
  SIGNAL Logical_Operator_out3218_out1            : std_logic;
  SIGNAL Logical_Operator_out3219_out1            : std_logic;
  SIGNAL Logical_Operator_out3220_out1            : std_logic;
  SIGNAL Logical_Operator_out3221_out1            : std_logic;
  SIGNAL Logical_Operator_out3222_out1            : std_logic;
  SIGNAL Logical_Operator_out3223_out1            : std_logic;
  SIGNAL Logical_Operator_out3224_out1            : std_logic;
  SIGNAL Logical_Operator_out3225_out1            : std_logic;
  SIGNAL Logical_Operator_out3226_out1            : std_logic;
  SIGNAL Logical_Operator_out3227_out1            : std_logic;
  SIGNAL Logical_Operator_out3228_out1            : std_logic;
  SIGNAL Logical_Operator_out3229_out1            : std_logic;
  SIGNAL Logical_Operator_out3230_out1            : std_logic;
  SIGNAL Logical_Operator_out3231_out1            : std_logic;
  SIGNAL Logical_Operator_out3232_out1            : std_logic;
  SIGNAL Logical_Operator_out3233_out1            : std_logic;
  SIGNAL Logical_Operator_out3234_out1            : std_logic;
  SIGNAL Logical_Operator_out3235_out1            : std_logic;
  SIGNAL Logical_Operator_out3236_out1            : std_logic;
  SIGNAL Logical_Operator_out3237_out1            : std_logic;
  SIGNAL Logical_Operator_out3238_out1            : std_logic;
  SIGNAL Logical_Operator_out3239_out1            : std_logic;
  SIGNAL Logical_Operator_out3240_out1            : std_logic;
  SIGNAL Logical_Operator_out3241_out1            : std_logic;
  SIGNAL Logical_Operator_out3242_out1            : std_logic;
  SIGNAL Logical_Operator_out3243_out1            : std_logic;
  SIGNAL Logical_Operator_out3244_out1            : std_logic;
  SIGNAL Logical_Operator_out3245_out1            : std_logic;
  SIGNAL Logical_Operator_out3246_out1            : std_logic;
  SIGNAL Logical_Operator_out3247_out1            : std_logic;
  SIGNAL Logical_Operator_out3248_out1            : std_logic;
  SIGNAL Logical_Operator_out3249_out1            : std_logic;
  SIGNAL Logical_Operator_out3250_out1            : std_logic;
  SIGNAL Logical_Operator_out3251_out1            : std_logic;
  SIGNAL Logical_Operator_out3252_out1            : std_logic;
  SIGNAL Logical_Operator_out3253_out1            : std_logic;
  SIGNAL Logical_Operator_out3254_out1            : std_logic;
  SIGNAL Logical_Operator_out3255_out1            : std_logic;
  SIGNAL Logical_Operator_out3256_out1            : std_logic;
  SIGNAL Logical_Operator_out3257_out1            : std_logic;
  SIGNAL Logical_Operator_out3258_out1            : std_logic;
  SIGNAL Logical_Operator_out3259_out1            : std_logic;
  SIGNAL Logical_Operator_out3260_out1            : std_logic;
  SIGNAL Logical_Operator_out3261_out1            : std_logic;
  SIGNAL Logical_Operator_out3262_out1            : std_logic;
  SIGNAL Logical_Operator_out3263_out1            : std_logic;
  SIGNAL Logical_Operator_out3264_out1            : std_logic;
  SIGNAL Logical_Operator_out3265_out1            : std_logic;
  SIGNAL Logical_Operator_out3266_out1            : std_logic;
  SIGNAL Logical_Operator_out3267_out1            : std_logic;
  SIGNAL Logical_Operator_out3268_out1            : std_logic;
  SIGNAL Logical_Operator_out3269_out1            : std_logic;
  SIGNAL Logical_Operator_out3270_out1            : std_logic;
  SIGNAL Logical_Operator_out3271_out1            : std_logic;
  SIGNAL Logical_Operator_out3272_out1            : std_logic;
  SIGNAL Logical_Operator_out3273_out1            : std_logic;
  SIGNAL Logical_Operator_out3274_out1            : std_logic;
  SIGNAL Logical_Operator_out3275_out1            : std_logic;
  SIGNAL Logical_Operator_out3276_out1            : std_logic;
  SIGNAL Logical_Operator_out3277_out1            : std_logic;
  SIGNAL Logical_Operator_out3278_out1            : std_logic;
  SIGNAL Logical_Operator_out3279_out1            : std_logic;
  SIGNAL Logical_Operator_out3280_out1            : std_logic;
  SIGNAL Logical_Operator_out3281_out1            : std_logic;
  SIGNAL Logical_Operator_out3282_out1            : std_logic;
  SIGNAL Logical_Operator_out3283_out1            : std_logic;
  SIGNAL Logical_Operator_out3284_out1            : std_logic;
  SIGNAL Logical_Operator_out3285_out1            : std_logic;
  SIGNAL Logical_Operator_out3286_out1            : std_logic;
  SIGNAL Logical_Operator_out3287_out1            : std_logic;
  SIGNAL Logical_Operator_out3288_out1            : std_logic;
  SIGNAL Logical_Operator_out3289_out1            : std_logic;
  SIGNAL Logical_Operator_out3290_out1            : std_logic;
  SIGNAL Logical_Operator_out3291_out1            : std_logic;
  SIGNAL Logical_Operator_out3292_out1            : std_logic;
  SIGNAL Logical_Operator_out3293_out1            : std_logic;
  SIGNAL Logical_Operator_out3294_out1            : std_logic;
  SIGNAL Logical_Operator_out3295_out1            : std_logic;
  SIGNAL Logical_Operator_out3296_out1            : std_logic;
  SIGNAL Logical_Operator_out3297_out1            : std_logic;
  SIGNAL Logical_Operator_out3298_out1            : std_logic;
  SIGNAL Logical_Operator_out3299_out1            : std_logic;
  SIGNAL Logical_Operator_out3300_out1            : std_logic;
  SIGNAL Logical_Operator_out3301_out1            : std_logic;
  SIGNAL Logical_Operator_out3302_out1            : std_logic;
  SIGNAL Logical_Operator_out3303_out1            : std_logic;
  SIGNAL Logical_Operator_out3304_out1            : std_logic;
  SIGNAL Logical_Operator_out3305_out1            : std_logic;
  SIGNAL Logical_Operator_out3306_out1            : std_logic;
  SIGNAL Logical_Operator_out3307_out1            : std_logic;
  SIGNAL Logical_Operator_out3308_out1            : std_logic;
  SIGNAL Logical_Operator_out3309_out1            : std_logic;
  SIGNAL Logical_Operator_out3310_out1            : std_logic;
  SIGNAL Logical_Operator_out3311_out1            : std_logic;
  SIGNAL Logical_Operator_out3312_out1            : std_logic;
  SIGNAL Logical_Operator_out3313_out1            : std_logic;
  SIGNAL Logical_Operator_out3314_out1            : std_logic;
  SIGNAL Logical_Operator_out3315_out1            : std_logic;
  SIGNAL Logical_Operator_out3316_out1            : std_logic;
  SIGNAL Logical_Operator_out3317_out1            : std_logic;
  SIGNAL Logical_Operator_out3318_out1            : std_logic;
  SIGNAL Logical_Operator_out3319_out1            : std_logic;
  SIGNAL Logical_Operator_out3320_out1            : std_logic;
  SIGNAL Logical_Operator_out3321_out1            : std_logic;
  SIGNAL Logical_Operator_out3322_out1            : std_logic;
  SIGNAL Logical_Operator_out3323_out1            : std_logic;
  SIGNAL Logical_Operator_out3324_out1            : std_logic;
  SIGNAL Logical_Operator_out3325_out1            : std_logic;
  SIGNAL Logical_Operator_out3326_out1            : std_logic;
  SIGNAL Logical_Operator_out3327_out1            : std_logic;
  SIGNAL Logical_Operator_out3328_out1            : std_logic;
  SIGNAL Logical_Operator_out3329_out1            : std_logic;
  SIGNAL Logical_Operator_out3330_out1            : std_logic;
  SIGNAL Logical_Operator_out3331_out1            : std_logic;
  SIGNAL Logical_Operator_out3332_out1            : std_logic;
  SIGNAL Logical_Operator_out3333_out1            : std_logic;
  SIGNAL Logical_Operator_out3334_out1            : std_logic;
  SIGNAL Logical_Operator_out3335_out1            : std_logic;
  SIGNAL Logical_Operator_out3336_out1            : std_logic;
  SIGNAL Logical_Operator_out3337_out1            : std_logic;
  SIGNAL Logical_Operator_out3338_out1            : std_logic;
  SIGNAL Logical_Operator_out3339_out1            : std_logic;
  SIGNAL Logical_Operator_out3340_out1            : std_logic;
  SIGNAL Logical_Operator_out3341_out1            : std_logic;
  SIGNAL Logical_Operator_out3342_out1            : std_logic;
  SIGNAL Logical_Operator_out3343_out1            : std_logic;
  SIGNAL Logical_Operator_out3344_out1            : std_logic;
  SIGNAL Logical_Operator_out3345_out1            : std_logic;
  SIGNAL Logical_Operator_out3346_out1            : std_logic;
  SIGNAL Logical_Operator_out3347_out1            : std_logic;
  SIGNAL Logical_Operator_out3348_out1            : std_logic;
  SIGNAL Logical_Operator_out3349_out1            : std_logic;
  SIGNAL Logical_Operator_out3350_out1            : std_logic;
  SIGNAL Logical_Operator_out3351_out1            : std_logic;
  SIGNAL Logical_Operator_out3352_out1            : std_logic;
  SIGNAL Logical_Operator_out3353_out1            : std_logic;
  SIGNAL Logical_Operator_out3354_out1            : std_logic;
  SIGNAL Logical_Operator_out3355_out1            : std_logic;
  SIGNAL Logical_Operator_out3356_out1            : std_logic;
  SIGNAL Logical_Operator_out3357_out1            : std_logic;
  SIGNAL Logical_Operator_out3358_out1            : std_logic;
  SIGNAL Logical_Operator_out3359_out1            : std_logic;
  SIGNAL Logical_Operator_out3360_out1            : std_logic;
  SIGNAL Logical_Operator_out3361_out1            : std_logic;
  SIGNAL Logical_Operator_out3362_out1            : std_logic;
  SIGNAL Logical_Operator_out3363_out1            : std_logic;
  SIGNAL Logical_Operator_out3364_out1            : std_logic;
  SIGNAL Logical_Operator_out3365_out1            : std_logic;
  SIGNAL Logical_Operator_out3366_out1            : std_logic;
  SIGNAL Logical_Operator_out3367_out1            : std_logic;
  SIGNAL Logical_Operator_out3368_out1            : std_logic;
  SIGNAL Logical_Operator_out3369_out1            : std_logic;
  SIGNAL Logical_Operator_out3370_out1            : std_logic;
  SIGNAL Logical_Operator_out3371_out1            : std_logic;
  SIGNAL Logical_Operator_out3372_out1            : std_logic;
  SIGNAL Logical_Operator_out3373_out1            : std_logic;
  SIGNAL Logical_Operator_out3374_out1            : std_logic;
  SIGNAL Logical_Operator_out3375_out1            : std_logic;
  SIGNAL Logical_Operator_out3376_out1            : std_logic;
  SIGNAL Logical_Operator_out3377_out1            : std_logic;
  SIGNAL Logical_Operator_out3378_out1            : std_logic;
  SIGNAL Logical_Operator_out3379_out1            : std_logic;
  SIGNAL Logical_Operator_out3380_out1            : std_logic;
  SIGNAL Logical_Operator_out3381_out1            : std_logic;
  SIGNAL Logical_Operator_out3382_out1            : std_logic;
  SIGNAL Logical_Operator_out3383_out1            : std_logic;
  SIGNAL Logical_Operator_out3384_out1            : std_logic;
  SIGNAL Logical_Operator_out3385_out1            : std_logic;
  SIGNAL Logical_Operator_out3386_out1            : std_logic;
  SIGNAL Logical_Operator_out3387_out1            : std_logic;
  SIGNAL Logical_Operator_out3388_out1            : std_logic;
  SIGNAL Logical_Operator_out3389_out1            : std_logic;
  SIGNAL Logical_Operator_out3390_out1            : std_logic;
  SIGNAL Logical_Operator_out3391_out1            : std_logic;
  SIGNAL Logical_Operator_out3392_out1            : std_logic;
  SIGNAL Logical_Operator_out3393_out1            : std_logic;
  SIGNAL Logical_Operator_out3394_out1            : std_logic;
  SIGNAL Logical_Operator_out3395_out1            : std_logic;
  SIGNAL Logical_Operator_out3396_out1            : std_logic;
  SIGNAL Logical_Operator_out3397_out1            : std_logic;
  SIGNAL Logical_Operator_out3398_out1            : std_logic;
  SIGNAL Logical_Operator_out3399_out1            : std_logic;
  SIGNAL Logical_Operator_out3400_out1            : std_logic;
  SIGNAL Logical_Operator_out3401_out1            : std_logic;
  SIGNAL Logical_Operator_out3402_out1            : std_logic;
  SIGNAL Logical_Operator_out3403_out1            : std_logic;
  SIGNAL Logical_Operator_out3404_out1            : std_logic;
  SIGNAL Logical_Operator_out3405_out1            : std_logic;
  SIGNAL Logical_Operator_out3406_out1            : std_logic;
  SIGNAL Logical_Operator_out3407_out1            : std_logic;
  SIGNAL Logical_Operator_out3408_out1            : std_logic;
  SIGNAL Logical_Operator_out3409_out1            : std_logic;
  SIGNAL Logical_Operator_out3410_out1            : std_logic;
  SIGNAL Logical_Operator_out3411_out1            : std_logic;
  SIGNAL Logical_Operator_out3412_out1            : std_logic;
  SIGNAL Logical_Operator_out3413_out1            : std_logic;
  SIGNAL Logical_Operator_out3414_out1            : std_logic;
  SIGNAL Logical_Operator_out3415_out1            : std_logic;
  SIGNAL Logical_Operator_out3416_out1            : std_logic;
  SIGNAL Logical_Operator_out3417_out1            : std_logic;
  SIGNAL Logical_Operator_out3418_out1            : std_logic;
  SIGNAL Logical_Operator_out3419_out1            : std_logic;
  SIGNAL Logical_Operator_out3420_out1            : std_logic;
  SIGNAL Logical_Operator_out3421_out1            : std_logic;
  SIGNAL Logical_Operator_out3422_out1            : std_logic;
  SIGNAL Logical_Operator_out3423_out1            : std_logic;
  SIGNAL Logical_Operator_out3424_out1            : std_logic;
  SIGNAL Logical_Operator_out3425_out1            : std_logic;
  SIGNAL Logical_Operator_out3426_out1            : std_logic;
  SIGNAL Logical_Operator_out3427_out1            : std_logic;
  SIGNAL Logical_Operator_out3428_out1            : std_logic;
  SIGNAL Logical_Operator_out3429_out1            : std_logic;
  SIGNAL Logical_Operator_out3430_out1            : std_logic;
  SIGNAL Logical_Operator_out3431_out1            : std_logic;
  SIGNAL Logical_Operator_out3432_out1            : std_logic;
  SIGNAL Logical_Operator_out3433_out1            : std_logic;
  SIGNAL Logical_Operator_out3434_out1            : std_logic;
  SIGNAL Logical_Operator_out3435_out1            : std_logic;
  SIGNAL Logical_Operator_out3436_out1            : std_logic;
  SIGNAL Logical_Operator_out3437_out1            : std_logic;
  SIGNAL Logical_Operator_out3438_out1            : std_logic;
  SIGNAL Logical_Operator_out3439_out1            : std_logic;
  SIGNAL Logical_Operator_out3440_out1            : std_logic;
  SIGNAL Logical_Operator_out3441_out1            : std_logic;
  SIGNAL Logical_Operator_out3442_out1            : std_logic;
  SIGNAL Logical_Operator_out3443_out1            : std_logic;
  SIGNAL Logical_Operator_out3444_out1            : std_logic;
  SIGNAL Logical_Operator_out3445_out1            : std_logic;
  SIGNAL Logical_Operator_out3446_out1            : std_logic;
  SIGNAL Logical_Operator_out3447_out1            : std_logic;
  SIGNAL Logical_Operator_out3448_out1            : std_logic;
  SIGNAL Logical_Operator_out3449_out1            : std_logic;
  SIGNAL Logical_Operator_out3450_out1            : std_logic;
  SIGNAL Logical_Operator_out3451_out1            : std_logic;
  SIGNAL Logical_Operator_out3452_out1            : std_logic;
  SIGNAL Logical_Operator_out3453_out1            : std_logic;
  SIGNAL Logical_Operator_out3454_out1            : std_logic;
  SIGNAL Logical_Operator_out3455_out1            : std_logic;
  SIGNAL Logical_Operator_out3456_out1            : std_logic;
  SIGNAL Logical_Operator_out3457_out1            : std_logic;
  SIGNAL Logical_Operator_out3458_out1            : std_logic;
  SIGNAL Logical_Operator_out3459_out1            : std_logic;
  SIGNAL Logical_Operator_out3460_out1            : std_logic;
  SIGNAL Logical_Operator_out3461_out1            : std_logic;
  SIGNAL Logical_Operator_out3462_out1            : std_logic;
  SIGNAL Logical_Operator_out3463_out1            : std_logic;
  SIGNAL Logical_Operator_out3464_out1            : std_logic;
  SIGNAL Logical_Operator_out3465_out1            : std_logic;
  SIGNAL Logical_Operator_out3466_out1            : std_logic;
  SIGNAL Logical_Operator_out3467_out1            : std_logic;
  SIGNAL Logical_Operator_out3468_out1            : std_logic;
  SIGNAL Logical_Operator_out3469_out1            : std_logic;
  SIGNAL Logical_Operator_out3470_out1            : std_logic;
  SIGNAL Logical_Operator_out3471_out1            : std_logic;
  SIGNAL Logical_Operator_out3472_out1            : std_logic;
  SIGNAL Logical_Operator_out3473_out1            : std_logic;
  SIGNAL Logical_Operator_out3474_out1            : std_logic;
  SIGNAL Logical_Operator_out3475_out1            : std_logic;
  SIGNAL Logical_Operator_out3476_out1            : std_logic;
  SIGNAL Logical_Operator_out3477_out1            : std_logic;
  SIGNAL Logical_Operator_out3478_out1            : std_logic;
  SIGNAL Logical_Operator_out3479_out1            : std_logic;
  SIGNAL Logical_Operator_out3480_out1            : std_logic;
  SIGNAL Logical_Operator_out3481_out1            : std_logic;
  SIGNAL Logical_Operator_out3482_out1            : std_logic;
  SIGNAL Logical_Operator_out3483_out1            : std_logic;
  SIGNAL Logical_Operator_out3484_out1            : std_logic;
  SIGNAL Logical_Operator_out3485_out1            : std_logic;
  SIGNAL Logical_Operator_out3486_out1            : std_logic;
  SIGNAL Logical_Operator_out3487_out1            : std_logic;
  SIGNAL Logical_Operator_out3488_out1            : std_logic;
  SIGNAL Logical_Operator_out3489_out1            : std_logic;
  SIGNAL Logical_Operator_out3490_out1            : std_logic;
  SIGNAL Logical_Operator_out3491_out1            : std_logic;
  SIGNAL Logical_Operator_out3492_out1            : std_logic;
  SIGNAL Logical_Operator_out3493_out1            : std_logic;
  SIGNAL Logical_Operator_out3494_out1            : std_logic;
  SIGNAL Logical_Operator_out3495_out1            : std_logic;
  SIGNAL Logical_Operator_out3496_out1            : std_logic;
  SIGNAL Logical_Operator_out3497_out1            : std_logic;
  SIGNAL Logical_Operator_out3498_out1            : std_logic;
  SIGNAL Logical_Operator_out3499_out1            : std_logic;
  SIGNAL Logical_Operator_out3500_out1            : std_logic;
  SIGNAL Logical_Operator_out3501_out1            : std_logic;
  SIGNAL Logical_Operator_out3502_out1            : std_logic;
  SIGNAL Logical_Operator_out3503_out1            : std_logic;
  SIGNAL Logical_Operator_out3504_out1            : std_logic;
  SIGNAL Logical_Operator_out3505_out1            : std_logic;
  SIGNAL Logical_Operator_out3506_out1            : std_logic;
  SIGNAL Logical_Operator_out3507_out1            : std_logic;
  SIGNAL Logical_Operator_out3508_out1            : std_logic;
  SIGNAL Logical_Operator_out3509_out1            : std_logic;
  SIGNAL Logical_Operator_out3510_out1            : std_logic;
  SIGNAL Logical_Operator_out3511_out1            : std_logic;
  SIGNAL Logical_Operator_out3512_out1            : std_logic;
  SIGNAL Logical_Operator_out3513_out1            : std_logic;
  SIGNAL Logical_Operator_out3514_out1            : std_logic;
  SIGNAL Logical_Operator_out3515_out1            : std_logic;
  SIGNAL Logical_Operator_out3516_out1            : std_logic;
  SIGNAL Logical_Operator_out3517_out1            : std_logic;
  SIGNAL Logical_Operator_out3518_out1            : std_logic;
  SIGNAL Logical_Operator_out3519_out1            : std_logic;
  SIGNAL Logical_Operator_out3520_out1            : std_logic;
  SIGNAL Logical_Operator_out3521_out1            : std_logic;
  SIGNAL Logical_Operator_out3522_out1            : std_logic;
  SIGNAL Logical_Operator_out3523_out1            : std_logic;
  SIGNAL Logical_Operator_out3524_out1            : std_logic;
  SIGNAL Logical_Operator_out3525_out1            : std_logic;
  SIGNAL Logical_Operator_out3526_out1            : std_logic;
  SIGNAL Logical_Operator_out3527_out1            : std_logic;
  SIGNAL Logical_Operator_out3528_out1            : std_logic;
  SIGNAL Logical_Operator_out3529_out1            : std_logic;
  SIGNAL Logical_Operator_out3530_out1            : std_logic;
  SIGNAL Logical_Operator_out3531_out1            : std_logic;
  SIGNAL Logical_Operator_out3532_out1            : std_logic;
  SIGNAL Logical_Operator_out3533_out1            : std_logic;
  SIGNAL Logical_Operator_out3534_out1            : std_logic;
  SIGNAL Logical_Operator_out3535_out1            : std_logic;
  SIGNAL Logical_Operator_out3536_out1            : std_logic;
  SIGNAL Logical_Operator_out3537_out1            : std_logic;
  SIGNAL Logical_Operator_out3538_out1            : std_logic;
  SIGNAL Logical_Operator_out3539_out1            : std_logic;
  SIGNAL Logical_Operator_out3540_out1            : std_logic;
  SIGNAL Logical_Operator_out3541_out1            : std_logic;
  SIGNAL Logical_Operator_out3542_out1            : std_logic;
  SIGNAL Logical_Operator_out3543_out1            : std_logic;
  SIGNAL Logical_Operator_out3544_out1            : std_logic;
  SIGNAL Logical_Operator_out3545_out1            : std_logic;
  SIGNAL Logical_Operator_out3546_out1            : std_logic;
  SIGNAL Logical_Operator_out3547_out1            : std_logic;
  SIGNAL Logical_Operator_out3548_out1            : std_logic;
  SIGNAL Logical_Operator_out3549_out1            : std_logic;
  SIGNAL Logical_Operator_out3550_out1            : std_logic;
  SIGNAL Logical_Operator_out3551_out1            : std_logic;
  SIGNAL Logical_Operator_out3552_out1            : std_logic;
  SIGNAL Logical_Operator_out3553_out1            : std_logic;
  SIGNAL Logical_Operator_out3554_out1            : std_logic;
  SIGNAL Logical_Operator_out3555_out1            : std_logic;
  SIGNAL Logical_Operator_out3556_out1            : std_logic;
  SIGNAL Logical_Operator_out3557_out1            : std_logic;
  SIGNAL Logical_Operator_out3558_out1            : std_logic;
  SIGNAL Logical_Operator_out3559_out1            : std_logic;
  SIGNAL Logical_Operator_out3560_out1            : std_logic;
  SIGNAL Logical_Operator_out3561_out1            : std_logic;
  SIGNAL Logical_Operator_out3562_out1            : std_logic;
  SIGNAL Logical_Operator_out3563_out1            : std_logic;
  SIGNAL Logical_Operator_out3564_out1            : std_logic;
  SIGNAL Logical_Operator_out3565_out1            : std_logic;
  SIGNAL Logical_Operator_out3566_out1            : std_logic;
  SIGNAL Logical_Operator_out3567_out1            : std_logic;
  SIGNAL Logical_Operator_out3568_out1            : std_logic;
  SIGNAL Logical_Operator_out3569_out1            : std_logic;
  SIGNAL Logical_Operator_out3570_out1            : std_logic;
  SIGNAL Logical_Operator_out3571_out1            : std_logic;
  SIGNAL Logical_Operator_out3572_out1            : std_logic;
  SIGNAL Logical_Operator_out3573_out1            : std_logic;
  SIGNAL Logical_Operator_out3574_out1            : std_logic;
  SIGNAL Logical_Operator_out3575_out1            : std_logic;
  SIGNAL Logical_Operator_out3576_out1            : std_logic;
  SIGNAL Logical_Operator_out3577_out1            : std_logic;
  SIGNAL Logical_Operator_out3578_out1            : std_logic;
  SIGNAL Logical_Operator_out3579_out1            : std_logic;
  SIGNAL Logical_Operator_out3580_out1            : std_logic;
  SIGNAL Logical_Operator_out3581_out1            : std_logic;
  SIGNAL Logical_Operator_out3582_out1            : std_logic;
  SIGNAL Logical_Operator_out3583_out1            : std_logic;
  SIGNAL Logical_Operator_out3584_out1            : std_logic;
  SIGNAL Logical_Operator_out3585_out1            : std_logic;
  SIGNAL Logical_Operator_out3586_out1            : std_logic;
  SIGNAL Logical_Operator_out3587_out1            : std_logic;
  SIGNAL Logical_Operator_out3588_out1            : std_logic;
  SIGNAL Logical_Operator_out3589_out1            : std_logic;
  SIGNAL Logical_Operator_out3590_out1            : std_logic;
  SIGNAL Logical_Operator_out3591_out1            : std_logic;
  SIGNAL Logical_Operator_out3592_out1            : std_logic;
  SIGNAL Logical_Operator_out3593_out1            : std_logic;
  SIGNAL Logical_Operator_out3594_out1            : std_logic;
  SIGNAL Logical_Operator_out3595_out1            : std_logic;
  SIGNAL Logical_Operator_out3596_out1            : std_logic;
  SIGNAL Logical_Operator_out3597_out1            : std_logic;
  SIGNAL Logical_Operator_out3598_out1            : std_logic;
  SIGNAL Logical_Operator_out3599_out1            : std_logic;
  SIGNAL Logical_Operator_out3600_out1            : std_logic;
  SIGNAL Logical_Operator_out3601_out1            : std_logic;
  SIGNAL Logical_Operator_out3602_out1            : std_logic;
  SIGNAL Logical_Operator_out3603_out1            : std_logic;
  SIGNAL Logical_Operator_out3604_out1            : std_logic;
  SIGNAL Logical_Operator_out3605_out1            : std_logic;
  SIGNAL Logical_Operator_out3606_out1            : std_logic;
  SIGNAL Logical_Operator_out3607_out1            : std_logic;
  SIGNAL Logical_Operator_out3608_out1            : std_logic;
  SIGNAL Logical_Operator_out3609_out1            : std_logic;
  SIGNAL Logical_Operator_out3610_out1            : std_logic;
  SIGNAL Logical_Operator_out3611_out1            : std_logic;
  SIGNAL Logical_Operator_out3612_out1            : std_logic;
  SIGNAL Logical_Operator_out3613_out1            : std_logic;
  SIGNAL Logical_Operator_out3614_out1            : std_logic;
  SIGNAL Logical_Operator_out3615_out1            : std_logic;
  SIGNAL Logical_Operator_out3616_out1            : std_logic;
  SIGNAL Logical_Operator_out3617_out1            : std_logic;
  SIGNAL Logical_Operator_out3618_out1            : std_logic;
  SIGNAL Logical_Operator_out3619_out1            : std_logic;
  SIGNAL Logical_Operator_out3620_out1            : std_logic;
  SIGNAL Logical_Operator_out3621_out1            : std_logic;
  SIGNAL Logical_Operator_out3622_out1            : std_logic;
  SIGNAL Logical_Operator_out3623_out1            : std_logic;
  SIGNAL Logical_Operator_out3624_out1            : std_logic;
  SIGNAL Logical_Operator_out3625_out1            : std_logic;
  SIGNAL Logical_Operator_out3626_out1            : std_logic;
  SIGNAL Logical_Operator_out3627_out1            : std_logic;
  SIGNAL Logical_Operator_out3628_out1            : std_logic;
  SIGNAL Logical_Operator_out3629_out1            : std_logic;
  SIGNAL Logical_Operator_out3630_out1            : std_logic;
  SIGNAL Logical_Operator_out3631_out1            : std_logic;
  SIGNAL Logical_Operator_out3632_out1            : std_logic;
  SIGNAL Logical_Operator_out3633_out1            : std_logic;
  SIGNAL Logical_Operator_out3634_out1            : std_logic;
  SIGNAL Logical_Operator_out3635_out1            : std_logic;
  SIGNAL Logical_Operator_out3636_out1            : std_logic;
  SIGNAL Logical_Operator_out3637_out1            : std_logic;
  SIGNAL Logical_Operator_out3638_out1            : std_logic;
  SIGNAL Logical_Operator_out3639_out1            : std_logic;
  SIGNAL Logical_Operator_out3640_out1            : std_logic;
  SIGNAL Logical_Operator_out3641_out1            : std_logic;
  SIGNAL Logical_Operator_out3642_out1            : std_logic;
  SIGNAL Logical_Operator_out3643_out1            : std_logic;
  SIGNAL Logical_Operator_out3644_out1            : std_logic;
  SIGNAL Logical_Operator_out3645_out1            : std_logic;
  SIGNAL Logical_Operator_out3646_out1            : std_logic;
  SIGNAL Logical_Operator_out3647_out1            : std_logic;
  SIGNAL Logical_Operator_out3648_out1            : std_logic;
  SIGNAL Logical_Operator_out3649_out1            : std_logic;
  SIGNAL Logical_Operator_out3650_out1            : std_logic;
  SIGNAL Logical_Operator_out3651_out1            : std_logic;
  SIGNAL Logical_Operator_out3652_out1            : std_logic;
  SIGNAL Logical_Operator_out3653_out1            : std_logic;
  SIGNAL Logical_Operator_out3654_out1            : std_logic;
  SIGNAL Logical_Operator_out3655_out1            : std_logic;
  SIGNAL Logical_Operator_out3656_out1            : std_logic;
  SIGNAL Logical_Operator_out3657_out1            : std_logic;
  SIGNAL Logical_Operator_out3658_out1            : std_logic;
  SIGNAL Logical_Operator_out3659_out1            : std_logic;
  SIGNAL Logical_Operator_out3660_out1            : std_logic;
  SIGNAL Logical_Operator_out3661_out1            : std_logic;
  SIGNAL Logical_Operator_out3662_out1            : std_logic;
  SIGNAL Logical_Operator_out3663_out1            : std_logic;
  SIGNAL Logical_Operator_out3664_out1            : std_logic;
  SIGNAL Logical_Operator_out3665_out1            : std_logic;
  SIGNAL Logical_Operator_out3666_out1            : std_logic;
  SIGNAL Logical_Operator_out3667_out1            : std_logic;
  SIGNAL Logical_Operator_out3668_out1            : std_logic;
  SIGNAL Logical_Operator_out3669_out1            : std_logic;
  SIGNAL Logical_Operator_out3670_out1            : std_logic;
  SIGNAL Logical_Operator_out3671_out1            : std_logic;
  SIGNAL Logical_Operator_out3672_out1            : std_logic;
  SIGNAL Logical_Operator_out3673_out1            : std_logic;
  SIGNAL Logical_Operator_out3674_out1            : std_logic;
  SIGNAL Logical_Operator_out3675_out1            : std_logic;
  SIGNAL Logical_Operator_out3676_out1            : std_logic;
  SIGNAL Logical_Operator_out3677_out1            : std_logic;
  SIGNAL Logical_Operator_out3678_out1            : std_logic;
  SIGNAL Logical_Operator_out3679_out1            : std_logic;
  SIGNAL Logical_Operator_out3680_out1            : std_logic;
  SIGNAL Logical_Operator_out3681_out1            : std_logic;
  SIGNAL Logical_Operator_out3682_out1            : std_logic;
  SIGNAL Logical_Operator_out3683_out1            : std_logic;
  SIGNAL Logical_Operator_out3684_out1            : std_logic;
  SIGNAL Logical_Operator_out3685_out1            : std_logic;
  SIGNAL Logical_Operator_out3686_out1            : std_logic;
  SIGNAL Logical_Operator_out3687_out1            : std_logic;
  SIGNAL Logical_Operator_out3688_out1            : std_logic;
  SIGNAL Logical_Operator_out3689_out1            : std_logic;
  SIGNAL Logical_Operator_out3690_out1            : std_logic;
  SIGNAL Logical_Operator_out3691_out1            : std_logic;
  SIGNAL Logical_Operator_out3692_out1            : std_logic;
  SIGNAL Logical_Operator_out3693_out1            : std_logic;
  SIGNAL Logical_Operator_out3694_out1            : std_logic;
  SIGNAL Logical_Operator_out3695_out1            : std_logic;
  SIGNAL Logical_Operator_out3696_out1            : std_logic;
  SIGNAL Logical_Operator_out3697_out1            : std_logic;
  SIGNAL Logical_Operator_out3698_out1            : std_logic;
  SIGNAL Logical_Operator_out3699_out1            : std_logic;
  SIGNAL Logical_Operator_out3700_out1            : std_logic;
  SIGNAL Logical_Operator_out3701_out1            : std_logic;
  SIGNAL Logical_Operator_out3702_out1            : std_logic;
  SIGNAL Logical_Operator_out3703_out1            : std_logic;
  SIGNAL Logical_Operator_out3704_out1            : std_logic;
  SIGNAL Logical_Operator_out3705_out1            : std_logic;
  SIGNAL Logical_Operator_out3706_out1            : std_logic;
  SIGNAL Logical_Operator_out3707_out1            : std_logic;
  SIGNAL Logical_Operator_out3708_out1            : std_logic;
  SIGNAL Logical_Operator_out3709_out1            : std_logic;
  SIGNAL Logical_Operator_out3710_out1            : std_logic;
  SIGNAL Logical_Operator_out3711_out1            : std_logic;
  SIGNAL Logical_Operator_out3712_out1            : std_logic;
  SIGNAL Logical_Operator_out3713_out1            : std_logic;
  SIGNAL Logical_Operator_out3714_out1            : std_logic;
  SIGNAL Logical_Operator_out3715_out1            : std_logic;
  SIGNAL Logical_Operator_out3716_out1            : std_logic;
  SIGNAL Logical_Operator_out3717_out1            : std_logic;
  SIGNAL Logical_Operator_out3718_out1            : std_logic;
  SIGNAL Logical_Operator_out3719_out1            : std_logic;
  SIGNAL Logical_Operator_out3720_out1            : std_logic;
  SIGNAL Logical_Operator_out3721_out1            : std_logic;
  SIGNAL Logical_Operator_out3722_out1            : std_logic;
  SIGNAL Logical_Operator_out3723_out1            : std_logic;
  SIGNAL Logical_Operator_out3724_out1            : std_logic;
  SIGNAL Logical_Operator_out3725_out1            : std_logic;
  SIGNAL Logical_Operator_out3726_out1            : std_logic;
  SIGNAL Logical_Operator_out3727_out1            : std_logic;
  SIGNAL Logical_Operator_out3728_out1            : std_logic;
  SIGNAL Logical_Operator_out3729_out1            : std_logic;
  SIGNAL Logical_Operator_out3730_out1            : std_logic;
  SIGNAL Logical_Operator_out3731_out1            : std_logic;
  SIGNAL Logical_Operator_out3732_out1            : std_logic;
  SIGNAL Logical_Operator_out3733_out1            : std_logic;
  SIGNAL Logical_Operator_out3734_out1            : std_logic;
  SIGNAL Logical_Operator_out3735_out1            : std_logic;
  SIGNAL Logical_Operator_out3736_out1            : std_logic;
  SIGNAL Logical_Operator_out3737_out1            : std_logic;
  SIGNAL Logical_Operator_out3738_out1            : std_logic;
  SIGNAL Logical_Operator_out3739_out1            : std_logic;
  SIGNAL Logical_Operator_out3740_out1            : std_logic;
  SIGNAL Logical_Operator_out3741_out1            : std_logic;
  SIGNAL Logical_Operator_out3742_out1            : std_logic;
  SIGNAL Logical_Operator_out3743_out1            : std_logic;
  SIGNAL Logical_Operator_out3744_out1            : std_logic;
  SIGNAL Logical_Operator_out3745_out1            : std_logic;
  SIGNAL Logical_Operator_out3746_out1            : std_logic;
  SIGNAL Logical_Operator_out3747_out1            : std_logic;
  SIGNAL Logical_Operator_out3748_out1            : std_logic;
  SIGNAL Logical_Operator_out3749_out1            : std_logic;
  SIGNAL Logical_Operator_out3750_out1            : std_logic;
  SIGNAL Logical_Operator_out3751_out1            : std_logic;
  SIGNAL Logical_Operator_out3752_out1            : std_logic;
  SIGNAL Logical_Operator_out3753_out1            : std_logic;
  SIGNAL Logical_Operator_out3754_out1            : std_logic;
  SIGNAL Logical_Operator_out3755_out1            : std_logic;
  SIGNAL Logical_Operator_out3756_out1            : std_logic;
  SIGNAL Logical_Operator_out3757_out1            : std_logic;
  SIGNAL Logical_Operator_out3758_out1            : std_logic;
  SIGNAL Logical_Operator_out3759_out1            : std_logic;
  SIGNAL Logical_Operator_out3760_out1            : std_logic;
  SIGNAL Logical_Operator_out3761_out1            : std_logic;
  SIGNAL Logical_Operator_out3762_out1            : std_logic;
  SIGNAL Logical_Operator_out3763_out1            : std_logic;
  SIGNAL Logical_Operator_out3764_out1            : std_logic;
  SIGNAL Logical_Operator_out3765_out1            : std_logic;
  SIGNAL Logical_Operator_out3766_out1            : std_logic;
  SIGNAL Logical_Operator_out3767_out1            : std_logic;
  SIGNAL Logical_Operator_out3768_out1            : std_logic;
  SIGNAL Logical_Operator_out3769_out1            : std_logic;
  SIGNAL Logical_Operator_out3770_out1            : std_logic;
  SIGNAL Logical_Operator_out3771_out1            : std_logic;
  SIGNAL Logical_Operator_out3772_out1            : std_logic;
  SIGNAL Logical_Operator_out3773_out1            : std_logic;
  SIGNAL Logical_Operator_out3774_out1            : std_logic;
  SIGNAL Logical_Operator_out3775_out1            : std_logic;
  SIGNAL Logical_Operator_out3776_out1            : std_logic;
  SIGNAL Logical_Operator_out3777_out1            : std_logic;
  SIGNAL Logical_Operator_out3778_out1            : std_logic;
  SIGNAL Logical_Operator_out3779_out1            : std_logic;
  SIGNAL Logical_Operator_out3780_out1            : std_logic;
  SIGNAL Logical_Operator_out3781_out1            : std_logic;
  SIGNAL Logical_Operator_out3782_out1            : std_logic;
  SIGNAL Logical_Operator_out3783_out1            : std_logic;
  SIGNAL Logical_Operator_out3784_out1            : std_logic;
  SIGNAL Logical_Operator_out3785_out1            : std_logic;
  SIGNAL Logical_Operator_out3786_out1            : std_logic;
  SIGNAL Logical_Operator_out3787_out1            : std_logic;
  SIGNAL Logical_Operator_out3788_out1            : std_logic;
  SIGNAL Logical_Operator_out3789_out1            : std_logic;
  SIGNAL Logical_Operator_out3790_out1            : std_logic;
  SIGNAL Logical_Operator_out3791_out1            : std_logic;
  SIGNAL Logical_Operator_out3792_out1            : std_logic;
  SIGNAL Logical_Operator_out3793_out1            : std_logic;
  SIGNAL Logical_Operator_out3794_out1            : std_logic;
  SIGNAL Logical_Operator_out3795_out1            : std_logic;
  SIGNAL Logical_Operator_out3796_out1            : std_logic;
  SIGNAL Logical_Operator_out3797_out1            : std_logic;
  SIGNAL Logical_Operator_out3798_out1            : std_logic;
  SIGNAL Logical_Operator_out3799_out1            : std_logic;
  SIGNAL Logical_Operator_out3800_out1            : std_logic;
  SIGNAL Logical_Operator_out3801_out1            : std_logic;
  SIGNAL Logical_Operator_out3802_out1            : std_logic;
  SIGNAL Logical_Operator_out3803_out1            : std_logic;
  SIGNAL Logical_Operator_out3804_out1            : std_logic;
  SIGNAL Logical_Operator_out3805_out1            : std_logic;
  SIGNAL Logical_Operator_out3806_out1            : std_logic;
  SIGNAL Logical_Operator_out3807_out1            : std_logic;
  SIGNAL Logical_Operator_out3808_out1            : std_logic;
  SIGNAL Logical_Operator_out3809_out1            : std_logic;
  SIGNAL Logical_Operator_out3810_out1            : std_logic;
  SIGNAL Logical_Operator_out3811_out1            : std_logic;
  SIGNAL Logical_Operator_out3812_out1            : std_logic;
  SIGNAL Logical_Operator_out3813_out1            : std_logic;
  SIGNAL Logical_Operator_out3814_out1            : std_logic;
  SIGNAL Logical_Operator_out3815_out1            : std_logic;
  SIGNAL Logical_Operator_out3816_out1            : std_logic;
  SIGNAL Logical_Operator_out3817_out1            : std_logic;
  SIGNAL Logical_Operator_out3818_out1            : std_logic;
  SIGNAL Logical_Operator_out3819_out1            : std_logic;
  SIGNAL Logical_Operator_out3820_out1            : std_logic;
  SIGNAL Logical_Operator_out3821_out1            : std_logic;
  SIGNAL Logical_Operator_out3822_out1            : std_logic;
  SIGNAL Logical_Operator_out3823_out1            : std_logic;
  SIGNAL Logical_Operator_out3824_out1            : std_logic;
  SIGNAL Logical_Operator_out3825_out1            : std_logic;
  SIGNAL Logical_Operator_out3826_out1            : std_logic;
  SIGNAL Logical_Operator_out3827_out1            : std_logic;
  SIGNAL Logical_Operator_out3828_out1            : std_logic;
  SIGNAL Logical_Operator_out3829_out1            : std_logic;
  SIGNAL Logical_Operator_out3830_out1            : std_logic;
  SIGNAL Logical_Operator_out3831_out1            : std_logic;
  SIGNAL Logical_Operator_out3832_out1            : std_logic;
  SIGNAL Logical_Operator_out3833_out1            : std_logic;
  SIGNAL Logical_Operator_out3834_out1            : std_logic;
  SIGNAL Logical_Operator_out3835_out1            : std_logic;
  SIGNAL Logical_Operator_out3836_out1            : std_logic;
  SIGNAL Logical_Operator_out3837_out1            : std_logic;
  SIGNAL Logical_Operator_out3838_out1            : std_logic;
  SIGNAL Logical_Operator_out3839_out1            : std_logic;
  SIGNAL Logical_Operator_out3840_out1            : std_logic;
  SIGNAL Logical_Operator_out3841_out1            : std_logic;
  SIGNAL Logical_Operator_out3842_out1            : std_logic;
  SIGNAL Logical_Operator_out3843_out1            : std_logic;
  SIGNAL Logical_Operator_out3844_out1            : std_logic;
  SIGNAL Logical_Operator_out3845_out1            : std_logic;
  SIGNAL Logical_Operator_out3846_out1            : std_logic;
  SIGNAL Logical_Operator_out3847_out1            : std_logic;
  SIGNAL Logical_Operator_out3848_out1            : std_logic;
  SIGNAL Logical_Operator_out3849_out1            : std_logic;
  SIGNAL Logical_Operator_out3850_out1            : std_logic;
  SIGNAL Logical_Operator_out3851_out1            : std_logic;
  SIGNAL Logical_Operator_out3852_out1            : std_logic;
  SIGNAL Logical_Operator_out3853_out1            : std_logic;
  SIGNAL Logical_Operator_out3854_out1            : std_logic;
  SIGNAL Logical_Operator_out3855_out1            : std_logic;
  SIGNAL Logical_Operator_out3856_out1            : std_logic;
  SIGNAL Logical_Operator_out3857_out1            : std_logic;
  SIGNAL Logical_Operator_out3858_out1            : std_logic;
  SIGNAL Logical_Operator_out3859_out1            : std_logic;
  SIGNAL Logical_Operator_out3860_out1            : std_logic;
  SIGNAL Logical_Operator_out3861_out1            : std_logic;
  SIGNAL Logical_Operator_out3862_out1            : std_logic;
  SIGNAL Logical_Operator_out3863_out1            : std_logic;
  SIGNAL Logical_Operator_out3864_out1            : std_logic;
  SIGNAL Logical_Operator_out3865_out1            : std_logic;
  SIGNAL Logical_Operator_out3866_out1            : std_logic;
  SIGNAL Logical_Operator_out3867_out1            : std_logic;
  SIGNAL Logical_Operator_out3868_out1            : std_logic;
  SIGNAL Logical_Operator_out3869_out1            : std_logic;
  SIGNAL Logical_Operator_out3870_out1            : std_logic;
  SIGNAL Logical_Operator_out3871_out1            : std_logic;
  SIGNAL Logical_Operator_out3872_out1            : std_logic;
  SIGNAL Logical_Operator_out3873_out1            : std_logic;
  SIGNAL Logical_Operator_out3874_out1            : std_logic;
  SIGNAL Logical_Operator_out3875_out1            : std_logic;
  SIGNAL Logical_Operator_out3876_out1            : std_logic;
  SIGNAL Logical_Operator_out3877_out1            : std_logic;
  SIGNAL Logical_Operator_out3878_out1            : std_logic;
  SIGNAL Logical_Operator_out3879_out1            : std_logic;
  SIGNAL Logical_Operator_out3880_out1            : std_logic;
  SIGNAL Logical_Operator_out3881_out1            : std_logic;
  SIGNAL Logical_Operator_out3882_out1            : std_logic;
  SIGNAL Logical_Operator_out3883_out1            : std_logic;
  SIGNAL Logical_Operator_out3884_out1            : std_logic;
  SIGNAL Logical_Operator_out3885_out1            : std_logic;
  SIGNAL Logical_Operator_out3886_out1            : std_logic;
  SIGNAL Logical_Operator_out3887_out1            : std_logic;
  SIGNAL Logical_Operator_out3888_out1            : std_logic;
  SIGNAL Logical_Operator_out3889_out1            : std_logic;
  SIGNAL Logical_Operator_out3890_out1            : std_logic;
  SIGNAL Logical_Operator_out3891_out1            : std_logic;
  SIGNAL Logical_Operator_out3892_out1            : std_logic;
  SIGNAL Logical_Operator_out3893_out1            : std_logic;
  SIGNAL Logical_Operator_out3894_out1            : std_logic;
  SIGNAL Logical_Operator_out3895_out1            : std_logic;
  SIGNAL Logical_Operator_out3896_out1            : std_logic;
  SIGNAL Logical_Operator_out3897_out1            : std_logic;
  SIGNAL Logical_Operator_out3898_out1            : std_logic;
  SIGNAL Logical_Operator_out3899_out1            : std_logic;
  SIGNAL Logical_Operator_out3900_out1            : std_logic;
  SIGNAL Logical_Operator_out3901_out1            : std_logic;
  SIGNAL Logical_Operator_out3902_out1            : std_logic;
  SIGNAL Logical_Operator_out3903_out1            : std_logic;
  SIGNAL Logical_Operator_out3904_out1            : std_logic;
  SIGNAL Logical_Operator_out3905_out1            : std_logic;
  SIGNAL Logical_Operator_out3906_out1            : std_logic;
  SIGNAL Logical_Operator_out3907_out1            : std_logic;
  SIGNAL Logical_Operator_out3908_out1            : std_logic;
  SIGNAL Logical_Operator_out3909_out1            : std_logic;
  SIGNAL Logical_Operator_out3910_out1            : std_logic;
  SIGNAL Logical_Operator_out3911_out1            : std_logic;
  SIGNAL Logical_Operator_out3912_out1            : std_logic;
  SIGNAL Logical_Operator_out3913_out1            : std_logic;
  SIGNAL Logical_Operator_out3914_out1            : std_logic;
  SIGNAL Logical_Operator_out3915_out1            : std_logic;
  SIGNAL Logical_Operator_out3916_out1            : std_logic;
  SIGNAL Logical_Operator_out3917_out1            : std_logic;
  SIGNAL Logical_Operator_out3918_out1            : std_logic;
  SIGNAL Logical_Operator_out3919_out1            : std_logic;
  SIGNAL Logical_Operator_out3920_out1            : std_logic;
  SIGNAL Logical_Operator_out3921_out1            : std_logic;
  SIGNAL Logical_Operator_out3922_out1            : std_logic;
  SIGNAL Logical_Operator_out3923_out1            : std_logic;
  SIGNAL Logical_Operator_out3924_out1            : std_logic;
  SIGNAL Logical_Operator_out3925_out1            : std_logic;
  SIGNAL Logical_Operator_out3926_out1            : std_logic;
  SIGNAL Logical_Operator_out3927_out1            : std_logic;
  SIGNAL Logical_Operator_out3928_out1            : std_logic;
  SIGNAL Logical_Operator_out3929_out1            : std_logic;
  SIGNAL Logical_Operator_out3930_out1            : std_logic;
  SIGNAL Logical_Operator_out3931_out1            : std_logic;
  SIGNAL Logical_Operator_out3932_out1            : std_logic;
  SIGNAL Logical_Operator_out3933_out1            : std_logic;
  SIGNAL Logical_Operator_out3934_out1            : std_logic;
  SIGNAL Logical_Operator_out3935_out1            : std_logic;
  SIGNAL Logical_Operator_out3936_out1            : std_logic;
  SIGNAL Logical_Operator_out3937_out1            : std_logic;
  SIGNAL Logical_Operator_out3938_out1            : std_logic;
  SIGNAL Logical_Operator_out3939_out1            : std_logic;
  SIGNAL Logical_Operator_out3940_out1            : std_logic;
  SIGNAL Logical_Operator_out3941_out1            : std_logic;
  SIGNAL Logical_Operator_out3942_out1            : std_logic;
  SIGNAL Logical_Operator_out3943_out1            : std_logic;
  SIGNAL Logical_Operator_out3944_out1            : std_logic;
  SIGNAL Logical_Operator_out3945_out1            : std_logic;
  SIGNAL Logical_Operator_out3946_out1            : std_logic;
  SIGNAL Logical_Operator_out3947_out1            : std_logic;
  SIGNAL Logical_Operator_out3948_out1            : std_logic;
  SIGNAL Logical_Operator_out3949_out1            : std_logic;
  SIGNAL Logical_Operator_out3950_out1            : std_logic;
  SIGNAL Logical_Operator_out3951_out1            : std_logic;
  SIGNAL Logical_Operator_out3952_out1            : std_logic;
  SIGNAL Logical_Operator_out3953_out1            : std_logic;
  SIGNAL Logical_Operator_out3954_out1            : std_logic;
  SIGNAL Logical_Operator_out3955_out1            : std_logic;
  SIGNAL Logical_Operator_out3956_out1            : std_logic;
  SIGNAL Logical_Operator_out3957_out1            : std_logic;
  SIGNAL Logical_Operator_out3958_out1            : std_logic;
  SIGNAL Logical_Operator_out3959_out1            : std_logic;
  SIGNAL Logical_Operator_out3960_out1            : std_logic;
  SIGNAL Logical_Operator_out3961_out1            : std_logic;
  SIGNAL Logical_Operator_out3962_out1            : std_logic;
  SIGNAL Logical_Operator_out3963_out1            : std_logic;
  SIGNAL Logical_Operator_out3964_out1            : std_logic;
  SIGNAL Logical_Operator_out3965_out1            : std_logic;
  SIGNAL Logical_Operator_out3966_out1            : std_logic;
  SIGNAL Logical_Operator_out3967_out1            : std_logic;
  SIGNAL Logical_Operator_out3968_out1            : std_logic;
  SIGNAL Logical_Operator_out3969_out1            : std_logic;
  SIGNAL Logical_Operator_out3970_out1            : std_logic;
  SIGNAL Logical_Operator_out3971_out1            : std_logic;
  SIGNAL Logical_Operator_out3972_out1            : std_logic;
  SIGNAL Logical_Operator_out3973_out1            : std_logic;
  SIGNAL Logical_Operator_out3974_out1            : std_logic;
  SIGNAL Logical_Operator_out3975_out1            : std_logic;
  SIGNAL Logical_Operator_out3976_out1            : std_logic;
  SIGNAL Logical_Operator_out3977_out1            : std_logic;
  SIGNAL Logical_Operator_out3978_out1            : std_logic;
  SIGNAL Logical_Operator_out3979_out1            : std_logic;
  SIGNAL Logical_Operator_out3980_out1            : std_logic;
  SIGNAL Logical_Operator_out3981_out1            : std_logic;
  SIGNAL Logical_Operator_out3982_out1            : std_logic;
  SIGNAL Logical_Operator_out3983_out1            : std_logic;
  SIGNAL Logical_Operator_out3984_out1            : std_logic;
  SIGNAL Logical_Operator_out3985_out1            : std_logic;
  SIGNAL Logical_Operator_out3986_out1            : std_logic;
  SIGNAL Logical_Operator_out3987_out1            : std_logic;
  SIGNAL Logical_Operator_out3988_out1            : std_logic;
  SIGNAL Logical_Operator_out3989_out1            : std_logic;
  SIGNAL Logical_Operator_out3990_out1            : std_logic;
  SIGNAL Logical_Operator_out3991_out1            : std_logic;
  SIGNAL Logical_Operator_out3992_out1            : std_logic;
  SIGNAL Logical_Operator_out3993_out1            : std_logic;
  SIGNAL Logical_Operator_out3994_out1            : std_logic;
  SIGNAL Logical_Operator_out3995_out1            : std_logic;
  SIGNAL Logical_Operator_out3996_out1            : std_logic;
  SIGNAL Logical_Operator_out3997_out1            : std_logic;
  SIGNAL Logical_Operator_out3998_out1            : std_logic;
  SIGNAL Logical_Operator_out3999_out1            : std_logic;
  SIGNAL Logical_Operator_out4000_out1            : std_logic;
  SIGNAL Logical_Operator_out4001_out1            : std_logic;
  SIGNAL Logical_Operator_out4002_out1            : std_logic;
  SIGNAL Logical_Operator_out4003_out1            : std_logic;
  SIGNAL Logical_Operator_out4004_out1            : std_logic;
  SIGNAL Logical_Operator_out4005_out1            : std_logic;
  SIGNAL Logical_Operator_out4006_out1            : std_logic;
  SIGNAL Logical_Operator_out4007_out1            : std_logic;
  SIGNAL Logical_Operator_out4008_out1            : std_logic;
  SIGNAL Logical_Operator_out4009_out1            : std_logic;
  SIGNAL Logical_Operator_out4010_out1            : std_logic;
  SIGNAL Logical_Operator_out4011_out1            : std_logic;
  SIGNAL Logical_Operator_out4012_out1            : std_logic;
  SIGNAL Logical_Operator_out4013_out1            : std_logic;
  SIGNAL Logical_Operator_out4014_out1            : std_logic;
  SIGNAL Logical_Operator_out4015_out1            : std_logic;
  SIGNAL Logical_Operator_out4016_out1            : std_logic;
  SIGNAL Logical_Operator_out4017_out1            : std_logic;
  SIGNAL Logical_Operator_out4018_out1            : std_logic;
  SIGNAL Logical_Operator_out4019_out1            : std_logic;
  SIGNAL Logical_Operator_out4020_out1            : std_logic;
  SIGNAL Logical_Operator_out4021_out1            : std_logic;
  SIGNAL Logical_Operator_out4022_out1            : std_logic;
  SIGNAL Logical_Operator_out4023_out1            : std_logic;
  SIGNAL Logical_Operator_out4024_out1            : std_logic;
  SIGNAL Logical_Operator_out4025_out1            : std_logic;
  SIGNAL Logical_Operator_out4026_out1            : std_logic;
  SIGNAL Logical_Operator_out4027_out1            : std_logic;
  SIGNAL Logical_Operator_out4028_out1            : std_logic;
  SIGNAL Logical_Operator_out4029_out1            : std_logic;
  SIGNAL Logical_Operator_out4030_out1            : std_logic;
  SIGNAL Logical_Operator_out4031_out1            : std_logic;
  SIGNAL Logical_Operator_out4032_out1            : std_logic;
  SIGNAL Logical_Operator_out4033_out1            : std_logic;
  SIGNAL Logical_Operator_out4034_out1            : std_logic;
  SIGNAL Logical_Operator_out4035_out1            : std_logic;
  SIGNAL Logical_Operator_out4036_out1            : std_logic;
  SIGNAL Logical_Operator_out4037_out1            : std_logic;
  SIGNAL Logical_Operator_out4038_out1            : std_logic;
  SIGNAL Logical_Operator_out4039_out1            : std_logic;
  SIGNAL Logical_Operator_out4040_out1            : std_logic;
  SIGNAL Logical_Operator_out4041_out1            : std_logic;
  SIGNAL Logical_Operator_out4042_out1            : std_logic;
  SIGNAL Logical_Operator_out4043_out1            : std_logic;
  SIGNAL Logical_Operator_out4044_out1            : std_logic;
  SIGNAL Logical_Operator_out4045_out1            : std_logic;
  SIGNAL Logical_Operator_out4046_out1            : std_logic;
  SIGNAL Logical_Operator_out4047_out1            : std_logic;
  SIGNAL Logical_Operator_out4048_out1            : std_logic;
  SIGNAL Logical_Operator_out4049_out1            : std_logic;
  SIGNAL Logical_Operator_out4050_out1            : std_logic;
  SIGNAL Logical_Operator_out4051_out1            : std_logic;
  SIGNAL Logical_Operator_out4052_out1            : std_logic;
  SIGNAL Logical_Operator_out4053_out1            : std_logic;
  SIGNAL Logical_Operator_out4054_out1            : std_logic;
  SIGNAL Logical_Operator_out4055_out1            : std_logic;
  SIGNAL Logical_Operator_out4056_out1            : std_logic;
  SIGNAL Logical_Operator_out4057_out1            : std_logic;
  SIGNAL Logical_Operator_out4058_out1            : std_logic;
  SIGNAL Logical_Operator_out4059_out1            : std_logic;
  SIGNAL Logical_Operator_out4060_out1            : std_logic;
  SIGNAL Logical_Operator_out4061_out1            : std_logic;
  SIGNAL Logical_Operator_out4062_out1            : std_logic;
  SIGNAL Logical_Operator_out4063_out1            : std_logic;
  SIGNAL Logical_Operator_out4064_out1            : std_logic;
  SIGNAL Logical_Operator_out4065_out1            : std_logic;
  SIGNAL Logical_Operator_out4066_out1            : std_logic;
  SIGNAL Logical_Operator_out4067_out1            : std_logic;
  SIGNAL Logical_Operator_out4068_out1            : std_logic;
  SIGNAL Logical_Operator_out4069_out1            : std_logic;
  SIGNAL Logical_Operator_out4070_out1            : std_logic;
  SIGNAL Logical_Operator_out4071_out1            : std_logic;
  SIGNAL Logical_Operator_out4072_out1            : std_logic;
  SIGNAL Logical_Operator_out4073_out1            : std_logic;
  SIGNAL Logical_Operator_out4074_out1            : std_logic;
  SIGNAL Logical_Operator_out4075_out1            : std_logic;
  SIGNAL Logical_Operator_out4076_out1            : std_logic;
  SIGNAL Logical_Operator_out4077_out1            : std_logic;
  SIGNAL Logical_Operator_out4078_out1            : std_logic;
  SIGNAL Logical_Operator_out4079_out1            : std_logic;
  SIGNAL Logical_Operator_out4080_out1            : std_logic;
  SIGNAL Logical_Operator_out4081_out1            : std_logic;
  SIGNAL Logical_Operator_out4082_out1            : std_logic;
  SIGNAL Logical_Operator_out4083_out1            : std_logic;
  SIGNAL Logical_Operator_out4084_out1            : std_logic;
  SIGNAL Logical_Operator_out4085_out1            : std_logic;
  SIGNAL Logical_Operator_out4086_out1            : std_logic;
  SIGNAL Logical_Operator_out4087_out1            : std_logic;
  SIGNAL Logical_Operator_out4088_out1            : std_logic;
  SIGNAL Logical_Operator_out4089_out1            : std_logic;
  SIGNAL Logical_Operator_out4090_out1            : std_logic;
  SIGNAL Logical_Operator_out4091_out1            : std_logic;
  SIGNAL Logical_Operator_out4092_out1            : std_logic;
  SIGNAL Logical_Operator_out4093_out1            : std_logic;
  SIGNAL Logical_Operator_out4094_out1            : std_logic;
  SIGNAL Logical_Operator_out4095_out1            : std_logic;
  SIGNAL Logical_Operator_out4096_out1            : std_logic;
  SIGNAL Logical_Operator_out4097_out1            : std_logic;
  SIGNAL Logical_Operator_out4098_out1            : std_logic;
  SIGNAL Logical_Operator_out4099_out1            : std_logic;
  SIGNAL Logical_Operator_out4100_out1            : std_logic;
  SIGNAL Logical_Operator_out4101_out1            : std_logic;
  SIGNAL Logical_Operator_out4102_out1            : std_logic;
  SIGNAL Logical_Operator_out4103_out1            : std_logic;
  SIGNAL Logical_Operator_out4104_out1            : std_logic;
  SIGNAL Logical_Operator_out4105_out1            : std_logic;
  SIGNAL Logical_Operator_out4106_out1            : std_logic;
  SIGNAL Logical_Operator_out4107_out1            : std_logic;
  SIGNAL Logical_Operator_out4108_out1            : std_logic;
  SIGNAL Logical_Operator_out4109_out1            : std_logic;
  SIGNAL Logical_Operator_out4110_out1            : std_logic;
  SIGNAL Logical_Operator_out4111_out1            : std_logic;
  SIGNAL Logical_Operator_out4112_out1            : std_logic;
  SIGNAL Logical_Operator_out4113_out1            : std_logic;
  SIGNAL Logical_Operator_out4114_out1            : std_logic;
  SIGNAL Logical_Operator_out4115_out1            : std_logic;
  SIGNAL Logical_Operator_out4116_out1            : std_logic;
  SIGNAL Logical_Operator_out4117_out1            : std_logic;
  SIGNAL Logical_Operator_out4118_out1            : std_logic;
  SIGNAL Logical_Operator_out4119_out1            : std_logic;
  SIGNAL Logical_Operator_out4120_out1            : std_logic;
  SIGNAL Logical_Operator_out4121_out1            : std_logic;
  SIGNAL Logical_Operator_out4122_out1            : std_logic;
  SIGNAL Logical_Operator_out4123_out1            : std_logic;
  SIGNAL Logical_Operator_out4124_out1            : std_logic;
  SIGNAL Logical_Operator_out4125_out1            : std_logic;
  SIGNAL Logical_Operator_out4126_out1            : std_logic;
  SIGNAL Logical_Operator_out4127_out1            : std_logic;
  SIGNAL Logical_Operator_out4128_out1            : std_logic;
  SIGNAL Logical_Operator_out4129_out1            : std_logic;
  SIGNAL Logical_Operator_out4130_out1            : std_logic;
  SIGNAL Logical_Operator_out4131_out1            : std_logic;
  SIGNAL Logical_Operator_out4132_out1            : std_logic;
  SIGNAL Logical_Operator_out4133_out1            : std_logic;
  SIGNAL Logical_Operator_out4134_out1            : std_logic;
  SIGNAL Logical_Operator_out4135_out1            : std_logic;
  SIGNAL Logical_Operator_out4136_out1            : std_logic;
  SIGNAL Logical_Operator_out4137_out1            : std_logic;
  SIGNAL Logical_Operator_out4138_out1            : std_logic;
  SIGNAL Logical_Operator_out4139_out1            : std_logic;
  SIGNAL Logical_Operator_out4140_out1            : std_logic;
  SIGNAL Logical_Operator_out4141_out1            : std_logic;
  SIGNAL Logical_Operator_out4142_out1            : std_logic;
  SIGNAL Logical_Operator_out4143_out1            : std_logic;
  SIGNAL Logical_Operator_out4144_out1            : std_logic;
  SIGNAL Logical_Operator_out4145_out1            : std_logic;
  SIGNAL Logical_Operator_out4146_out1            : std_logic;
  SIGNAL Logical_Operator_out4147_out1            : std_logic;
  SIGNAL Logical_Operator_out4148_out1            : std_logic;
  SIGNAL Logical_Operator_out4149_out1            : std_logic;
  SIGNAL Logical_Operator_out4150_out1            : std_logic;
  SIGNAL Logical_Operator_out4151_out1            : std_logic;
  SIGNAL Logical_Operator_out4152_out1            : std_logic;
  SIGNAL Logical_Operator_out4153_out1            : std_logic;
  SIGNAL Logical_Operator_out4154_out1            : std_logic;
  SIGNAL Logical_Operator_out4155_out1            : std_logic;
  SIGNAL Logical_Operator_out4156_out1            : std_logic;
  SIGNAL Logical_Operator_out4157_out1            : std_logic;
  SIGNAL Logical_Operator_out4158_out1            : std_logic;
  SIGNAL Logical_Operator_out4159_out1            : std_logic;
  SIGNAL Logical_Operator_out4160_out1            : std_logic;
  SIGNAL Logical_Operator_out4161_out1            : std_logic;
  SIGNAL Logical_Operator_out4162_out1            : std_logic;
  SIGNAL Logical_Operator_out4163_out1            : std_logic;
  SIGNAL Logical_Operator_out4164_out1            : std_logic;
  SIGNAL Logical_Operator_out4165_out1            : std_logic;
  SIGNAL Logical_Operator_out4166_out1            : std_logic;
  SIGNAL Logical_Operator_out4167_out1            : std_logic;
  SIGNAL Logical_Operator_out4168_out1            : std_logic;
  SIGNAL Logical_Operator_out4169_out1            : std_logic;
  SIGNAL Logical_Operator_out4170_out1            : std_logic;
  SIGNAL Logical_Operator_out4171_out1            : std_logic;
  SIGNAL Logical_Operator_out4172_out1            : std_logic;
  SIGNAL Logical_Operator_out4173_out1            : std_logic;
  SIGNAL Logical_Operator_out4174_out1            : std_logic;
  SIGNAL Logical_Operator_out4175_out1            : std_logic;
  SIGNAL Logical_Operator_out4176_out1            : std_logic;
  SIGNAL Logical_Operator_out4177_out1            : std_logic;
  SIGNAL Logical_Operator_out4178_out1            : std_logic;
  SIGNAL Logical_Operator_out4179_out1            : std_logic;
  SIGNAL Logical_Operator_out4180_out1            : std_logic;
  SIGNAL Logical_Operator_out4181_out1            : std_logic;
  SIGNAL Logical_Operator_out4182_out1            : std_logic;
  SIGNAL Logical_Operator_out4183_out1            : std_logic;
  SIGNAL Logical_Operator_out4184_out1            : std_logic;
  SIGNAL Logical_Operator_out4185_out1            : std_logic;
  SIGNAL Logical_Operator_out4186_out1            : std_logic;
  SIGNAL Logical_Operator_out4187_out1            : std_logic;
  SIGNAL Logical_Operator_out4188_out1            : std_logic;
  SIGNAL Logical_Operator_out4189_out1            : std_logic;
  SIGNAL Logical_Operator_out4190_out1            : std_logic;
  SIGNAL Logical_Operator_out4191_out1            : std_logic;
  SIGNAL Logical_Operator_out4192_out1            : std_logic;
  SIGNAL Logical_Operator_out4193_out1            : std_logic;
  SIGNAL Logical_Operator_out4194_out1            : std_logic;
  SIGNAL Logical_Operator_out4195_out1            : std_logic;
  SIGNAL Logical_Operator_out4196_out1            : std_logic;
  SIGNAL Logical_Operator_out4197_out1            : std_logic;
  SIGNAL Logical_Operator_out4198_out1            : std_logic;
  SIGNAL Logical_Operator_out4199_out1            : std_logic;
  SIGNAL Logical_Operator_out4200_out1            : std_logic;
  SIGNAL Logical_Operator_out4201_out1            : std_logic;
  SIGNAL Logical_Operator_out4202_out1            : std_logic;
  SIGNAL Logical_Operator_out4203_out1            : std_logic;
  SIGNAL Logical_Operator_out4204_out1            : std_logic;
  SIGNAL Logical_Operator_out4205_out1            : std_logic;
  SIGNAL Logical_Operator_out4206_out1            : std_logic;
  SIGNAL Logical_Operator_out4207_out1            : std_logic;
  SIGNAL Logical_Operator_out4208_out1            : std_logic;
  SIGNAL Logical_Operator_out4209_out1            : std_logic;
  SIGNAL Logical_Operator_out4210_out1            : std_logic;
  SIGNAL Logical_Operator_out4211_out1            : std_logic;
  SIGNAL Logical_Operator_out4212_out1            : std_logic;
  SIGNAL Logical_Operator_out4213_out1            : std_logic;
  SIGNAL Logical_Operator_out4214_out1            : std_logic;
  SIGNAL Logical_Operator_out4215_out1            : std_logic;
  SIGNAL Logical_Operator_out4216_out1            : std_logic;
  SIGNAL Logical_Operator_out4217_out1            : std_logic;
  SIGNAL Logical_Operator_out4218_out1            : std_logic;
  SIGNAL Logical_Operator_out4219_out1            : std_logic;
  SIGNAL Logical_Operator_out4220_out1            : std_logic;
  SIGNAL Logical_Operator_out4221_out1            : std_logic;
  SIGNAL Logical_Operator_out4222_out1            : std_logic;
  SIGNAL Logical_Operator_out4223_out1            : std_logic;
  SIGNAL Logical_Operator_out4224_out1            : std_logic;
  SIGNAL Logical_Operator_out4225_out1            : std_logic;
  SIGNAL Logical_Operator_out4226_out1            : std_logic;
  SIGNAL Logical_Operator_out4227_out1            : std_logic;
  SIGNAL Logical_Operator_out4228_out1            : std_logic;
  SIGNAL Logical_Operator_out4229_out1            : std_logic;
  SIGNAL Logical_Operator_out4230_out1            : std_logic;
  SIGNAL Logical_Operator_out4231_out1            : std_logic;
  SIGNAL Logical_Operator_out4232_out1            : std_logic;
  SIGNAL Logical_Operator_out4233_out1            : std_logic;
  SIGNAL Logical_Operator_out4234_out1            : std_logic;
  SIGNAL Logical_Operator_out4235_out1            : std_logic;
  SIGNAL Logical_Operator_out4236_out1            : std_logic;
  SIGNAL Logical_Operator_out4237_out1            : std_logic;
  SIGNAL Logical_Operator_out4238_out1            : std_logic;
  SIGNAL Logical_Operator_out4239_out1            : std_logic;
  SIGNAL Logical_Operator_out4240_out1            : std_logic;
  SIGNAL Logical_Operator_out4241_out1            : std_logic;
  SIGNAL Logical_Operator_out4242_out1            : std_logic;
  SIGNAL Logical_Operator_out4243_out1            : std_logic;
  SIGNAL Logical_Operator_out4244_out1            : std_logic;
  SIGNAL Logical_Operator_out4245_out1            : std_logic;
  SIGNAL Logical_Operator_out4246_out1            : std_logic;
  SIGNAL Logical_Operator_out4247_out1            : std_logic;
  SIGNAL Logical_Operator_out4248_out1            : std_logic;
  SIGNAL Logical_Operator_out4249_out1            : std_logic;
  SIGNAL Logical_Operator_out4250_out1            : std_logic;
  SIGNAL Logical_Operator_out4251_out1            : std_logic;
  SIGNAL Logical_Operator_out4252_out1            : std_logic;
  SIGNAL Logical_Operator_out4253_out1            : std_logic;
  SIGNAL Logical_Operator_out4254_out1            : std_logic;
  SIGNAL Logical_Operator_out4255_out1            : std_logic;
  SIGNAL Logical_Operator_out4256_out1            : std_logic;
  SIGNAL Logical_Operator_out4257_out1            : std_logic;
  SIGNAL Logical_Operator_out4258_out1            : std_logic;
  SIGNAL Logical_Operator_out4259_out1            : std_logic;
  SIGNAL Logical_Operator_out4260_out1            : std_logic;
  SIGNAL Logical_Operator_out4261_out1            : std_logic;
  SIGNAL Logical_Operator_out4262_out1            : std_logic;
  SIGNAL Logical_Operator_out4263_out1            : std_logic;
  SIGNAL Logical_Operator_out4264_out1            : std_logic;
  SIGNAL Logical_Operator_out4265_out1            : std_logic;
  SIGNAL Logical_Operator_out4266_out1            : std_logic;
  SIGNAL Logical_Operator_out4267_out1            : std_logic;
  SIGNAL Logical_Operator_out4268_out1            : std_logic;
  SIGNAL Logical_Operator_out4269_out1            : std_logic;
  SIGNAL Logical_Operator_out4270_out1            : std_logic;
  SIGNAL Logical_Operator_out4271_out1            : std_logic;
  SIGNAL Logical_Operator_out4272_out1            : std_logic;
  SIGNAL Logical_Operator_out4273_out1            : std_logic;
  SIGNAL Logical_Operator_out4274_out1            : std_logic;
  SIGNAL Logical_Operator_out4275_out1            : std_logic;
  SIGNAL Logical_Operator_out4276_out1            : std_logic;
  SIGNAL Logical_Operator_out4277_out1            : std_logic;
  SIGNAL Logical_Operator_out4278_out1            : std_logic;
  SIGNAL Logical_Operator_out4279_out1            : std_logic;
  SIGNAL Logical_Operator_out4280_out1            : std_logic;
  SIGNAL Logical_Operator_out4281_out1            : std_logic;
  SIGNAL Logical_Operator_out4282_out1            : std_logic;
  SIGNAL Logical_Operator_out4283_out1            : std_logic;
  SIGNAL Logical_Operator_out4284_out1            : std_logic;
  SIGNAL Logical_Operator_out4285_out1            : std_logic;
  SIGNAL Logical_Operator_out4286_out1            : std_logic;
  SIGNAL Logical_Operator_out4287_out1            : std_logic;
  SIGNAL Logical_Operator_out4288_out1            : std_logic;
  SIGNAL Logical_Operator_out4289_out1            : std_logic;
  SIGNAL Logical_Operator_out4290_out1            : std_logic;
  SIGNAL Logical_Operator_out4291_out1            : std_logic;
  SIGNAL Logical_Operator_out4292_out1            : std_logic;
  SIGNAL Logical_Operator_out4293_out1            : std_logic;
  SIGNAL Logical_Operator_out4294_out1            : std_logic;
  SIGNAL Logical_Operator_out4295_out1            : std_logic;
  SIGNAL Logical_Operator_out4296_out1            : std_logic;
  SIGNAL Logical_Operator_out4297_out1            : std_logic;
  SIGNAL Logical_Operator_out4298_out1            : std_logic;
  SIGNAL Logical_Operator_out4299_out1            : std_logic;
  SIGNAL Logical_Operator_out4300_out1            : std_logic;
  SIGNAL Logical_Operator_out4301_out1            : std_logic;
  SIGNAL Logical_Operator_out4302_out1            : std_logic;
  SIGNAL Logical_Operator_out4303_out1            : std_logic;
  SIGNAL Logical_Operator_out4304_out1            : std_logic;
  SIGNAL Logical_Operator_out4305_out1            : std_logic;
  SIGNAL Logical_Operator_out4306_out1            : std_logic;
  SIGNAL Logical_Operator_out4307_out1            : std_logic;
  SIGNAL Logical_Operator_out4308_out1            : std_logic;
  SIGNAL Logical_Operator_out4309_out1            : std_logic;
  SIGNAL Logical_Operator_out4310_out1            : std_logic;
  SIGNAL Logical_Operator_out4311_out1            : std_logic;
  SIGNAL Logical_Operator_out4312_out1            : std_logic;
  SIGNAL Logical_Operator_out4313_out1            : std_logic;
  SIGNAL Logical_Operator_out4314_out1            : std_logic;
  SIGNAL Logical_Operator_out4315_out1            : std_logic;
  SIGNAL Logical_Operator_out4316_out1            : std_logic;
  SIGNAL Logical_Operator_out4317_out1            : std_logic;
  SIGNAL Logical_Operator_out4318_out1            : std_logic;
  SIGNAL Logical_Operator_out4319_out1            : std_logic;
  SIGNAL Logical_Operator_out4320_out1            : std_logic;
  SIGNAL Logical_Operator_out4321_out1            : std_logic;
  SIGNAL Logical_Operator_out4322_out1            : std_logic;
  SIGNAL Logical_Operator_out4323_out1            : std_logic;
  SIGNAL Logical_Operator_out4324_out1            : std_logic;
  SIGNAL Logical_Operator_out4325_out1            : std_logic;
  SIGNAL Logical_Operator_out4326_out1            : std_logic;
  SIGNAL Logical_Operator_out4327_out1            : std_logic;
  SIGNAL Logical_Operator_out4328_out1            : std_logic;
  SIGNAL Logical_Operator_out4329_out1            : std_logic;
  SIGNAL Logical_Operator_out4330_out1            : std_logic;
  SIGNAL Logical_Operator_out4331_out1            : std_logic;
  SIGNAL Logical_Operator_out4332_out1            : std_logic;
  SIGNAL Logical_Operator_out4333_out1            : std_logic;
  SIGNAL Logical_Operator_out4334_out1            : std_logic;
  SIGNAL Logical_Operator_out4335_out1            : std_logic;
  SIGNAL Logical_Operator_out4336_out1            : std_logic;
  SIGNAL Logical_Operator_out4337_out1            : std_logic;
  SIGNAL Logical_Operator_out4338_out1            : std_logic;
  SIGNAL Logical_Operator_out4339_out1            : std_logic;
  SIGNAL Logical_Operator_out4340_out1            : std_logic;
  SIGNAL Logical_Operator_out4341_out1            : std_logic;
  SIGNAL Logical_Operator_out4342_out1            : std_logic;
  SIGNAL Logical_Operator_out4343_out1            : std_logic;
  SIGNAL Logical_Operator_out4344_out1            : std_logic;
  SIGNAL Logical_Operator_out4345_out1            : std_logic;
  SIGNAL Logical_Operator_out4346_out1            : std_logic;
  SIGNAL Logical_Operator_out4347_out1            : std_logic;
  SIGNAL Logical_Operator_out4348_out1            : std_logic;
  SIGNAL Logical_Operator_out4349_out1            : std_logic;
  SIGNAL Logical_Operator_out4350_out1            : std_logic;
  SIGNAL Logical_Operator_out4351_out1            : std_logic;
  SIGNAL Logical_Operator_out4352_out1            : std_logic;
  SIGNAL Logical_Operator_out4353_out1            : std_logic;
  SIGNAL Logical_Operator_out4354_out1            : std_logic;
  SIGNAL Logical_Operator_out4355_out1            : std_logic;
  SIGNAL Logical_Operator_out4356_out1            : std_logic;
  SIGNAL Logical_Operator_out4357_out1            : std_logic;
  SIGNAL Logical_Operator_out4358_out1            : std_logic;
  SIGNAL Logical_Operator_out4359_out1            : std_logic;
  SIGNAL Logical_Operator_out4360_out1            : std_logic;
  SIGNAL Logical_Operator_out4361_out1            : std_logic;
  SIGNAL Logical_Operator_out4362_out1            : std_logic;
  SIGNAL Logical_Operator_out4363_out1            : std_logic;
  SIGNAL Logical_Operator_out4364_out1            : std_logic;
  SIGNAL Logical_Operator_out4365_out1            : std_logic;
  SIGNAL Logical_Operator_out4366_out1            : std_logic;
  SIGNAL Logical_Operator_out4367_out1            : std_logic;
  SIGNAL Logical_Operator_out4368_out1            : std_logic;
  SIGNAL Logical_Operator_out4369_out1            : std_logic;
  SIGNAL Logical_Operator_out4370_out1            : std_logic;
  SIGNAL Logical_Operator_out4371_out1            : std_logic;
  SIGNAL Logical_Operator_out4372_out1            : std_logic;
  SIGNAL Logical_Operator_out4373_out1            : std_logic;
  SIGNAL Logical_Operator_out4374_out1            : std_logic;
  SIGNAL Logical_Operator_out4375_out1            : std_logic;
  SIGNAL Logical_Operator_out4376_out1            : std_logic;
  SIGNAL Logical_Operator_out4377_out1            : std_logic;
  SIGNAL Logical_Operator_out4378_out1            : std_logic;
  SIGNAL Logical_Operator_out4379_out1            : std_logic;
  SIGNAL Logical_Operator_out4380_out1            : std_logic;
  SIGNAL Logical_Operator_out4381_out1            : std_logic;
  SIGNAL Logical_Operator_out4382_out1            : std_logic;
  SIGNAL Logical_Operator_out4383_out1            : std_logic;
  SIGNAL Logical_Operator_out4384_out1            : std_logic;
  SIGNAL Logical_Operator_out4385_out1            : std_logic;
  SIGNAL Logical_Operator_out4386_out1            : std_logic;
  SIGNAL Logical_Operator_out4387_out1            : std_logic;
  SIGNAL Logical_Operator_out4388_out1            : std_logic;
  SIGNAL Logical_Operator_out4389_out1            : std_logic;
  SIGNAL Logical_Operator_out4390_out1            : std_logic;
  SIGNAL Logical_Operator_out4391_out1            : std_logic;
  SIGNAL Logical_Operator_out4392_out1            : std_logic;
  SIGNAL Logical_Operator_out4393_out1            : std_logic;
  SIGNAL Logical_Operator_out4394_out1            : std_logic;
  SIGNAL Logical_Operator_out4395_out1            : std_logic;
  SIGNAL Logical_Operator_out4396_out1            : std_logic;
  SIGNAL Logical_Operator_out4397_out1            : std_logic;
  SIGNAL Logical_Operator_out4398_out1            : std_logic;
  SIGNAL Logical_Operator_out4399_out1            : std_logic;
  SIGNAL Logical_Operator_out4400_out1            : std_logic;
  SIGNAL Logical_Operator_out4401_out1            : std_logic;
  SIGNAL Logical_Operator_out4402_out1            : std_logic;
  SIGNAL Logical_Operator_out4403_out1            : std_logic;
  SIGNAL Logical_Operator_out4404_out1            : std_logic;
  SIGNAL Logical_Operator_out4405_out1            : std_logic;
  SIGNAL Logical_Operator_out4406_out1            : std_logic;
  SIGNAL Logical_Operator_out4407_out1            : std_logic;
  SIGNAL Logical_Operator_out4408_out1            : std_logic;
  SIGNAL Logical_Operator_out4409_out1            : std_logic;
  SIGNAL Logical_Operator_out4410_out1            : std_logic;
  SIGNAL Logical_Operator_out4411_out1            : std_logic;
  SIGNAL Logical_Operator_out4412_out1            : std_logic;
  SIGNAL Logical_Operator_out4413_out1            : std_logic;
  SIGNAL Logical_Operator_out4414_out1            : std_logic;
  SIGNAL Logical_Operator_out4415_out1            : std_logic;
  SIGNAL Logical_Operator_out4416_out1            : std_logic;
  SIGNAL Logical_Operator_out4417_out1            : std_logic;
  SIGNAL Logical_Operator_out4418_out1            : std_logic;
  SIGNAL Logical_Operator_out4419_out1            : std_logic;
  SIGNAL Logical_Operator_out4420_out1            : std_logic;
  SIGNAL Logical_Operator_out4421_out1            : std_logic;
  SIGNAL Logical_Operator_out4422_out1            : std_logic;
  SIGNAL Logical_Operator_out4423_out1            : std_logic;
  SIGNAL Logical_Operator_out4424_out1            : std_logic;
  SIGNAL Logical_Operator_out4425_out1            : std_logic;
  SIGNAL Logical_Operator_out4426_out1            : std_logic;
  SIGNAL Logical_Operator_out4427_out1            : std_logic;
  SIGNAL Logical_Operator_out4428_out1            : std_logic;
  SIGNAL Logical_Operator_out4429_out1            : std_logic;
  SIGNAL Logical_Operator_out4430_out1            : std_logic;
  SIGNAL Logical_Operator_out4431_out1            : std_logic;
  SIGNAL Logical_Operator_out4432_out1            : std_logic;
  SIGNAL Logical_Operator_out4433_out1            : std_logic;
  SIGNAL Logical_Operator_out4434_out1            : std_logic;
  SIGNAL Logical_Operator_out4435_out1            : std_logic;
  SIGNAL Logical_Operator_out4436_out1            : std_logic;
  SIGNAL Logical_Operator_out4437_out1            : std_logic;
  SIGNAL Logical_Operator_out4438_out1            : std_logic;
  SIGNAL Logical_Operator_out4439_out1            : std_logic;
  SIGNAL Logical_Operator_out4440_out1            : std_logic;
  SIGNAL Logical_Operator_out4441_out1            : std_logic;
  SIGNAL Logical_Operator_out4442_out1            : std_logic;
  SIGNAL Logical_Operator_out4443_out1            : std_logic;
  SIGNAL Logical_Operator_out4444_out1            : std_logic;
  SIGNAL Logical_Operator_out4445_out1            : std_logic;
  SIGNAL Logical_Operator_out4446_out1            : std_logic;
  SIGNAL Logical_Operator_out4447_out1            : std_logic;
  SIGNAL Logical_Operator_out4448_out1            : std_logic;
  SIGNAL Logical_Operator_out4449_out1            : std_logic;
  SIGNAL Logical_Operator_out4450_out1            : std_logic;
  SIGNAL Logical_Operator_out4451_out1            : std_logic;
  SIGNAL Logical_Operator_out4452_out1            : std_logic;
  SIGNAL Logical_Operator_out4453_out1            : std_logic;
  SIGNAL Logical_Operator_out4454_out1            : std_logic;
  SIGNAL Logical_Operator_out4455_out1            : std_logic;
  SIGNAL Logical_Operator_out4456_out1            : std_logic;
  SIGNAL Logical_Operator_out4457_out1            : std_logic;
  SIGNAL Logical_Operator_out4458_out1            : std_logic;
  SIGNAL Logical_Operator_out4459_out1            : std_logic;
  SIGNAL Logical_Operator_out4460_out1            : std_logic;
  SIGNAL Logical_Operator_out4461_out1            : std_logic;
  SIGNAL Logical_Operator_out4462_out1            : std_logic;
  SIGNAL Logical_Operator_out4463_out1            : std_logic;
  SIGNAL Logical_Operator_out4464_out1            : std_logic;
  SIGNAL Logical_Operator_out4465_out1            : std_logic;
  SIGNAL Logical_Operator_out4466_out1            : std_logic;
  SIGNAL Logical_Operator_out4467_out1            : std_logic;
  SIGNAL Logical_Operator_out4468_out1            : std_logic;
  SIGNAL Logical_Operator_out4469_out1            : std_logic;
  SIGNAL Logical_Operator_out4470_out1            : std_logic;
  SIGNAL Logical_Operator_out4471_out1            : std_logic;
  SIGNAL Logical_Operator_out4472_out1            : std_logic;
  SIGNAL Logical_Operator_out4473_out1            : std_logic;
  SIGNAL Logical_Operator_out4474_out1            : std_logic;
  SIGNAL Logical_Operator_out4475_out1            : std_logic;
  SIGNAL Logical_Operator_out4476_out1            : std_logic;
  SIGNAL Logical_Operator_out4477_out1            : std_logic;
  SIGNAL Logical_Operator_out4478_out1            : std_logic;
  SIGNAL Logical_Operator_out4479_out1            : std_logic;
  SIGNAL Logical_Operator_out4480_out1            : std_logic;
  SIGNAL Logical_Operator_out4481_out1            : std_logic;
  SIGNAL Logical_Operator_out4482_out1            : std_logic;
  SIGNAL Logical_Operator_out4483_out1            : std_logic;
  SIGNAL Logical_Operator_out4484_out1            : std_logic;
  SIGNAL Logical_Operator_out4485_out1            : std_logic;
  SIGNAL Logical_Operator_out4486_out1            : std_logic;
  SIGNAL Logical_Operator_out4487_out1            : std_logic;
  SIGNAL Logical_Operator_out4488_out1            : std_logic;
  SIGNAL Logical_Operator_out4489_out1            : std_logic;
  SIGNAL Logical_Operator_out4490_out1            : std_logic;
  SIGNAL Logical_Operator_out4491_out1            : std_logic;
  SIGNAL Logical_Operator_out4492_out1            : std_logic;
  SIGNAL Logical_Operator_out4493_out1            : std_logic;
  SIGNAL Logical_Operator_out4494_out1            : std_logic;
  SIGNAL Logical_Operator_out4495_out1            : std_logic;
  SIGNAL Logical_Operator_out4496_out1            : std_logic;
  SIGNAL Logical_Operator_out4497_out1            : std_logic;
  SIGNAL Logical_Operator_out4498_out1            : std_logic;
  SIGNAL Logical_Operator_out4499_out1            : std_logic;
  SIGNAL Logical_Operator_out4500_out1            : std_logic;
  SIGNAL Logical_Operator_out4501_out1            : std_logic;
  SIGNAL Logical_Operator_out4502_out1            : std_logic;
  SIGNAL Logical_Operator_out4503_out1            : std_logic;
  SIGNAL Logical_Operator_out4504_out1            : std_logic;
  SIGNAL Logical_Operator_out4505_out1            : std_logic;
  SIGNAL Logical_Operator_out4506_out1            : std_logic;
  SIGNAL Logical_Operator_out4507_out1            : std_logic;
  SIGNAL Logical_Operator_out4508_out1            : std_logic;
  SIGNAL Logical_Operator_out4509_out1            : std_logic;
  SIGNAL Logical_Operator_out4510_out1            : std_logic;
  SIGNAL Logical_Operator_out4511_out1            : std_logic;
  SIGNAL Logical_Operator_out4512_out1            : std_logic;
  SIGNAL Logical_Operator_out4513_out1            : std_logic;
  SIGNAL Logical_Operator_out4514_out1            : std_logic;
  SIGNAL Logical_Operator_out4515_out1            : std_logic;
  SIGNAL Logical_Operator_out4516_out1            : std_logic;
  SIGNAL Logical_Operator_out4517_out1            : std_logic;
  SIGNAL Logical_Operator_out4518_out1            : std_logic;
  SIGNAL Logical_Operator_out4519_out1            : std_logic;
  SIGNAL Logical_Operator_out4520_out1            : std_logic;
  SIGNAL Logical_Operator_out4521_out1            : std_logic;
  SIGNAL Logical_Operator_out4522_out1            : std_logic;
  SIGNAL Logical_Operator_out4523_out1            : std_logic;
  SIGNAL Logical_Operator_out4524_out1            : std_logic;
  SIGNAL Logical_Operator_out4525_out1            : std_logic;
  SIGNAL Logical_Operator_out4526_out1            : std_logic;
  SIGNAL Logical_Operator_out4527_out1            : std_logic;
  SIGNAL Logical_Operator_out4528_out1            : std_logic;
  SIGNAL Logical_Operator_out4529_out1            : std_logic;
  SIGNAL Logical_Operator_out4530_out1            : std_logic;
  SIGNAL Logical_Operator_out4531_out1            : std_logic;
  SIGNAL Logical_Operator_out4532_out1            : std_logic;
  SIGNAL Logical_Operator_out4533_out1            : std_logic;
  SIGNAL Logical_Operator_out4534_out1            : std_logic;
  SIGNAL Logical_Operator_out4535_out1            : std_logic;
  SIGNAL Logical_Operator_out4536_out1            : std_logic;
  SIGNAL Logical_Operator_out4537_out1            : std_logic;
  SIGNAL Logical_Operator_out4538_out1            : std_logic;
  SIGNAL Logical_Operator_out4539_out1            : std_logic;
  SIGNAL Logical_Operator_out4540_out1            : std_logic;
  SIGNAL Logical_Operator_out4541_out1            : std_logic;
  SIGNAL Logical_Operator_out4542_out1            : std_logic;
  SIGNAL Logical_Operator_out4543_out1            : std_logic;
  SIGNAL Logical_Operator_out4544_out1            : std_logic;
  SIGNAL Logical_Operator_out4545_out1            : std_logic;
  SIGNAL Logical_Operator_out4546_out1            : std_logic;
  SIGNAL Logical_Operator_out4547_out1            : std_logic;
  SIGNAL Logical_Operator_out4548_out1            : std_logic;
  SIGNAL Logical_Operator_out4549_out1            : std_logic;
  SIGNAL Logical_Operator_out4550_out1            : std_logic;
  SIGNAL Logical_Operator_out4551_out1            : std_logic;
  SIGNAL Logical_Operator_out4552_out1            : std_logic;
  SIGNAL Logical_Operator_out4553_out1            : std_logic;
  SIGNAL Logical_Operator_out4554_out1            : std_logic;
  SIGNAL Logical_Operator_out4555_out1            : std_logic;
  SIGNAL Logical_Operator_out4556_out1            : std_logic;
  SIGNAL Logical_Operator_out4557_out1            : std_logic;
  SIGNAL Logical_Operator_out4558_out1            : std_logic;
  SIGNAL Logical_Operator_out4559_out1            : std_logic;
  SIGNAL Logical_Operator_out4560_out1            : std_logic;
  SIGNAL Logical_Operator_out4561_out1            : std_logic;
  SIGNAL Logical_Operator_out4562_out1            : std_logic;
  SIGNAL Logical_Operator_out4563_out1            : std_logic;
  SIGNAL Logical_Operator_out4564_out1            : std_logic;
  SIGNAL Logical_Operator_out4565_out1            : std_logic;
  SIGNAL Logical_Operator_out4566_out1            : std_logic;
  SIGNAL Logical_Operator_out4567_out1            : std_logic;
  SIGNAL Logical_Operator_out4568_out1            : std_logic;
  SIGNAL Logical_Operator_out4569_out1            : std_logic;
  SIGNAL Logical_Operator_out4570_out1            : std_logic;
  SIGNAL Logical_Operator_out4571_out1            : std_logic;
  SIGNAL Logical_Operator_out4572_out1            : std_logic;
  SIGNAL Logical_Operator_out4573_out1            : std_logic;
  SIGNAL Logical_Operator_out4574_out1            : std_logic;
  SIGNAL Logical_Operator_out4575_out1            : std_logic;
  SIGNAL Logical_Operator_out4576_out1            : std_logic;
  SIGNAL Logical_Operator_out4577_out1            : std_logic;
  SIGNAL Logical_Operator_out4578_out1            : std_logic;
  SIGNAL Logical_Operator_out4579_out1            : std_logic;
  SIGNAL Logical_Operator_out4580_out1            : std_logic;
  SIGNAL Logical_Operator_out4581_out1            : std_logic;
  SIGNAL Logical_Operator_out4582_out1            : std_logic;
  SIGNAL Logical_Operator_out4583_out1            : std_logic;
  SIGNAL Logical_Operator_out4584_out1            : std_logic;
  SIGNAL Logical_Operator_out4585_out1            : std_logic;
  SIGNAL Logical_Operator_out4586_out1            : std_logic;
  SIGNAL Logical_Operator_out4587_out1            : std_logic;
  SIGNAL Logical_Operator_out4588_out1            : std_logic;
  SIGNAL Logical_Operator_out4589_out1            : std_logic;
  SIGNAL Logical_Operator_out4590_out1            : std_logic;
  SIGNAL Logical_Operator_out4591_out1            : std_logic;
  SIGNAL Logical_Operator_out4592_out1            : std_logic;
  SIGNAL Logical_Operator_out4593_out1            : std_logic;
  SIGNAL Logical_Operator_out4594_out1            : std_logic;
  SIGNAL Logical_Operator_out4595_out1            : std_logic;
  SIGNAL Logical_Operator_out4596_out1            : std_logic;
  SIGNAL Logical_Operator_out4597_out1            : std_logic;
  SIGNAL Logical_Operator_out4598_out1            : std_logic;
  SIGNAL Logical_Operator_out4599_out1            : std_logic;
  SIGNAL Logical_Operator_out4600_out1            : std_logic;
  SIGNAL Logical_Operator_out4601_out1            : std_logic;
  SIGNAL Logical_Operator_out4602_out1            : std_logic;
  SIGNAL Logical_Operator_out4603_out1            : std_logic;
  SIGNAL Logical_Operator_out4604_out1            : std_logic;
  SIGNAL Logical_Operator_out4605_out1            : std_logic;
  SIGNAL Logical_Operator_out4606_out1            : std_logic;
  SIGNAL Logical_Operator_out4607_out1            : std_logic;
  SIGNAL Logical_Operator_out4608_out1            : std_logic;
  SIGNAL Logical_Operator_out4609_out1            : std_logic;
  SIGNAL Logical_Operator_out4610_out1            : std_logic;
  SIGNAL Logical_Operator_out4611_out1            : std_logic;
  SIGNAL Logical_Operator_out4612_out1            : std_logic;
  SIGNAL Logical_Operator_out4613_out1            : std_logic;
  SIGNAL Logical_Operator_out4614_out1            : std_logic;
  SIGNAL Logical_Operator_out4615_out1            : std_logic;
  SIGNAL Logical_Operator_out4616_out1            : std_logic;
  SIGNAL Logical_Operator_out4617_out1            : std_logic;
  SIGNAL Logical_Operator_out4618_out1            : std_logic;
  SIGNAL Logical_Operator_out4619_out1            : std_logic;
  SIGNAL Logical_Operator_out4620_out1            : std_logic;
  SIGNAL Logical_Operator_out4621_out1            : std_logic;
  SIGNAL Logical_Operator_out4622_out1            : std_logic;
  SIGNAL Logical_Operator_out4623_out1            : std_logic;
  SIGNAL Logical_Operator_out4624_out1            : std_logic;
  SIGNAL Logical_Operator_out4625_out1            : std_logic;
  SIGNAL Logical_Operator_out4626_out1            : std_logic;
  SIGNAL Logical_Operator_out4627_out1            : std_logic;
  SIGNAL Logical_Operator_out4628_out1            : std_logic;
  SIGNAL Logical_Operator_out4629_out1            : std_logic;
  SIGNAL Logical_Operator_out4630_out1            : std_logic;
  SIGNAL Logical_Operator_out4631_out1            : std_logic;
  SIGNAL Logical_Operator_out4632_out1            : std_logic;
  SIGNAL Logical_Operator_out4633_out1            : std_logic;
  SIGNAL Logical_Operator_out4634_out1            : std_logic;
  SIGNAL Logical_Operator_out4635_out1            : std_logic;
  SIGNAL Logical_Operator_out4636_out1            : std_logic;
  SIGNAL Logical_Operator_out4637_out1            : std_logic;
  SIGNAL Logical_Operator_out4638_out1            : std_logic;
  SIGNAL Logical_Operator_out4639_out1            : std_logic;
  SIGNAL Logical_Operator_out4640_out1            : std_logic;
  SIGNAL Logical_Operator_out4641_out1            : std_logic;
  SIGNAL Logical_Operator_out4642_out1            : std_logic;
  SIGNAL Logical_Operator_out4643_out1            : std_logic;
  SIGNAL Logical_Operator_out4644_out1            : std_logic;
  SIGNAL Logical_Operator_out4645_out1            : std_logic;
  SIGNAL Logical_Operator_out4646_out1            : std_logic;
  SIGNAL Logical_Operator_out4647_out1            : std_logic;
  SIGNAL Logical_Operator_out4648_out1            : std_logic;
  SIGNAL Logical_Operator_out4649_out1            : std_logic;
  SIGNAL Logical_Operator_out4650_out1            : std_logic;
  SIGNAL Logical_Operator_out4651_out1            : std_logic;
  SIGNAL Logical_Operator_out4652_out1            : std_logic;
  SIGNAL Logical_Operator_out4653_out1            : std_logic;
  SIGNAL Logical_Operator_out4654_out1            : std_logic;
  SIGNAL Logical_Operator_out4655_out1            : std_logic;
  SIGNAL Logical_Operator_out4656_out1            : std_logic;
  SIGNAL Logical_Operator_out4657_out1            : std_logic;
  SIGNAL Logical_Operator_out4658_out1            : std_logic;
  SIGNAL Logical_Operator_out4659_out1            : std_logic;
  SIGNAL Logical_Operator_out4660_out1            : std_logic;
  SIGNAL Logical_Operator_out4661_out1            : std_logic;
  SIGNAL Logical_Operator_out4662_out1            : std_logic;
  SIGNAL Logical_Operator_out4663_out1            : std_logic;
  SIGNAL Logical_Operator_out4664_out1            : std_logic;
  SIGNAL Logical_Operator_out4665_out1            : std_logic;
  SIGNAL Logical_Operator_out4666_out1            : std_logic;
  SIGNAL Logical_Operator_out4667_out1            : std_logic;
  SIGNAL Logical_Operator_out4668_out1            : std_logic;
  SIGNAL Logical_Operator_out4669_out1            : std_logic;
  SIGNAL Logical_Operator_out4670_out1            : std_logic;
  SIGNAL Logical_Operator_out4671_out1            : std_logic;
  SIGNAL Logical_Operator_out4672_out1            : std_logic;
  SIGNAL Logical_Operator_out4673_out1            : std_logic;
  SIGNAL Logical_Operator_out4674_out1            : std_logic;
  SIGNAL Logical_Operator_out4675_out1            : std_logic;
  SIGNAL Logical_Operator_out4676_out1            : std_logic;
  SIGNAL Logical_Operator_out4677_out1            : std_logic;
  SIGNAL Logical_Operator_out4678_out1            : std_logic;
  SIGNAL Logical_Operator_out4679_out1            : std_logic;
  SIGNAL Logical_Operator_out4680_out1            : std_logic;
  SIGNAL Logical_Operator_out4681_out1            : std_logic;
  SIGNAL Logical_Operator_out4682_out1            : std_logic;
  SIGNAL Logical_Operator_out4683_out1            : std_logic;
  SIGNAL Logical_Operator_out4684_out1            : std_logic;
  SIGNAL Logical_Operator_out4685_out1            : std_logic;
  SIGNAL Logical_Operator_out4686_out1            : std_logic;
  SIGNAL Logical_Operator_out4687_out1            : std_logic;
  SIGNAL Logical_Operator_out4688_out1            : std_logic;
  SIGNAL Logical_Operator_out4689_out1            : std_logic;
  SIGNAL Logical_Operator_out4690_out1            : std_logic;
  SIGNAL Logical_Operator_out4691_out1            : std_logic;
  SIGNAL Logical_Operator_out4692_out1            : std_logic;
  SIGNAL Logical_Operator_out4693_out1            : std_logic;
  SIGNAL Logical_Operator_out4694_out1            : std_logic;
  SIGNAL Logical_Operator_out4695_out1            : std_logic;
  SIGNAL Logical_Operator_out4696_out1            : std_logic;
  SIGNAL Logical_Operator_out4697_out1            : std_logic;
  SIGNAL Logical_Operator_out4698_out1            : std_logic;
  SIGNAL Logical_Operator_out4699_out1            : std_logic;
  SIGNAL Logical_Operator_out4700_out1            : std_logic;
  SIGNAL Logical_Operator_out4701_out1            : std_logic;
  SIGNAL Logical_Operator_out4702_out1            : std_logic;
  SIGNAL Logical_Operator_out4703_out1            : std_logic;
  SIGNAL Logical_Operator_out4704_out1            : std_logic;
  SIGNAL Logical_Operator_out4705_out1            : std_logic;
  SIGNAL Logical_Operator_out4706_out1            : std_logic;
  SIGNAL Logical_Operator_out4707_out1            : std_logic;
  SIGNAL Logical_Operator_out4708_out1            : std_logic;
  SIGNAL Logical_Operator_out4709_out1            : std_logic;
  SIGNAL Logical_Operator_out4710_out1            : std_logic;
  SIGNAL Logical_Operator_out4711_out1            : std_logic;
  SIGNAL Logical_Operator_out4712_out1            : std_logic;
  SIGNAL Logical_Operator_out4713_out1            : std_logic;
  SIGNAL Logical_Operator_out4714_out1            : std_logic;
  SIGNAL Logical_Operator_out4715_out1            : std_logic;
  SIGNAL Logical_Operator_out4716_out1            : std_logic;
  SIGNAL Logical_Operator_out4717_out1            : std_logic;
  SIGNAL Logical_Operator_out4718_out1            : std_logic;
  SIGNAL Logical_Operator_out4719_out1            : std_logic;
  SIGNAL Logical_Operator_out4720_out1            : std_logic;
  SIGNAL Logical_Operator_out4721_out1            : std_logic;
  SIGNAL Logical_Operator_out4722_out1            : std_logic;
  SIGNAL Logical_Operator_out4723_out1            : std_logic;
  SIGNAL Logical_Operator_out4724_out1            : std_logic;
  SIGNAL Logical_Operator_out4725_out1            : std_logic;
  SIGNAL Logical_Operator_out4726_out1            : std_logic;
  SIGNAL Logical_Operator_out4727_out1            : std_logic;
  SIGNAL Logical_Operator_out4728_out1            : std_logic;
  SIGNAL Logical_Operator_out4729_out1            : std_logic;
  SIGNAL Logical_Operator_out4730_out1            : std_logic;
  SIGNAL Logical_Operator_out4731_out1            : std_logic;
  SIGNAL Logical_Operator_out4732_out1            : std_logic;
  SIGNAL Logical_Operator_out4733_out1            : std_logic;
  SIGNAL Logical_Operator_out4734_out1            : std_logic;
  SIGNAL Logical_Operator_out4735_out1            : std_logic;
  SIGNAL Logical_Operator_out4736_out1            : std_logic;
  SIGNAL Logical_Operator_out4737_out1            : std_logic;
  SIGNAL Logical_Operator_out4738_out1            : std_logic;
  SIGNAL Logical_Operator_out4739_out1            : std_logic;
  SIGNAL Logical_Operator_out4740_out1            : std_logic;
  SIGNAL Logical_Operator_out4741_out1            : std_logic;
  SIGNAL Logical_Operator_out4742_out1            : std_logic;
  SIGNAL Logical_Operator_out4743_out1            : std_logic;
  SIGNAL Logical_Operator_out4744_out1            : std_logic;
  SIGNAL Logical_Operator_out4745_out1            : std_logic;
  SIGNAL Logical_Operator_out4746_out1            : std_logic;
  SIGNAL Logical_Operator_out4747_out1            : std_logic;
  SIGNAL Logical_Operator_out4748_out1            : std_logic;
  SIGNAL Logical_Operator_out4749_out1            : std_logic;
  SIGNAL Logical_Operator_out4750_out1            : std_logic;
  SIGNAL Logical_Operator_out4751_out1            : std_logic;
  SIGNAL Logical_Operator_out4752_out1            : std_logic;
  SIGNAL Logical_Operator_out4753_out1            : std_logic;
  SIGNAL Logical_Operator_out4754_out1            : std_logic;
  SIGNAL Logical_Operator_out4755_out1            : std_logic;
  SIGNAL Logical_Operator_out4756_out1            : std_logic;
  SIGNAL Logical_Operator_out4757_out1            : std_logic;
  SIGNAL Logical_Operator_out4758_out1            : std_logic;
  SIGNAL Logical_Operator_out4759_out1            : std_logic;
  SIGNAL Logical_Operator_out4760_out1            : std_logic;
  SIGNAL Logical_Operator_out4761_out1            : std_logic;
  SIGNAL Logical_Operator_out4762_out1            : std_logic;
  SIGNAL Logical_Operator_out4763_out1            : std_logic;
  SIGNAL Logical_Operator_out4764_out1            : std_logic;
  SIGNAL Logical_Operator_out4765_out1            : std_logic;
  SIGNAL Logical_Operator_out4766_out1            : std_logic;
  SIGNAL Logical_Operator_out4767_out1            : std_logic;
  SIGNAL Logical_Operator_out4768_out1            : std_logic;
  SIGNAL Logical_Operator_out4769_out1            : std_logic;
  SIGNAL Logical_Operator_out4770_out1            : std_logic;
  SIGNAL Logical_Operator_out4771_out1            : std_logic;
  SIGNAL Logical_Operator_out4772_out1            : std_logic;
  SIGNAL Logical_Operator_out4773_out1            : std_logic;
  SIGNAL Logical_Operator_out4774_out1            : std_logic;
  SIGNAL Logical_Operator_out4775_out1            : std_logic;
  SIGNAL Logical_Operator_out4776_out1            : std_logic;
  SIGNAL Logical_Operator_out4777_out1            : std_logic;
  SIGNAL Logical_Operator_out4778_out1            : std_logic;
  SIGNAL Logical_Operator_out4779_out1            : std_logic;
  SIGNAL Logical_Operator_out4780_out1            : std_logic;
  SIGNAL Logical_Operator_out4781_out1            : std_logic;
  SIGNAL Logical_Operator_out4782_out1            : std_logic;
  SIGNAL Logical_Operator_out4783_out1            : std_logic;
  SIGNAL Logical_Operator_out4784_out1            : std_logic;
  SIGNAL Logical_Operator_out4785_out1            : std_logic;
  SIGNAL Logical_Operator_out4786_out1            : std_logic;
  SIGNAL Logical_Operator_out4787_out1            : std_logic;
  SIGNAL Logical_Operator_out4788_out1            : std_logic;
  SIGNAL Logical_Operator_out4789_out1            : std_logic;
  SIGNAL Logical_Operator_out4790_out1            : std_logic;
  SIGNAL Logical_Operator_out4791_out1            : std_logic;
  SIGNAL Logical_Operator_out4792_out1            : std_logic;
  SIGNAL Logical_Operator_out4793_out1            : std_logic;
  SIGNAL Logical_Operator_out4794_out1            : std_logic;
  SIGNAL Logical_Operator_out4795_out1            : std_logic;
  SIGNAL Logical_Operator_out4796_out1            : std_logic;
  SIGNAL Logical_Operator_out4797_out1            : std_logic;
  SIGNAL Logical_Operator_out4798_out1            : std_logic;
  SIGNAL Logical_Operator_out4799_out1            : std_logic;
  SIGNAL Logical_Operator_out4800_out1            : std_logic;
  SIGNAL Logical_Operator_out4801_out1            : std_logic;
  SIGNAL Logical_Operator_out4802_out1            : std_logic;
  SIGNAL Logical_Operator_out4803_out1            : std_logic;
  SIGNAL Logical_Operator_out4804_out1            : std_logic;
  SIGNAL Logical_Operator_out4805_out1            : std_logic;
  SIGNAL Logical_Operator_out4806_out1            : std_logic;
  SIGNAL Logical_Operator_out4807_out1            : std_logic;
  SIGNAL Logical_Operator_out4808_out1            : std_logic;
  SIGNAL Logical_Operator_out4809_out1            : std_logic;
  SIGNAL Logical_Operator_out4810_out1            : std_logic;
  SIGNAL Logical_Operator_out4811_out1            : std_logic;
  SIGNAL Logical_Operator_out4812_out1            : std_logic;
  SIGNAL Logical_Operator_out4813_out1            : std_logic;
  SIGNAL Logical_Operator_out4814_out1            : std_logic;
  SIGNAL Logical_Operator_out4815_out1            : std_logic;
  SIGNAL Logical_Operator_out4816_out1            : std_logic;
  SIGNAL Logical_Operator_out4817_out1            : std_logic;
  SIGNAL Logical_Operator_out4818_out1            : std_logic;
  SIGNAL Logical_Operator_out4819_out1            : std_logic;
  SIGNAL Logical_Operator_out4820_out1            : std_logic;
  SIGNAL Logical_Operator_out4821_out1            : std_logic;
  SIGNAL Logical_Operator_out4822_out1            : std_logic;
  SIGNAL Logical_Operator_out4823_out1            : std_logic;
  SIGNAL Logical_Operator_out4824_out1            : std_logic;
  SIGNAL Logical_Operator_out4825_out1            : std_logic;
  SIGNAL Logical_Operator_out4826_out1            : std_logic;
  SIGNAL Logical_Operator_out4827_out1            : std_logic;
  SIGNAL Logical_Operator_out4828_out1            : std_logic;
  SIGNAL Logical_Operator_out4829_out1            : std_logic;
  SIGNAL Logical_Operator_out4830_out1            : std_logic;
  SIGNAL Logical_Operator_out4831_out1            : std_logic;
  SIGNAL Logical_Operator_out4832_out1            : std_logic;
  SIGNAL Logical_Operator_out4833_out1            : std_logic;
  SIGNAL Logical_Operator_out4834_out1            : std_logic;
  SIGNAL Logical_Operator_out4835_out1            : std_logic;
  SIGNAL Logical_Operator_out4836_out1            : std_logic;
  SIGNAL Logical_Operator_out4837_out1            : std_logic;
  SIGNAL Logical_Operator_out4838_out1            : std_logic;
  SIGNAL Logical_Operator_out4839_out1            : std_logic;
  SIGNAL Logical_Operator_out4840_out1            : std_logic;
  SIGNAL Logical_Operator_out4841_out1            : std_logic;
  SIGNAL Logical_Operator_out4842_out1            : std_logic;
  SIGNAL Logical_Operator_out4843_out1            : std_logic;
  SIGNAL Logical_Operator_out4844_out1            : std_logic;
  SIGNAL Logical_Operator_out4845_out1            : std_logic;
  SIGNAL Logical_Operator_out4846_out1            : std_logic;
  SIGNAL Logical_Operator_out4847_out1            : std_logic;
  SIGNAL Logical_Operator_out4848_out1            : std_logic;
  SIGNAL Logical_Operator_out4849_out1            : std_logic;
  SIGNAL Logical_Operator_out4850_out1            : std_logic;
  SIGNAL Logical_Operator_out4851_out1            : std_logic;
  SIGNAL Logical_Operator_out4852_out1            : std_logic;
  SIGNAL Logical_Operator_out4853_out1            : std_logic;
  SIGNAL Logical_Operator_out4854_out1            : std_logic;
  SIGNAL Logical_Operator_out4855_out1            : std_logic;
  SIGNAL Logical_Operator_out4856_out1            : std_logic;
  SIGNAL Logical_Operator_out4857_out1            : std_logic;
  SIGNAL Logical_Operator_out4858_out1            : std_logic;
  SIGNAL Logical_Operator_out4859_out1            : std_logic;
  SIGNAL Logical_Operator_out4860_out1            : std_logic;
  SIGNAL Logical_Operator_out4861_out1            : std_logic;
  SIGNAL Logical_Operator_out4862_out1            : std_logic;
  SIGNAL Logical_Operator_out4863_out1            : std_logic;
  SIGNAL Logical_Operator_out4864_out1            : std_logic;
  SIGNAL Logical_Operator_out4865_out1            : std_logic;
  SIGNAL Logical_Operator_out4866_out1            : std_logic;
  SIGNAL Logical_Operator_out4867_out1            : std_logic;
  SIGNAL Logical_Operator_out4868_out1            : std_logic;
  SIGNAL Logical_Operator_out4869_out1            : std_logic;
  SIGNAL Logical_Operator_out4870_out1            : std_logic;
  SIGNAL Logical_Operator_out4871_out1            : std_logic;
  SIGNAL Logical_Operator_out4872_out1            : std_logic;
  SIGNAL Logical_Operator_out4873_out1            : std_logic;
  SIGNAL Logical_Operator_out4874_out1            : std_logic;
  SIGNAL Logical_Operator_out4875_out1            : std_logic;
  SIGNAL Logical_Operator_out4876_out1            : std_logic;
  SIGNAL Logical_Operator_out4877_out1            : std_logic;
  SIGNAL Logical_Operator_out4878_out1            : std_logic;
  SIGNAL Logical_Operator_out4879_out1            : std_logic;
  SIGNAL Logical_Operator_out4880_out1            : std_logic;
  SIGNAL Logical_Operator_out4881_out1            : std_logic;
  SIGNAL Logical_Operator_out4882_out1            : std_logic;
  SIGNAL Logical_Operator_out4883_out1            : std_logic;
  SIGNAL Logical_Operator_out4884_out1            : std_logic;
  SIGNAL Logical_Operator_out4885_out1            : std_logic;
  SIGNAL Logical_Operator_out4886_out1            : std_logic;
  SIGNAL Logical_Operator_out4887_out1            : std_logic;
  SIGNAL Logical_Operator_out4888_out1            : std_logic;
  SIGNAL Logical_Operator_out4889_out1            : std_logic;
  SIGNAL Logical_Operator_out4890_out1            : std_logic;
  SIGNAL Logical_Operator_out4891_out1            : std_logic;
  SIGNAL Logical_Operator_out4892_out1            : std_logic;
  SIGNAL Logical_Operator_out4893_out1            : std_logic;
  SIGNAL Logical_Operator_out4894_out1            : std_logic;
  SIGNAL Logical_Operator_out4895_out1            : std_logic;
  SIGNAL Logical_Operator_out4896_out1            : std_logic;
  SIGNAL Logical_Operator_out4897_out1            : std_logic;
  SIGNAL Logical_Operator_out4898_out1            : std_logic;
  SIGNAL Logical_Operator_out4899_out1            : std_logic;
  SIGNAL Logical_Operator_out4900_out1            : std_logic;
  SIGNAL Logical_Operator_out4901_out1            : std_logic;
  SIGNAL Logical_Operator_out4902_out1            : std_logic;
  SIGNAL Logical_Operator_out4903_out1            : std_logic;
  SIGNAL Logical_Operator_out4904_out1            : std_logic;
  SIGNAL Logical_Operator_out4905_out1            : std_logic;
  SIGNAL Logical_Operator_out4906_out1            : std_logic;
  SIGNAL Logical_Operator_out4907_out1            : std_logic;
  SIGNAL Logical_Operator_out4908_out1            : std_logic;
  SIGNAL Logical_Operator_out4909_out1            : std_logic;
  SIGNAL Logical_Operator_out4910_out1            : std_logic;
  SIGNAL Logical_Operator_out4911_out1            : std_logic;
  SIGNAL Logical_Operator_out4912_out1            : std_logic;
  SIGNAL Logical_Operator_out4913_out1            : std_logic;
  SIGNAL Logical_Operator_out4914_out1            : std_logic;
  SIGNAL Logical_Operator_out4915_out1            : std_logic;
  SIGNAL Logical_Operator_out4916_out1            : std_logic;
  SIGNAL Logical_Operator_out4917_out1            : std_logic;
  SIGNAL Logical_Operator_out4918_out1            : std_logic;
  SIGNAL Logical_Operator_out4919_out1            : std_logic;
  SIGNAL Logical_Operator_out4920_out1            : std_logic;
  SIGNAL Logical_Operator_out4921_out1            : std_logic;
  SIGNAL Logical_Operator_out4922_out1            : std_logic;
  SIGNAL Logical_Operator_out4923_out1            : std_logic;
  SIGNAL Logical_Operator_out4924_out1            : std_logic;
  SIGNAL Logical_Operator_out4925_out1            : std_logic;
  SIGNAL Logical_Operator_out4926_out1            : std_logic;
  SIGNAL Logical_Operator_out4927_out1            : std_logic;
  SIGNAL Logical_Operator_out4928_out1            : std_logic;
  SIGNAL Logical_Operator_out4929_out1            : std_logic;
  SIGNAL Logical_Operator_out4930_out1            : std_logic;
  SIGNAL Logical_Operator_out4931_out1            : std_logic;
  SIGNAL Logical_Operator_out4932_out1            : std_logic;
  SIGNAL Logical_Operator_out4933_out1            : std_logic;
  SIGNAL Logical_Operator_out4934_out1            : std_logic;
  SIGNAL Logical_Operator_out4935_out1            : std_logic;
  SIGNAL Logical_Operator_out4936_out1            : std_logic;
  SIGNAL Logical_Operator_out4937_out1            : std_logic;
  SIGNAL Logical_Operator_out4938_out1            : std_logic;
  SIGNAL Logical_Operator_out4939_out1            : std_logic;
  SIGNAL Logical_Operator_out4940_out1            : std_logic;
  SIGNAL Logical_Operator_out4941_out1            : std_logic;
  SIGNAL Logical_Operator_out4942_out1            : std_logic;
  SIGNAL Logical_Operator_out4943_out1            : std_logic;
  SIGNAL Logical_Operator_out4944_out1            : std_logic;
  SIGNAL Logical_Operator_out4945_out1            : std_logic;
  SIGNAL Logical_Operator_out4946_out1            : std_logic;
  SIGNAL Logical_Operator_out4947_out1            : std_logic;
  SIGNAL Logical_Operator_out4948_out1            : std_logic;
  SIGNAL Logical_Operator_out4949_out1            : std_logic;
  SIGNAL Logical_Operator_out4950_out1            : std_logic;
  SIGNAL Logical_Operator_out4951_out1            : std_logic;
  SIGNAL Logical_Operator_out4952_out1            : std_logic;
  SIGNAL Logical_Operator_out4953_out1            : std_logic;
  SIGNAL Logical_Operator_out4954_out1            : std_logic;
  SIGNAL Logical_Operator_out4955_out1            : std_logic;
  SIGNAL Logical_Operator_out4956_out1            : std_logic;
  SIGNAL Logical_Operator_out4957_out1            : std_logic;
  SIGNAL Logical_Operator_out4958_out1            : std_logic;
  SIGNAL Logical_Operator_out4959_out1            : std_logic;
  SIGNAL Logical_Operator_out4960_out1            : std_logic;
  SIGNAL Logical_Operator_out4961_out1            : std_logic;
  SIGNAL Logical_Operator_out4962_out1            : std_logic;
  SIGNAL Logical_Operator_out4963_out1            : std_logic;
  SIGNAL Logical_Operator_out4964_out1            : std_logic;
  SIGNAL Logical_Operator_out4965_out1            : std_logic;
  SIGNAL Logical_Operator_out4966_out1            : std_logic;
  SIGNAL Logical_Operator_out4967_out1            : std_logic;
  SIGNAL Logical_Operator_out4968_out1            : std_logic;
  SIGNAL Logical_Operator_out4969_out1            : std_logic;
  SIGNAL Logical_Operator_out4970_out1            : std_logic;
  SIGNAL Logical_Operator_out4971_out1            : std_logic;
  SIGNAL Logical_Operator_out4972_out1            : std_logic;
  SIGNAL Logical_Operator_out4973_out1            : std_logic;
  SIGNAL Logical_Operator_out4974_out1            : std_logic;
  SIGNAL Logical_Operator_out4975_out1            : std_logic;
  SIGNAL Logical_Operator_out4976_out1            : std_logic;
  SIGNAL Logical_Operator_out4977_out1            : std_logic;
  SIGNAL Logical_Operator_out4978_out1            : std_logic;
  SIGNAL Logical_Operator_out4979_out1            : std_logic;
  SIGNAL Logical_Operator_out4980_out1            : std_logic;
  SIGNAL Logical_Operator_out4981_out1            : std_logic;
  SIGNAL Logical_Operator_out4982_out1            : std_logic;
  SIGNAL Logical_Operator_out4983_out1            : std_logic;
  SIGNAL Logical_Operator_out4984_out1            : std_logic;
  SIGNAL Logical_Operator_out4985_out1            : std_logic;
  SIGNAL Logical_Operator_out4986_out1            : std_logic;
  SIGNAL Logical_Operator_out4987_out1            : std_logic;
  SIGNAL Logical_Operator_out4988_out1            : std_logic;
  SIGNAL Logical_Operator_out4989_out1            : std_logic;
  SIGNAL Logical_Operator_out4990_out1            : std_logic;
  SIGNAL Logical_Operator_out4991_out1            : std_logic;
  SIGNAL Logical_Operator_out4992_out1            : std_logic;
  SIGNAL Logical_Operator_out4993_out1            : std_logic;
  SIGNAL Logical_Operator_out4994_out1            : std_logic;
  SIGNAL Logical_Operator_out4995_out1            : std_logic;
  SIGNAL Logical_Operator_out4996_out1            : std_logic;
  SIGNAL Logical_Operator_out4997_out1            : std_logic;
  SIGNAL Logical_Operator_out4998_out1            : std_logic;
  SIGNAL Logical_Operator_out4999_out1            : std_logic;
  SIGNAL Logical_Operator_out5000_out1            : std_logic;
  SIGNAL Logical_Operator_out5001_out1            : std_logic;
  SIGNAL Logical_Operator_out5002_out1            : std_logic;
  SIGNAL Logical_Operator_out5003_out1            : std_logic;
  SIGNAL Logical_Operator_out5004_out1            : std_logic;
  SIGNAL Logical_Operator_out5005_out1            : std_logic;
  SIGNAL Logical_Operator_out5006_out1            : std_logic;
  SIGNAL Logical_Operator_out5007_out1            : std_logic;
  SIGNAL Logical_Operator_out5008_out1            : std_logic;
  SIGNAL Logical_Operator_out5009_out1            : std_logic;
  SIGNAL Logical_Operator_out5010_out1            : std_logic;
  SIGNAL Logical_Operator_out5011_out1            : std_logic;
  SIGNAL Logical_Operator_out5012_out1            : std_logic;
  SIGNAL Logical_Operator_out5013_out1            : std_logic;
  SIGNAL Logical_Operator_out5014_out1            : std_logic;
  SIGNAL Logical_Operator_out5015_out1            : std_logic;
  SIGNAL Logical_Operator_out5016_out1            : std_logic;
  SIGNAL Logical_Operator_out5017_out1            : std_logic;
  SIGNAL Logical_Operator_out5018_out1            : std_logic;
  SIGNAL Logical_Operator_out5019_out1            : std_logic;
  SIGNAL Logical_Operator_out5020_out1            : std_logic;
  SIGNAL Logical_Operator_out5021_out1            : std_logic;
  SIGNAL Logical_Operator_out5022_out1            : std_logic;
  SIGNAL Logical_Operator_out5023_out1            : std_logic;
  SIGNAL Logical_Operator_out5024_out1            : std_logic;
  SIGNAL Logical_Operator_out5025_out1            : std_logic;
  SIGNAL Logical_Operator_out5026_out1            : std_logic;
  SIGNAL Logical_Operator_out5027_out1            : std_logic;
  SIGNAL Logical_Operator_out5028_out1            : std_logic;
  SIGNAL Logical_Operator_out5029_out1            : std_logic;
  SIGNAL Logical_Operator_out5030_out1            : std_logic;
  SIGNAL Logical_Operator_out5031_out1            : std_logic;
  SIGNAL Logical_Operator_out5032_out1            : std_logic;
  SIGNAL Logical_Operator_out5033_out1            : std_logic;
  SIGNAL Logical_Operator_out5034_out1            : std_logic;
  SIGNAL Logical_Operator_out5035_out1            : std_logic;
  SIGNAL Logical_Operator_out5036_out1            : std_logic;
  SIGNAL Logical_Operator_out5037_out1            : std_logic;
  SIGNAL Logical_Operator_out5038_out1            : std_logic;
  SIGNAL Logical_Operator_out5039_out1            : std_logic;
  SIGNAL Logical_Operator_out5040_out1            : std_logic;
  SIGNAL Logical_Operator_out5041_out1            : std_logic;
  SIGNAL Logical_Operator_out5042_out1            : std_logic;
  SIGNAL Logical_Operator_out5043_out1            : std_logic;
  SIGNAL Logical_Operator_out5044_out1            : std_logic;
  SIGNAL Logical_Operator_out5045_out1            : std_logic;
  SIGNAL Logical_Operator_out5046_out1            : std_logic;
  SIGNAL Logical_Operator_out5047_out1            : std_logic;
  SIGNAL Logical_Operator_out5048_out1            : std_logic;
  SIGNAL Logical_Operator_out5049_out1            : std_logic;
  SIGNAL Logical_Operator_out5050_out1            : std_logic;
  SIGNAL Logical_Operator_out5051_out1            : std_logic;
  SIGNAL Logical_Operator_out5052_out1            : std_logic;
  SIGNAL Logical_Operator_out5053_out1            : std_logic;
  SIGNAL Logical_Operator_out5054_out1            : std_logic;
  SIGNAL Logical_Operator_out5055_out1            : std_logic;
  SIGNAL Logical_Operator_out5056_out1            : std_logic;
  SIGNAL Logical_Operator_out5057_out1            : std_logic;
  SIGNAL Logical_Operator_out5058_out1            : std_logic;
  SIGNAL Logical_Operator_out5059_out1            : std_logic;
  SIGNAL Logical_Operator_out5060_out1            : std_logic;
  SIGNAL Logical_Operator_out5061_out1            : std_logic;
  SIGNAL Logical_Operator_out5062_out1            : std_logic;
  SIGNAL Logical_Operator_out5063_out1            : std_logic;
  SIGNAL Logical_Operator_out5064_out1            : std_logic;
  SIGNAL Logical_Operator_out5065_out1            : std_logic;
  SIGNAL Logical_Operator_out5066_out1            : std_logic;
  SIGNAL Logical_Operator_out5067_out1            : std_logic;
  SIGNAL Logical_Operator_out5068_out1            : std_logic;
  SIGNAL Logical_Operator_out5069_out1            : std_logic;
  SIGNAL Logical_Operator_out5070_out1            : std_logic;
  SIGNAL Logical_Operator_out5071_out1            : std_logic;
  SIGNAL Logical_Operator_out5072_out1            : std_logic;
  SIGNAL Logical_Operator_out5073_out1            : std_logic;
  SIGNAL Logical_Operator_out5074_out1            : std_logic;
  SIGNAL Logical_Operator_out5075_out1            : std_logic;
  SIGNAL Logical_Operator_out5076_out1            : std_logic;
  SIGNAL Logical_Operator_out5077_out1            : std_logic;
  SIGNAL Logical_Operator_out5078_out1            : std_logic;
  SIGNAL Logical_Operator_out5079_out1            : std_logic;
  SIGNAL Logical_Operator_out5080_out1            : std_logic;
  SIGNAL Logical_Operator_out5081_out1            : std_logic;
  SIGNAL Logical_Operator_out5082_out1            : std_logic;
  SIGNAL Logical_Operator_out5083_out1            : std_logic;
  SIGNAL Logical_Operator_out5084_out1            : std_logic;
  SIGNAL Logical_Operator_out5085_out1            : std_logic;
  SIGNAL Logical_Operator_out5086_out1            : std_logic;
  SIGNAL Logical_Operator_out5087_out1            : std_logic;
  SIGNAL Logical_Operator_out5088_out1            : std_logic;
  SIGNAL Logical_Operator_out5089_out1            : std_logic;
  SIGNAL Logical_Operator_out5090_out1            : std_logic;
  SIGNAL Logical_Operator_out5091_out1            : std_logic;
  SIGNAL Logical_Operator_out5092_out1            : std_logic;
  SIGNAL Logical_Operator_out5093_out1            : std_logic;
  SIGNAL Logical_Operator_out5094_out1            : std_logic;
  SIGNAL Logical_Operator_out5095_out1            : std_logic;
  SIGNAL Logical_Operator_out5096_out1            : std_logic;
  SIGNAL Logical_Operator_out5097_out1            : std_logic;
  SIGNAL Logical_Operator_out5098_out1            : std_logic;
  SIGNAL Logical_Operator_out5099_out1            : std_logic;
  SIGNAL Logical_Operator_out5100_out1            : std_logic;
  SIGNAL Logical_Operator_out5101_out1            : std_logic;
  SIGNAL Logical_Operator_out5102_out1            : std_logic;
  SIGNAL Logical_Operator_out5103_out1            : std_logic;
  SIGNAL Logical_Operator_out5104_out1            : std_logic;
  SIGNAL Logical_Operator_out5105_out1            : std_logic;
  SIGNAL Logical_Operator_out5106_out1            : std_logic;
  SIGNAL Logical_Operator_out5107_out1            : std_logic;
  SIGNAL Logical_Operator_out5108_out1            : std_logic;
  SIGNAL Logical_Operator_out5109_out1            : std_logic;
  SIGNAL Logical_Operator_out5110_out1            : std_logic;
  SIGNAL Logical_Operator_out5111_out1            : std_logic;
  SIGNAL Logical_Operator_out5112_out1            : std_logic;
  SIGNAL Logical_Operator_out5113_out1            : std_logic;
  SIGNAL Logical_Operator_out5114_out1            : std_logic;
  SIGNAL Logical_Operator_out5115_out1            : std_logic;
  SIGNAL Logical_Operator_out5116_out1            : std_logic;
  SIGNAL Logical_Operator_out5117_out1            : std_logic;
  SIGNAL Logical_Operator_out5118_out1            : std_logic;
  SIGNAL Logical_Operator_out5119_out1            : std_logic;
  SIGNAL Logical_Operator_out5120_out1            : std_logic;

BEGIN

  Logical_Operator_out1_out1 <= in1 XOR in2;

  Logical_Operator_out2_out1 <= in3 XOR in4;

  Logical_Operator_out3_out1 <= in5 XOR in6;

  Logical_Operator_out4_out1 <= in7 XOR in8;

  Logical_Operator_out5_out1 <= in9 XOR in10;

  Logical_Operator_out6_out1 <= in11 XOR in12;

  Logical_Operator_out7_out1 <= in13 XOR in14;

  Logical_Operator_out8_out1 <= in15 XOR in16;

  Logical_Operator_out9_out1 <= in17 XOR in18;

  Logical_Operator_out10_out1 <= in19 XOR in20;

  Logical_Operator_out11_out1 <= in21 XOR in22;

  Logical_Operator_out12_out1 <= in23 XOR in24;

  Logical_Operator_out13_out1 <= in25 XOR in26;

  Logical_Operator_out14_out1 <= in27 XOR in28;

  Logical_Operator_out15_out1 <= in29 XOR in30;

  Logical_Operator_out16_out1 <= in31 XOR in32;

  Logical_Operator_out17_out1 <= in33 XOR in34;

  Logical_Operator_out18_out1 <= in35 XOR in36;

  Logical_Operator_out19_out1 <= in37 XOR in38;

  Logical_Operator_out20_out1 <= in39 XOR in40;

  Logical_Operator_out21_out1 <= in41 XOR in42;

  Logical_Operator_out22_out1 <= in43 XOR in44;

  Logical_Operator_out23_out1 <= in45 XOR in46;

  Logical_Operator_out24_out1 <= in47 XOR in48;

  Logical_Operator_out25_out1 <= in49 XOR in50;

  Logical_Operator_out26_out1 <= in51 XOR in52;

  Logical_Operator_out27_out1 <= in53 XOR in54;

  Logical_Operator_out28_out1 <= in55 XOR in56;

  Logical_Operator_out29_out1 <= in57 XOR in58;

  Logical_Operator_out30_out1 <= in59 XOR in60;

  Logical_Operator_out31_out1 <= in61 XOR in62;

  Logical_Operator_out32_out1 <= in63 XOR in64;

  Logical_Operator_out33_out1 <= in65 XOR in66;

  Logical_Operator_out34_out1 <= in67 XOR in68;

  Logical_Operator_out35_out1 <= in69 XOR in70;

  Logical_Operator_out36_out1 <= in71 XOR in72;

  Logical_Operator_out37_out1 <= in73 XOR in74;

  Logical_Operator_out38_out1 <= in75 XOR in76;

  Logical_Operator_out39_out1 <= in77 XOR in78;

  Logical_Operator_out40_out1 <= in79 XOR in80;

  Logical_Operator_out41_out1 <= in81 XOR in82;

  Logical_Operator_out42_out1 <= in83 XOR in84;

  Logical_Operator_out43_out1 <= in85 XOR in86;

  Logical_Operator_out44_out1 <= in87 XOR in88;

  Logical_Operator_out45_out1 <= in89 XOR in90;

  Logical_Operator_out46_out1 <= in91 XOR in92;

  Logical_Operator_out47_out1 <= in93 XOR in94;

  Logical_Operator_out48_out1 <= in95 XOR in96;

  Logical_Operator_out49_out1 <= in97 XOR in98;

  Logical_Operator_out50_out1 <= in99 XOR in100;

  Logical_Operator_out51_out1 <= in101 XOR in102;

  Logical_Operator_out52_out1 <= in103 XOR in104;

  Logical_Operator_out53_out1 <= in105 XOR in106;

  Logical_Operator_out54_out1 <= in107 XOR in108;

  Logical_Operator_out55_out1 <= in109 XOR in110;

  Logical_Operator_out56_out1 <= in111 XOR in112;

  Logical_Operator_out57_out1 <= in113 XOR in114;

  Logical_Operator_out58_out1 <= in115 XOR in116;

  Logical_Operator_out59_out1 <= in117 XOR in118;

  Logical_Operator_out60_out1 <= in119 XOR in120;

  Logical_Operator_out61_out1 <= in121 XOR in122;

  Logical_Operator_out62_out1 <= in123 XOR in124;

  Logical_Operator_out63_out1 <= in125 XOR in126;

  Logical_Operator_out64_out1 <= in127 XOR in128;

  Logical_Operator_out65_out1 <= in129 XOR in130;

  Logical_Operator_out66_out1 <= in131 XOR in132;

  Logical_Operator_out67_out1 <= in133 XOR in134;

  Logical_Operator_out68_out1 <= in135 XOR in136;

  Logical_Operator_out69_out1 <= in137 XOR in138;

  Logical_Operator_out70_out1 <= in139 XOR in140;

  Logical_Operator_out71_out1 <= in141 XOR in142;

  Logical_Operator_out72_out1 <= in143 XOR in144;

  Logical_Operator_out73_out1 <= in145 XOR in146;

  Logical_Operator_out74_out1 <= in147 XOR in148;

  Logical_Operator_out75_out1 <= in149 XOR in150;

  Logical_Operator_out76_out1 <= in151 XOR in152;

  Logical_Operator_out77_out1 <= in153 XOR in154;

  Logical_Operator_out78_out1 <= in155 XOR in156;

  Logical_Operator_out79_out1 <= in157 XOR in158;

  Logical_Operator_out80_out1 <= in159 XOR in160;

  Logical_Operator_out81_out1 <= in161 XOR in162;

  Logical_Operator_out82_out1 <= in163 XOR in164;

  Logical_Operator_out83_out1 <= in165 XOR in166;

  Logical_Operator_out84_out1 <= in167 XOR in168;

  Logical_Operator_out85_out1 <= in169 XOR in170;

  Logical_Operator_out86_out1 <= in171 XOR in172;

  Logical_Operator_out87_out1 <= in173 XOR in174;

  Logical_Operator_out88_out1 <= in175 XOR in176;

  Logical_Operator_out89_out1 <= in177 XOR in178;

  Logical_Operator_out90_out1 <= in179 XOR in180;

  Logical_Operator_out91_out1 <= in181 XOR in182;

  Logical_Operator_out92_out1 <= in183 XOR in184;

  Logical_Operator_out93_out1 <= in185 XOR in186;

  Logical_Operator_out94_out1 <= in187 XOR in188;

  Logical_Operator_out95_out1 <= in189 XOR in190;

  Logical_Operator_out96_out1 <= in191 XOR in192;

  Logical_Operator_out97_out1 <= in193 XOR in194;

  Logical_Operator_out98_out1 <= in195 XOR in196;

  Logical_Operator_out99_out1 <= in197 XOR in198;

  Logical_Operator_out100_out1 <= in199 XOR in200;

  Logical_Operator_out101_out1 <= in201 XOR in202;

  Logical_Operator_out102_out1 <= in203 XOR in204;

  Logical_Operator_out103_out1 <= in205 XOR in206;

  Logical_Operator_out104_out1 <= in207 XOR in208;

  Logical_Operator_out105_out1 <= in209 XOR in210;

  Logical_Operator_out106_out1 <= in211 XOR in212;

  Logical_Operator_out107_out1 <= in213 XOR in214;

  Logical_Operator_out108_out1 <= in215 XOR in216;

  Logical_Operator_out109_out1 <= in217 XOR in218;

  Logical_Operator_out110_out1 <= in219 XOR in220;

  Logical_Operator_out111_out1 <= in221 XOR in222;

  Logical_Operator_out112_out1 <= in223 XOR in224;

  Logical_Operator_out113_out1 <= in225 XOR in226;

  Logical_Operator_out114_out1 <= in227 XOR in228;

  Logical_Operator_out115_out1 <= in229 XOR in230;

  Logical_Operator_out116_out1 <= in231 XOR in232;

  Logical_Operator_out117_out1 <= in233 XOR in234;

  Logical_Operator_out118_out1 <= in235 XOR in236;

  Logical_Operator_out119_out1 <= in237 XOR in238;

  Logical_Operator_out120_out1 <= in239 XOR in240;

  Logical_Operator_out121_out1 <= in241 XOR in242;

  Logical_Operator_out122_out1 <= in243 XOR in244;

  Logical_Operator_out123_out1 <= in245 XOR in246;

  Logical_Operator_out124_out1 <= in247 XOR in248;

  Logical_Operator_out125_out1 <= in249 XOR in250;

  Logical_Operator_out126_out1 <= in251 XOR in252;

  Logical_Operator_out127_out1 <= in253 XOR in254;

  Logical_Operator_out128_out1 <= in255 XOR in256;

  Logical_Operator_out129_out1 <= in257 XOR in258;

  Logical_Operator_out130_out1 <= in259 XOR in260;

  Logical_Operator_out131_out1 <= in261 XOR in262;

  Logical_Operator_out132_out1 <= in263 XOR in264;

  Logical_Operator_out133_out1 <= in265 XOR in266;

  Logical_Operator_out134_out1 <= in267 XOR in268;

  Logical_Operator_out135_out1 <= in269 XOR in270;

  Logical_Operator_out136_out1 <= in271 XOR in272;

  Logical_Operator_out137_out1 <= in273 XOR in274;

  Logical_Operator_out138_out1 <= in275 XOR in276;

  Logical_Operator_out139_out1 <= in277 XOR in278;

  Logical_Operator_out140_out1 <= in279 XOR in280;

  Logical_Operator_out141_out1 <= in281 XOR in282;

  Logical_Operator_out142_out1 <= in283 XOR in284;

  Logical_Operator_out143_out1 <= in285 XOR in286;

  Logical_Operator_out144_out1 <= in287 XOR in288;

  Logical_Operator_out145_out1 <= in289 XOR in290;

  Logical_Operator_out146_out1 <= in291 XOR in292;

  Logical_Operator_out147_out1 <= in293 XOR in294;

  Logical_Operator_out148_out1 <= in295 XOR in296;

  Logical_Operator_out149_out1 <= in297 XOR in298;

  Logical_Operator_out150_out1 <= in299 XOR in300;

  Logical_Operator_out151_out1 <= in301 XOR in302;

  Logical_Operator_out152_out1 <= in303 XOR in304;

  Logical_Operator_out153_out1 <= in305 XOR in306;

  Logical_Operator_out154_out1 <= in307 XOR in308;

  Logical_Operator_out155_out1 <= in309 XOR in310;

  Logical_Operator_out156_out1 <= in311 XOR in312;

  Logical_Operator_out157_out1 <= in313 XOR in314;

  Logical_Operator_out158_out1 <= in315 XOR in316;

  Logical_Operator_out159_out1 <= in317 XOR in318;

  Logical_Operator_out160_out1 <= in319 XOR in320;

  Logical_Operator_out161_out1 <= in321 XOR in322;

  Logical_Operator_out162_out1 <= in323 XOR in324;

  Logical_Operator_out163_out1 <= in325 XOR in326;

  Logical_Operator_out164_out1 <= in327 XOR in328;

  Logical_Operator_out165_out1 <= in329 XOR in330;

  Logical_Operator_out166_out1 <= in331 XOR in332;

  Logical_Operator_out167_out1 <= in333 XOR in334;

  Logical_Operator_out168_out1 <= in335 XOR in336;

  Logical_Operator_out169_out1 <= in337 XOR in338;

  Logical_Operator_out170_out1 <= in339 XOR in340;

  Logical_Operator_out171_out1 <= in341 XOR in342;

  Logical_Operator_out172_out1 <= in343 XOR in344;

  Logical_Operator_out173_out1 <= in345 XOR in346;

  Logical_Operator_out174_out1 <= in347 XOR in348;

  Logical_Operator_out175_out1 <= in349 XOR in350;

  Logical_Operator_out176_out1 <= in351 XOR in352;

  Logical_Operator_out177_out1 <= in353 XOR in354;

  Logical_Operator_out178_out1 <= in355 XOR in356;

  Logical_Operator_out179_out1 <= in357 XOR in358;

  Logical_Operator_out180_out1 <= in359 XOR in360;

  Logical_Operator_out181_out1 <= in361 XOR in362;

  Logical_Operator_out182_out1 <= in363 XOR in364;

  Logical_Operator_out183_out1 <= in365 XOR in366;

  Logical_Operator_out184_out1 <= in367 XOR in368;

  Logical_Operator_out185_out1 <= in369 XOR in370;

  Logical_Operator_out186_out1 <= in371 XOR in372;

  Logical_Operator_out187_out1 <= in373 XOR in374;

  Logical_Operator_out188_out1 <= in375 XOR in376;

  Logical_Operator_out189_out1 <= in377 XOR in378;

  Logical_Operator_out190_out1 <= in379 XOR in380;

  Logical_Operator_out191_out1 <= in381 XOR in382;

  Logical_Operator_out192_out1 <= in383 XOR in384;

  Logical_Operator_out193_out1 <= in385 XOR in386;

  Logical_Operator_out194_out1 <= in387 XOR in388;

  Logical_Operator_out195_out1 <= in389 XOR in390;

  Logical_Operator_out196_out1 <= in391 XOR in392;

  Logical_Operator_out197_out1 <= in393 XOR in394;

  Logical_Operator_out198_out1 <= in395 XOR in396;

  Logical_Operator_out199_out1 <= in397 XOR in398;

  Logical_Operator_out200_out1 <= in399 XOR in400;

  Logical_Operator_out201_out1 <= in401 XOR in402;

  Logical_Operator_out202_out1 <= in403 XOR in404;

  Logical_Operator_out203_out1 <= in405 XOR in406;

  Logical_Operator_out204_out1 <= in407 XOR in408;

  Logical_Operator_out205_out1 <= in409 XOR in410;

  Logical_Operator_out206_out1 <= in411 XOR in412;

  Logical_Operator_out207_out1 <= in413 XOR in414;

  Logical_Operator_out208_out1 <= in415 XOR in416;

  Logical_Operator_out209_out1 <= in417 XOR in418;

  Logical_Operator_out210_out1 <= in419 XOR in420;

  Logical_Operator_out211_out1 <= in421 XOR in422;

  Logical_Operator_out212_out1 <= in423 XOR in424;

  Logical_Operator_out213_out1 <= in425 XOR in426;

  Logical_Operator_out214_out1 <= in427 XOR in428;

  Logical_Operator_out215_out1 <= in429 XOR in430;

  Logical_Operator_out216_out1 <= in431 XOR in432;

  Logical_Operator_out217_out1 <= in433 XOR in434;

  Logical_Operator_out218_out1 <= in435 XOR in436;

  Logical_Operator_out219_out1 <= in437 XOR in438;

  Logical_Operator_out220_out1 <= in439 XOR in440;

  Logical_Operator_out221_out1 <= in441 XOR in442;

  Logical_Operator_out222_out1 <= in443 XOR in444;

  Logical_Operator_out223_out1 <= in445 XOR in446;

  Logical_Operator_out224_out1 <= in447 XOR in448;

  Logical_Operator_out225_out1 <= in449 XOR in450;

  Logical_Operator_out226_out1 <= in451 XOR in452;

  Logical_Operator_out227_out1 <= in453 XOR in454;

  Logical_Operator_out228_out1 <= in455 XOR in456;

  Logical_Operator_out229_out1 <= in457 XOR in458;

  Logical_Operator_out230_out1 <= in459 XOR in460;

  Logical_Operator_out231_out1 <= in461 XOR in462;

  Logical_Operator_out232_out1 <= in463 XOR in464;

  Logical_Operator_out233_out1 <= in465 XOR in466;

  Logical_Operator_out234_out1 <= in467 XOR in468;

  Logical_Operator_out235_out1 <= in469 XOR in470;

  Logical_Operator_out236_out1 <= in471 XOR in472;

  Logical_Operator_out237_out1 <= in473 XOR in474;

  Logical_Operator_out238_out1 <= in475 XOR in476;

  Logical_Operator_out239_out1 <= in477 XOR in478;

  Logical_Operator_out240_out1 <= in479 XOR in480;

  Logical_Operator_out241_out1 <= in481 XOR in482;

  Logical_Operator_out242_out1 <= in483 XOR in484;

  Logical_Operator_out243_out1 <= in485 XOR in486;

  Logical_Operator_out244_out1 <= in487 XOR in488;

  Logical_Operator_out245_out1 <= in489 XOR in490;

  Logical_Operator_out246_out1 <= in491 XOR in492;

  Logical_Operator_out247_out1 <= in493 XOR in494;

  Logical_Operator_out248_out1 <= in495 XOR in496;

  Logical_Operator_out249_out1 <= in497 XOR in498;

  Logical_Operator_out250_out1 <= in499 XOR in500;

  Logical_Operator_out251_out1 <= in501 XOR in502;

  Logical_Operator_out252_out1 <= in503 XOR in504;

  Logical_Operator_out253_out1 <= in505 XOR in506;

  Logical_Operator_out254_out1 <= in507 XOR in508;

  Logical_Operator_out255_out1 <= in509 XOR in510;

  Logical_Operator_out256_out1 <= in511 XOR in512;

  Logical_Operator_out257_out1 <= in513 XOR in514;

  Logical_Operator_out258_out1 <= in515 XOR in516;

  Logical_Operator_out259_out1 <= in517 XOR in518;

  Logical_Operator_out260_out1 <= in519 XOR in520;

  Logical_Operator_out261_out1 <= in521 XOR in522;

  Logical_Operator_out262_out1 <= in523 XOR in524;

  Logical_Operator_out263_out1 <= in525 XOR in526;

  Logical_Operator_out264_out1 <= in527 XOR in528;

  Logical_Operator_out265_out1 <= in529 XOR in530;

  Logical_Operator_out266_out1 <= in531 XOR in532;

  Logical_Operator_out267_out1 <= in533 XOR in534;

  Logical_Operator_out268_out1 <= in535 XOR in536;

  Logical_Operator_out269_out1 <= in537 XOR in538;

  Logical_Operator_out270_out1 <= in539 XOR in540;

  Logical_Operator_out271_out1 <= in541 XOR in542;

  Logical_Operator_out272_out1 <= in543 XOR in544;

  Logical_Operator_out273_out1 <= in545 XOR in546;

  Logical_Operator_out274_out1 <= in547 XOR in548;

  Logical_Operator_out275_out1 <= in549 XOR in550;

  Logical_Operator_out276_out1 <= in551 XOR in552;

  Logical_Operator_out277_out1 <= in553 XOR in554;

  Logical_Operator_out278_out1 <= in555 XOR in556;

  Logical_Operator_out279_out1 <= in557 XOR in558;

  Logical_Operator_out280_out1 <= in559 XOR in560;

  Logical_Operator_out281_out1 <= in561 XOR in562;

  Logical_Operator_out282_out1 <= in563 XOR in564;

  Logical_Operator_out283_out1 <= in565 XOR in566;

  Logical_Operator_out284_out1 <= in567 XOR in568;

  Logical_Operator_out285_out1 <= in569 XOR in570;

  Logical_Operator_out286_out1 <= in571 XOR in572;

  Logical_Operator_out287_out1 <= in573 XOR in574;

  Logical_Operator_out288_out1 <= in575 XOR in576;

  Logical_Operator_out289_out1 <= in577 XOR in578;

  Logical_Operator_out290_out1 <= in579 XOR in580;

  Logical_Operator_out291_out1 <= in581 XOR in582;

  Logical_Operator_out292_out1 <= in583 XOR in584;

  Logical_Operator_out293_out1 <= in585 XOR in586;

  Logical_Operator_out294_out1 <= in587 XOR in588;

  Logical_Operator_out295_out1 <= in589 XOR in590;

  Logical_Operator_out296_out1 <= in591 XOR in592;

  Logical_Operator_out297_out1 <= in593 XOR in594;

  Logical_Operator_out298_out1 <= in595 XOR in596;

  Logical_Operator_out299_out1 <= in597 XOR in598;

  Logical_Operator_out300_out1 <= in599 XOR in600;

  Logical_Operator_out301_out1 <= in601 XOR in602;

  Logical_Operator_out302_out1 <= in603 XOR in604;

  Logical_Operator_out303_out1 <= in605 XOR in606;

  Logical_Operator_out304_out1 <= in607 XOR in608;

  Logical_Operator_out305_out1 <= in609 XOR in610;

  Logical_Operator_out306_out1 <= in611 XOR in612;

  Logical_Operator_out307_out1 <= in613 XOR in614;

  Logical_Operator_out308_out1 <= in615 XOR in616;

  Logical_Operator_out309_out1 <= in617 XOR in618;

  Logical_Operator_out310_out1 <= in619 XOR in620;

  Logical_Operator_out311_out1 <= in621 XOR in622;

  Logical_Operator_out312_out1 <= in623 XOR in624;

  Logical_Operator_out313_out1 <= in625 XOR in626;

  Logical_Operator_out314_out1 <= in627 XOR in628;

  Logical_Operator_out315_out1 <= in629 XOR in630;

  Logical_Operator_out316_out1 <= in631 XOR in632;

  Logical_Operator_out317_out1 <= in633 XOR in634;

  Logical_Operator_out318_out1 <= in635 XOR in636;

  Logical_Operator_out319_out1 <= in637 XOR in638;

  Logical_Operator_out320_out1 <= in639 XOR in640;

  Logical_Operator_out321_out1 <= in641 XOR in642;

  Logical_Operator_out322_out1 <= in643 XOR in644;

  Logical_Operator_out323_out1 <= in645 XOR in646;

  Logical_Operator_out324_out1 <= in647 XOR in648;

  Logical_Operator_out325_out1 <= in649 XOR in650;

  Logical_Operator_out326_out1 <= in651 XOR in652;

  Logical_Operator_out327_out1 <= in653 XOR in654;

  Logical_Operator_out328_out1 <= in655 XOR in656;

  Logical_Operator_out329_out1 <= in657 XOR in658;

  Logical_Operator_out330_out1 <= in659 XOR in660;

  Logical_Operator_out331_out1 <= in661 XOR in662;

  Logical_Operator_out332_out1 <= in663 XOR in664;

  Logical_Operator_out333_out1 <= in665 XOR in666;

  Logical_Operator_out334_out1 <= in667 XOR in668;

  Logical_Operator_out335_out1 <= in669 XOR in670;

  Logical_Operator_out336_out1 <= in671 XOR in672;

  Logical_Operator_out337_out1 <= in673 XOR in674;

  Logical_Operator_out338_out1 <= in675 XOR in676;

  Logical_Operator_out339_out1 <= in677 XOR in678;

  Logical_Operator_out340_out1 <= in679 XOR in680;

  Logical_Operator_out341_out1 <= in681 XOR in682;

  Logical_Operator_out342_out1 <= in683 XOR in684;

  Logical_Operator_out343_out1 <= in685 XOR in686;

  Logical_Operator_out344_out1 <= in687 XOR in688;

  Logical_Operator_out345_out1 <= in689 XOR in690;

  Logical_Operator_out346_out1 <= in691 XOR in692;

  Logical_Operator_out347_out1 <= in693 XOR in694;

  Logical_Operator_out348_out1 <= in695 XOR in696;

  Logical_Operator_out349_out1 <= in697 XOR in698;

  Logical_Operator_out350_out1 <= in699 XOR in700;

  Logical_Operator_out351_out1 <= in701 XOR in702;

  Logical_Operator_out352_out1 <= in703 XOR in704;

  Logical_Operator_out353_out1 <= in705 XOR in706;

  Logical_Operator_out354_out1 <= in707 XOR in708;

  Logical_Operator_out355_out1 <= in709 XOR in710;

  Logical_Operator_out356_out1 <= in711 XOR in712;

  Logical_Operator_out357_out1 <= in713 XOR in714;

  Logical_Operator_out358_out1 <= in715 XOR in716;

  Logical_Operator_out359_out1 <= in717 XOR in718;

  Logical_Operator_out360_out1 <= in719 XOR in720;

  Logical_Operator_out361_out1 <= in721 XOR in722;

  Logical_Operator_out362_out1 <= in723 XOR in724;

  Logical_Operator_out363_out1 <= in725 XOR in726;

  Logical_Operator_out364_out1 <= in727 XOR in728;

  Logical_Operator_out365_out1 <= in729 XOR in730;

  Logical_Operator_out366_out1 <= in731 XOR in732;

  Logical_Operator_out367_out1 <= in733 XOR in734;

  Logical_Operator_out368_out1 <= in735 XOR in736;

  Logical_Operator_out369_out1 <= in737 XOR in738;

  Logical_Operator_out370_out1 <= in739 XOR in740;

  Logical_Operator_out371_out1 <= in741 XOR in742;

  Logical_Operator_out372_out1 <= in743 XOR in744;

  Logical_Operator_out373_out1 <= in745 XOR in746;

  Logical_Operator_out374_out1 <= in747 XOR in748;

  Logical_Operator_out375_out1 <= in749 XOR in750;

  Logical_Operator_out376_out1 <= in751 XOR in752;

  Logical_Operator_out377_out1 <= in753 XOR in754;

  Logical_Operator_out378_out1 <= in755 XOR in756;

  Logical_Operator_out379_out1 <= in757 XOR in758;

  Logical_Operator_out380_out1 <= in759 XOR in760;

  Logical_Operator_out381_out1 <= in761 XOR in762;

  Logical_Operator_out382_out1 <= in763 XOR in764;

  Logical_Operator_out383_out1 <= in765 XOR in766;

  Logical_Operator_out384_out1 <= in767 XOR in768;

  Logical_Operator_out385_out1 <= in769 XOR in770;

  Logical_Operator_out386_out1 <= in771 XOR in772;

  Logical_Operator_out387_out1 <= in773 XOR in774;

  Logical_Operator_out388_out1 <= in775 XOR in776;

  Logical_Operator_out389_out1 <= in777 XOR in778;

  Logical_Operator_out390_out1 <= in779 XOR in780;

  Logical_Operator_out391_out1 <= in781 XOR in782;

  Logical_Operator_out392_out1 <= in783 XOR in784;

  Logical_Operator_out393_out1 <= in785 XOR in786;

  Logical_Operator_out394_out1 <= in787 XOR in788;

  Logical_Operator_out395_out1 <= in789 XOR in790;

  Logical_Operator_out396_out1 <= in791 XOR in792;

  Logical_Operator_out397_out1 <= in793 XOR in794;

  Logical_Operator_out398_out1 <= in795 XOR in796;

  Logical_Operator_out399_out1 <= in797 XOR in798;

  Logical_Operator_out400_out1 <= in799 XOR in800;

  Logical_Operator_out401_out1 <= in801 XOR in802;

  Logical_Operator_out402_out1 <= in803 XOR in804;

  Logical_Operator_out403_out1 <= in805 XOR in806;

  Logical_Operator_out404_out1 <= in807 XOR in808;

  Logical_Operator_out405_out1 <= in809 XOR in810;

  Logical_Operator_out406_out1 <= in811 XOR in812;

  Logical_Operator_out407_out1 <= in813 XOR in814;

  Logical_Operator_out408_out1 <= in815 XOR in816;

  Logical_Operator_out409_out1 <= in817 XOR in818;

  Logical_Operator_out410_out1 <= in819 XOR in820;

  Logical_Operator_out411_out1 <= in821 XOR in822;

  Logical_Operator_out412_out1 <= in823 XOR in824;

  Logical_Operator_out413_out1 <= in825 XOR in826;

  Logical_Operator_out414_out1 <= in827 XOR in828;

  Logical_Operator_out415_out1 <= in829 XOR in830;

  Logical_Operator_out416_out1 <= in831 XOR in832;

  Logical_Operator_out417_out1 <= in833 XOR in834;

  Logical_Operator_out418_out1 <= in835 XOR in836;

  Logical_Operator_out419_out1 <= in837 XOR in838;

  Logical_Operator_out420_out1 <= in839 XOR in840;

  Logical_Operator_out421_out1 <= in841 XOR in842;

  Logical_Operator_out422_out1 <= in843 XOR in844;

  Logical_Operator_out423_out1 <= in845 XOR in846;

  Logical_Operator_out424_out1 <= in847 XOR in848;

  Logical_Operator_out425_out1 <= in849 XOR in850;

  Logical_Operator_out426_out1 <= in851 XOR in852;

  Logical_Operator_out427_out1 <= in853 XOR in854;

  Logical_Operator_out428_out1 <= in855 XOR in856;

  Logical_Operator_out429_out1 <= in857 XOR in858;

  Logical_Operator_out430_out1 <= in859 XOR in860;

  Logical_Operator_out431_out1 <= in861 XOR in862;

  Logical_Operator_out432_out1 <= in863 XOR in864;

  Logical_Operator_out433_out1 <= in865 XOR in866;

  Logical_Operator_out434_out1 <= in867 XOR in868;

  Logical_Operator_out435_out1 <= in869 XOR in870;

  Logical_Operator_out436_out1 <= in871 XOR in872;

  Logical_Operator_out437_out1 <= in873 XOR in874;

  Logical_Operator_out438_out1 <= in875 XOR in876;

  Logical_Operator_out439_out1 <= in877 XOR in878;

  Logical_Operator_out440_out1 <= in879 XOR in880;

  Logical_Operator_out441_out1 <= in881 XOR in882;

  Logical_Operator_out442_out1 <= in883 XOR in884;

  Logical_Operator_out443_out1 <= in885 XOR in886;

  Logical_Operator_out444_out1 <= in887 XOR in888;

  Logical_Operator_out445_out1 <= in889 XOR in890;

  Logical_Operator_out446_out1 <= in891 XOR in892;

  Logical_Operator_out447_out1 <= in893 XOR in894;

  Logical_Operator_out448_out1 <= in895 XOR in896;

  Logical_Operator_out449_out1 <= in897 XOR in898;

  Logical_Operator_out450_out1 <= in899 XOR in900;

  Logical_Operator_out451_out1 <= in901 XOR in902;

  Logical_Operator_out452_out1 <= in903 XOR in904;

  Logical_Operator_out453_out1 <= in905 XOR in906;

  Logical_Operator_out454_out1 <= in907 XOR in908;

  Logical_Operator_out455_out1 <= in909 XOR in910;

  Logical_Operator_out456_out1 <= in911 XOR in912;

  Logical_Operator_out457_out1 <= in913 XOR in914;

  Logical_Operator_out458_out1 <= in915 XOR in916;

  Logical_Operator_out459_out1 <= in917 XOR in918;

  Logical_Operator_out460_out1 <= in919 XOR in920;

  Logical_Operator_out461_out1 <= in921 XOR in922;

  Logical_Operator_out462_out1 <= in923 XOR in924;

  Logical_Operator_out463_out1 <= in925 XOR in926;

  Logical_Operator_out464_out1 <= in927 XOR in928;

  Logical_Operator_out465_out1 <= in929 XOR in930;

  Logical_Operator_out466_out1 <= in931 XOR in932;

  Logical_Operator_out467_out1 <= in933 XOR in934;

  Logical_Operator_out468_out1 <= in935 XOR in936;

  Logical_Operator_out469_out1 <= in937 XOR in938;

  Logical_Operator_out470_out1 <= in939 XOR in940;

  Logical_Operator_out471_out1 <= in941 XOR in942;

  Logical_Operator_out472_out1 <= in943 XOR in944;

  Logical_Operator_out473_out1 <= in945 XOR in946;

  Logical_Operator_out474_out1 <= in947 XOR in948;

  Logical_Operator_out475_out1 <= in949 XOR in950;

  Logical_Operator_out476_out1 <= in951 XOR in952;

  Logical_Operator_out477_out1 <= in953 XOR in954;

  Logical_Operator_out478_out1 <= in955 XOR in956;

  Logical_Operator_out479_out1 <= in957 XOR in958;

  Logical_Operator_out480_out1 <= in959 XOR in960;

  Logical_Operator_out481_out1 <= in961 XOR in962;

  Logical_Operator_out482_out1 <= in963 XOR in964;

  Logical_Operator_out483_out1 <= in965 XOR in966;

  Logical_Operator_out484_out1 <= in967 XOR in968;

  Logical_Operator_out485_out1 <= in969 XOR in970;

  Logical_Operator_out486_out1 <= in971 XOR in972;

  Logical_Operator_out487_out1 <= in973 XOR in974;

  Logical_Operator_out488_out1 <= in975 XOR in976;

  Logical_Operator_out489_out1 <= in977 XOR in978;

  Logical_Operator_out490_out1 <= in979 XOR in980;

  Logical_Operator_out491_out1 <= in981 XOR in982;

  Logical_Operator_out492_out1 <= in983 XOR in984;

  Logical_Operator_out493_out1 <= in985 XOR in986;

  Logical_Operator_out494_out1 <= in987 XOR in988;

  Logical_Operator_out495_out1 <= in989 XOR in990;

  Logical_Operator_out496_out1 <= in991 XOR in992;

  Logical_Operator_out497_out1 <= in993 XOR in994;

  Logical_Operator_out498_out1 <= in995 XOR in996;

  Logical_Operator_out499_out1 <= in997 XOR in998;

  Logical_Operator_out500_out1 <= in999 XOR in1000;

  Logical_Operator_out501_out1 <= in1001 XOR in1002;

  Logical_Operator_out502_out1 <= in1003 XOR in1004;

  Logical_Operator_out503_out1 <= in1005 XOR in1006;

  Logical_Operator_out504_out1 <= in1007 XOR in1008;

  Logical_Operator_out505_out1 <= in1009 XOR in1010;

  Logical_Operator_out506_out1 <= in1011 XOR in1012;

  Logical_Operator_out507_out1 <= in1013 XOR in1014;

  Logical_Operator_out508_out1 <= in1015 XOR in1016;

  Logical_Operator_out509_out1 <= in1017 XOR in1018;

  Logical_Operator_out510_out1 <= in1019 XOR in1020;

  Logical_Operator_out511_out1 <= in1021 XOR in1022;

  Logical_Operator_out512_out1 <= in1023 XOR in1024;

  Logical_Operator_out513_out1 <= Logical_Operator_out1_out1 XOR Logical_Operator_out2_out1;

  Logical_Operator_out514_out1 <= in2 XOR in4;

  Logical_Operator_out515_out1 <= Logical_Operator_out3_out1 XOR Logical_Operator_out4_out1;

  Logical_Operator_out516_out1 <= in6 XOR in8;

  Logical_Operator_out517_out1 <= Logical_Operator_out5_out1 XOR Logical_Operator_out6_out1;

  Logical_Operator_out518_out1 <= in10 XOR in12;

  Logical_Operator_out519_out1 <= Logical_Operator_out7_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out520_out1 <= in14 XOR in16;

  Logical_Operator_out521_out1 <= Logical_Operator_out9_out1 XOR Logical_Operator_out10_out1;

  Logical_Operator_out522_out1 <= in18 XOR in20;

  Logical_Operator_out523_out1 <= Logical_Operator_out11_out1 XOR Logical_Operator_out12_out1;

  Logical_Operator_out524_out1 <= in22 XOR in24;

  Logical_Operator_out525_out1 <= Logical_Operator_out13_out1 XOR Logical_Operator_out14_out1;

  Logical_Operator_out526_out1 <= in26 XOR in28;

  Logical_Operator_out527_out1 <= Logical_Operator_out15_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out528_out1 <= in30 XOR in32;

  Logical_Operator_out529_out1 <= Logical_Operator_out17_out1 XOR Logical_Operator_out18_out1;

  Logical_Operator_out530_out1 <= in34 XOR in36;

  Logical_Operator_out531_out1 <= Logical_Operator_out19_out1 XOR Logical_Operator_out20_out1;

  Logical_Operator_out532_out1 <= in38 XOR in40;

  Logical_Operator_out533_out1 <= Logical_Operator_out21_out1 XOR Logical_Operator_out22_out1;

  Logical_Operator_out534_out1 <= in42 XOR in44;

  Logical_Operator_out535_out1 <= Logical_Operator_out23_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out536_out1 <= in46 XOR in48;

  Logical_Operator_out537_out1 <= Logical_Operator_out25_out1 XOR Logical_Operator_out26_out1;

  Logical_Operator_out538_out1 <= in50 XOR in52;

  Logical_Operator_out539_out1 <= Logical_Operator_out27_out1 XOR Logical_Operator_out28_out1;

  Logical_Operator_out540_out1 <= in54 XOR in56;

  Logical_Operator_out541_out1 <= Logical_Operator_out29_out1 XOR Logical_Operator_out30_out1;

  Logical_Operator_out542_out1 <= in58 XOR in60;

  Logical_Operator_out543_out1 <= Logical_Operator_out31_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out544_out1 <= in62 XOR in64;

  Logical_Operator_out545_out1 <= Logical_Operator_out33_out1 XOR Logical_Operator_out34_out1;

  Logical_Operator_out546_out1 <= in66 XOR in68;

  Logical_Operator_out547_out1 <= Logical_Operator_out35_out1 XOR Logical_Operator_out36_out1;

  Logical_Operator_out548_out1 <= in70 XOR in72;

  Logical_Operator_out549_out1 <= Logical_Operator_out37_out1 XOR Logical_Operator_out38_out1;

  Logical_Operator_out550_out1 <= in74 XOR in76;

  Logical_Operator_out551_out1 <= Logical_Operator_out39_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out552_out1 <= in78 XOR in80;

  Logical_Operator_out553_out1 <= Logical_Operator_out41_out1 XOR Logical_Operator_out42_out1;

  Logical_Operator_out554_out1 <= in82 XOR in84;

  Logical_Operator_out555_out1 <= Logical_Operator_out43_out1 XOR Logical_Operator_out44_out1;

  Logical_Operator_out556_out1 <= in86 XOR in88;

  Logical_Operator_out557_out1 <= Logical_Operator_out45_out1 XOR Logical_Operator_out46_out1;

  Logical_Operator_out558_out1 <= in90 XOR in92;

  Logical_Operator_out559_out1 <= Logical_Operator_out47_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out560_out1 <= in94 XOR in96;

  Logical_Operator_out561_out1 <= Logical_Operator_out49_out1 XOR Logical_Operator_out50_out1;

  Logical_Operator_out562_out1 <= in98 XOR in100;

  Logical_Operator_out563_out1 <= Logical_Operator_out51_out1 XOR Logical_Operator_out52_out1;

  Logical_Operator_out564_out1 <= in102 XOR in104;

  Logical_Operator_out565_out1 <= Logical_Operator_out53_out1 XOR Logical_Operator_out54_out1;

  Logical_Operator_out566_out1 <= in106 XOR in108;

  Logical_Operator_out567_out1 <= Logical_Operator_out55_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out568_out1 <= in110 XOR in112;

  Logical_Operator_out569_out1 <= Logical_Operator_out57_out1 XOR Logical_Operator_out58_out1;

  Logical_Operator_out570_out1 <= in114 XOR in116;

  Logical_Operator_out571_out1 <= Logical_Operator_out59_out1 XOR Logical_Operator_out60_out1;

  Logical_Operator_out572_out1 <= in118 XOR in120;

  Logical_Operator_out573_out1 <= Logical_Operator_out61_out1 XOR Logical_Operator_out62_out1;

  Logical_Operator_out574_out1 <= in122 XOR in124;

  Logical_Operator_out575_out1 <= Logical_Operator_out63_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out576_out1 <= in126 XOR in128;

  Logical_Operator_out577_out1 <= Logical_Operator_out65_out1 XOR Logical_Operator_out66_out1;

  Logical_Operator_out578_out1 <= in130 XOR in132;

  Logical_Operator_out579_out1 <= Logical_Operator_out67_out1 XOR Logical_Operator_out68_out1;

  Logical_Operator_out580_out1 <= in134 XOR in136;

  Logical_Operator_out581_out1 <= Logical_Operator_out69_out1 XOR Logical_Operator_out70_out1;

  Logical_Operator_out582_out1 <= in138 XOR in140;

  Logical_Operator_out583_out1 <= Logical_Operator_out71_out1 XOR Logical_Operator_out72_out1;

  Logical_Operator_out584_out1 <= in142 XOR in144;

  Logical_Operator_out585_out1 <= Logical_Operator_out73_out1 XOR Logical_Operator_out74_out1;

  Logical_Operator_out586_out1 <= in146 XOR in148;

  Logical_Operator_out587_out1 <= Logical_Operator_out75_out1 XOR Logical_Operator_out76_out1;

  Logical_Operator_out588_out1 <= in150 XOR in152;

  Logical_Operator_out589_out1 <= Logical_Operator_out77_out1 XOR Logical_Operator_out78_out1;

  Logical_Operator_out590_out1 <= in154 XOR in156;

  Logical_Operator_out591_out1 <= Logical_Operator_out79_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out592_out1 <= in158 XOR in160;

  Logical_Operator_out593_out1 <= Logical_Operator_out81_out1 XOR Logical_Operator_out82_out1;

  Logical_Operator_out594_out1 <= in162 XOR in164;

  Logical_Operator_out595_out1 <= Logical_Operator_out83_out1 XOR Logical_Operator_out84_out1;

  Logical_Operator_out596_out1 <= in166 XOR in168;

  Logical_Operator_out597_out1 <= Logical_Operator_out85_out1 XOR Logical_Operator_out86_out1;

  Logical_Operator_out598_out1 <= in170 XOR in172;

  Logical_Operator_out599_out1 <= Logical_Operator_out87_out1 XOR Logical_Operator_out88_out1;

  Logical_Operator_out600_out1 <= in174 XOR in176;

  Logical_Operator_out601_out1 <= Logical_Operator_out89_out1 XOR Logical_Operator_out90_out1;

  Logical_Operator_out602_out1 <= in178 XOR in180;

  Logical_Operator_out603_out1 <= Logical_Operator_out91_out1 XOR Logical_Operator_out92_out1;

  Logical_Operator_out604_out1 <= in182 XOR in184;

  Logical_Operator_out605_out1 <= Logical_Operator_out93_out1 XOR Logical_Operator_out94_out1;

  Logical_Operator_out606_out1 <= in186 XOR in188;

  Logical_Operator_out607_out1 <= Logical_Operator_out95_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out608_out1 <= in190 XOR in192;

  Logical_Operator_out609_out1 <= Logical_Operator_out97_out1 XOR Logical_Operator_out98_out1;

  Logical_Operator_out610_out1 <= in194 XOR in196;

  Logical_Operator_out611_out1 <= Logical_Operator_out99_out1 XOR Logical_Operator_out100_out1;

  Logical_Operator_out612_out1 <= in198 XOR in200;

  Logical_Operator_out613_out1 <= Logical_Operator_out101_out1 XOR Logical_Operator_out102_out1;

  Logical_Operator_out614_out1 <= in202 XOR in204;

  Logical_Operator_out615_out1 <= Logical_Operator_out103_out1 XOR Logical_Operator_out104_out1;

  Logical_Operator_out616_out1 <= in206 XOR in208;

  Logical_Operator_out617_out1 <= Logical_Operator_out105_out1 XOR Logical_Operator_out106_out1;

  Logical_Operator_out618_out1 <= in210 XOR in212;

  Logical_Operator_out619_out1 <= Logical_Operator_out107_out1 XOR Logical_Operator_out108_out1;

  Logical_Operator_out620_out1 <= in214 XOR in216;

  Logical_Operator_out621_out1 <= Logical_Operator_out109_out1 XOR Logical_Operator_out110_out1;

  Logical_Operator_out622_out1 <= in218 XOR in220;

  Logical_Operator_out623_out1 <= Logical_Operator_out111_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out624_out1 <= in222 XOR in224;

  Logical_Operator_out625_out1 <= Logical_Operator_out113_out1 XOR Logical_Operator_out114_out1;

  Logical_Operator_out626_out1 <= in226 XOR in228;

  Logical_Operator_out627_out1 <= Logical_Operator_out115_out1 XOR Logical_Operator_out116_out1;

  Logical_Operator_out628_out1 <= in230 XOR in232;

  Logical_Operator_out629_out1 <= Logical_Operator_out117_out1 XOR Logical_Operator_out118_out1;

  Logical_Operator_out630_out1 <= in234 XOR in236;

  Logical_Operator_out631_out1 <= Logical_Operator_out119_out1 XOR Logical_Operator_out120_out1;

  Logical_Operator_out632_out1 <= in238 XOR in240;

  Logical_Operator_out633_out1 <= Logical_Operator_out121_out1 XOR Logical_Operator_out122_out1;

  Logical_Operator_out634_out1 <= in242 XOR in244;

  Logical_Operator_out635_out1 <= Logical_Operator_out123_out1 XOR Logical_Operator_out124_out1;

  Logical_Operator_out636_out1 <= in246 XOR in248;

  Logical_Operator_out637_out1 <= Logical_Operator_out125_out1 XOR Logical_Operator_out126_out1;

  Logical_Operator_out638_out1 <= in250 XOR in252;

  Logical_Operator_out639_out1 <= Logical_Operator_out127_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out640_out1 <= in254 XOR in256;

  Logical_Operator_out641_out1 <= Logical_Operator_out129_out1 XOR Logical_Operator_out130_out1;

  Logical_Operator_out642_out1 <= in258 XOR in260;

  Logical_Operator_out643_out1 <= Logical_Operator_out131_out1 XOR Logical_Operator_out132_out1;

  Logical_Operator_out644_out1 <= in262 XOR in264;

  Logical_Operator_out645_out1 <= Logical_Operator_out133_out1 XOR Logical_Operator_out134_out1;

  Logical_Operator_out646_out1 <= in266 XOR in268;

  Logical_Operator_out647_out1 <= Logical_Operator_out135_out1 XOR Logical_Operator_out136_out1;

  Logical_Operator_out648_out1 <= in270 XOR in272;

  Logical_Operator_out649_out1 <= Logical_Operator_out137_out1 XOR Logical_Operator_out138_out1;

  Logical_Operator_out650_out1 <= in274 XOR in276;

  Logical_Operator_out651_out1 <= Logical_Operator_out139_out1 XOR Logical_Operator_out140_out1;

  Logical_Operator_out652_out1 <= in278 XOR in280;

  Logical_Operator_out653_out1 <= Logical_Operator_out141_out1 XOR Logical_Operator_out142_out1;

  Logical_Operator_out654_out1 <= in282 XOR in284;

  Logical_Operator_out655_out1 <= Logical_Operator_out143_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out656_out1 <= in286 XOR in288;

  Logical_Operator_out657_out1 <= Logical_Operator_out145_out1 XOR Logical_Operator_out146_out1;

  Logical_Operator_out658_out1 <= in290 XOR in292;

  Logical_Operator_out659_out1 <= Logical_Operator_out147_out1 XOR Logical_Operator_out148_out1;

  Logical_Operator_out660_out1 <= in294 XOR in296;

  Logical_Operator_out661_out1 <= Logical_Operator_out149_out1 XOR Logical_Operator_out150_out1;

  Logical_Operator_out662_out1 <= in298 XOR in300;

  Logical_Operator_out663_out1 <= Logical_Operator_out151_out1 XOR Logical_Operator_out152_out1;

  Logical_Operator_out664_out1 <= in302 XOR in304;

  Logical_Operator_out665_out1 <= Logical_Operator_out153_out1 XOR Logical_Operator_out154_out1;

  Logical_Operator_out666_out1 <= in306 XOR in308;

  Logical_Operator_out667_out1 <= Logical_Operator_out155_out1 XOR Logical_Operator_out156_out1;

  Logical_Operator_out668_out1 <= in310 XOR in312;

  Logical_Operator_out669_out1 <= Logical_Operator_out157_out1 XOR Logical_Operator_out158_out1;

  Logical_Operator_out670_out1 <= in314 XOR in316;

  Logical_Operator_out671_out1 <= Logical_Operator_out159_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out672_out1 <= in318 XOR in320;

  Logical_Operator_out673_out1 <= Logical_Operator_out161_out1 XOR Logical_Operator_out162_out1;

  Logical_Operator_out674_out1 <= in322 XOR in324;

  Logical_Operator_out675_out1 <= Logical_Operator_out163_out1 XOR Logical_Operator_out164_out1;

  Logical_Operator_out676_out1 <= in326 XOR in328;

  Logical_Operator_out677_out1 <= Logical_Operator_out165_out1 XOR Logical_Operator_out166_out1;

  Logical_Operator_out678_out1 <= in330 XOR in332;

  Logical_Operator_out679_out1 <= Logical_Operator_out167_out1 XOR Logical_Operator_out168_out1;

  Logical_Operator_out680_out1 <= in334 XOR in336;

  Logical_Operator_out681_out1 <= Logical_Operator_out169_out1 XOR Logical_Operator_out170_out1;

  Logical_Operator_out682_out1 <= in338 XOR in340;

  Logical_Operator_out683_out1 <= Logical_Operator_out171_out1 XOR Logical_Operator_out172_out1;

  Logical_Operator_out684_out1 <= in342 XOR in344;

  Logical_Operator_out685_out1 <= Logical_Operator_out173_out1 XOR Logical_Operator_out174_out1;

  Logical_Operator_out686_out1 <= in346 XOR in348;

  Logical_Operator_out687_out1 <= Logical_Operator_out175_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out688_out1 <= in350 XOR in352;

  Logical_Operator_out689_out1 <= Logical_Operator_out177_out1 XOR Logical_Operator_out178_out1;

  Logical_Operator_out690_out1 <= in354 XOR in356;

  Logical_Operator_out691_out1 <= Logical_Operator_out179_out1 XOR Logical_Operator_out180_out1;

  Logical_Operator_out692_out1 <= in358 XOR in360;

  Logical_Operator_out693_out1 <= Logical_Operator_out181_out1 XOR Logical_Operator_out182_out1;

  Logical_Operator_out694_out1 <= in362 XOR in364;

  Logical_Operator_out695_out1 <= Logical_Operator_out183_out1 XOR Logical_Operator_out184_out1;

  Logical_Operator_out696_out1 <= in366 XOR in368;

  Logical_Operator_out697_out1 <= Logical_Operator_out185_out1 XOR Logical_Operator_out186_out1;

  Logical_Operator_out698_out1 <= in370 XOR in372;

  Logical_Operator_out699_out1 <= Logical_Operator_out187_out1 XOR Logical_Operator_out188_out1;

  Logical_Operator_out700_out1 <= in374 XOR in376;

  Logical_Operator_out701_out1 <= Logical_Operator_out189_out1 XOR Logical_Operator_out190_out1;

  Logical_Operator_out702_out1 <= in378 XOR in380;

  Logical_Operator_out703_out1 <= Logical_Operator_out191_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out704_out1 <= in382 XOR in384;

  Logical_Operator_out705_out1 <= Logical_Operator_out193_out1 XOR Logical_Operator_out194_out1;

  Logical_Operator_out706_out1 <= in386 XOR in388;

  Logical_Operator_out707_out1 <= Logical_Operator_out195_out1 XOR Logical_Operator_out196_out1;

  Logical_Operator_out708_out1 <= in390 XOR in392;

  Logical_Operator_out709_out1 <= Logical_Operator_out197_out1 XOR Logical_Operator_out198_out1;

  Logical_Operator_out710_out1 <= in394 XOR in396;

  Logical_Operator_out711_out1 <= Logical_Operator_out199_out1 XOR Logical_Operator_out200_out1;

  Logical_Operator_out712_out1 <= in398 XOR in400;

  Logical_Operator_out713_out1 <= Logical_Operator_out201_out1 XOR Logical_Operator_out202_out1;

  Logical_Operator_out714_out1 <= in402 XOR in404;

  Logical_Operator_out715_out1 <= Logical_Operator_out203_out1 XOR Logical_Operator_out204_out1;

  Logical_Operator_out716_out1 <= in406 XOR in408;

  Logical_Operator_out717_out1 <= Logical_Operator_out205_out1 XOR Logical_Operator_out206_out1;

  Logical_Operator_out718_out1 <= in410 XOR in412;

  Logical_Operator_out719_out1 <= Logical_Operator_out207_out1 XOR Logical_Operator_out208_out1;

  Logical_Operator_out720_out1 <= in414 XOR in416;

  Logical_Operator_out721_out1 <= Logical_Operator_out209_out1 XOR Logical_Operator_out210_out1;

  Logical_Operator_out722_out1 <= in418 XOR in420;

  Logical_Operator_out723_out1 <= Logical_Operator_out211_out1 XOR Logical_Operator_out212_out1;

  Logical_Operator_out724_out1 <= in422 XOR in424;

  Logical_Operator_out725_out1 <= Logical_Operator_out213_out1 XOR Logical_Operator_out214_out1;

  Logical_Operator_out726_out1 <= in426 XOR in428;

  Logical_Operator_out727_out1 <= Logical_Operator_out215_out1 XOR Logical_Operator_out216_out1;

  Logical_Operator_out728_out1 <= in430 XOR in432;

  Logical_Operator_out729_out1 <= Logical_Operator_out217_out1 XOR Logical_Operator_out218_out1;

  Logical_Operator_out730_out1 <= in434 XOR in436;

  Logical_Operator_out731_out1 <= Logical_Operator_out219_out1 XOR Logical_Operator_out220_out1;

  Logical_Operator_out732_out1 <= in438 XOR in440;

  Logical_Operator_out733_out1 <= Logical_Operator_out221_out1 XOR Logical_Operator_out222_out1;

  Logical_Operator_out734_out1 <= in442 XOR in444;

  Logical_Operator_out735_out1 <= Logical_Operator_out223_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out736_out1 <= in446 XOR in448;

  Logical_Operator_out737_out1 <= Logical_Operator_out225_out1 XOR Logical_Operator_out226_out1;

  Logical_Operator_out738_out1 <= in450 XOR in452;

  Logical_Operator_out739_out1 <= Logical_Operator_out227_out1 XOR Logical_Operator_out228_out1;

  Logical_Operator_out740_out1 <= in454 XOR in456;

  Logical_Operator_out741_out1 <= Logical_Operator_out229_out1 XOR Logical_Operator_out230_out1;

  Logical_Operator_out742_out1 <= in458 XOR in460;

  Logical_Operator_out743_out1 <= Logical_Operator_out231_out1 XOR Logical_Operator_out232_out1;

  Logical_Operator_out744_out1 <= in462 XOR in464;

  Logical_Operator_out745_out1 <= Logical_Operator_out233_out1 XOR Logical_Operator_out234_out1;

  Logical_Operator_out746_out1 <= in466 XOR in468;

  Logical_Operator_out747_out1 <= Logical_Operator_out235_out1 XOR Logical_Operator_out236_out1;

  Logical_Operator_out748_out1 <= in470 XOR in472;

  Logical_Operator_out749_out1 <= Logical_Operator_out237_out1 XOR Logical_Operator_out238_out1;

  Logical_Operator_out750_out1 <= in474 XOR in476;

  Logical_Operator_out751_out1 <= Logical_Operator_out239_out1 XOR Logical_Operator_out240_out1;

  Logical_Operator_out752_out1 <= in478 XOR in480;

  Logical_Operator_out753_out1 <= Logical_Operator_out241_out1 XOR Logical_Operator_out242_out1;

  Logical_Operator_out754_out1 <= in482 XOR in484;

  Logical_Operator_out755_out1 <= Logical_Operator_out243_out1 XOR Logical_Operator_out244_out1;

  Logical_Operator_out756_out1 <= in486 XOR in488;

  Logical_Operator_out757_out1 <= Logical_Operator_out245_out1 XOR Logical_Operator_out246_out1;

  Logical_Operator_out758_out1 <= in490 XOR in492;

  Logical_Operator_out759_out1 <= Logical_Operator_out247_out1 XOR Logical_Operator_out248_out1;

  Logical_Operator_out760_out1 <= in494 XOR in496;

  Logical_Operator_out761_out1 <= Logical_Operator_out249_out1 XOR Logical_Operator_out250_out1;

  Logical_Operator_out762_out1 <= in498 XOR in500;

  Logical_Operator_out763_out1 <= Logical_Operator_out251_out1 XOR Logical_Operator_out252_out1;

  Logical_Operator_out764_out1 <= in502 XOR in504;

  Logical_Operator_out765_out1 <= Logical_Operator_out253_out1 XOR Logical_Operator_out254_out1;

  Logical_Operator_out766_out1 <= in506 XOR in508;

  Logical_Operator_out767_out1 <= Logical_Operator_out255_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out768_out1 <= in510 XOR in512;

  Logical_Operator_out769_out1 <= Logical_Operator_out257_out1 XOR Logical_Operator_out258_out1;

  Logical_Operator_out770_out1 <= in514 XOR in516;

  Logical_Operator_out771_out1 <= Logical_Operator_out259_out1 XOR Logical_Operator_out260_out1;

  Logical_Operator_out772_out1 <= in518 XOR in520;

  Logical_Operator_out773_out1 <= Logical_Operator_out261_out1 XOR Logical_Operator_out262_out1;

  Logical_Operator_out774_out1 <= in522 XOR in524;

  Logical_Operator_out775_out1 <= Logical_Operator_out263_out1 XOR Logical_Operator_out264_out1;

  Logical_Operator_out776_out1 <= in526 XOR in528;

  Logical_Operator_out777_out1 <= Logical_Operator_out265_out1 XOR Logical_Operator_out266_out1;

  Logical_Operator_out778_out1 <= in530 XOR in532;

  Logical_Operator_out779_out1 <= Logical_Operator_out267_out1 XOR Logical_Operator_out268_out1;

  Logical_Operator_out780_out1 <= in534 XOR in536;

  Logical_Operator_out781_out1 <= Logical_Operator_out269_out1 XOR Logical_Operator_out270_out1;

  Logical_Operator_out782_out1 <= in538 XOR in540;

  Logical_Operator_out783_out1 <= Logical_Operator_out271_out1 XOR Logical_Operator_out272_out1;

  Logical_Operator_out784_out1 <= in542 XOR in544;

  Logical_Operator_out785_out1 <= Logical_Operator_out273_out1 XOR Logical_Operator_out274_out1;

  Logical_Operator_out786_out1 <= in546 XOR in548;

  Logical_Operator_out787_out1 <= Logical_Operator_out275_out1 XOR Logical_Operator_out276_out1;

  Logical_Operator_out788_out1 <= in550 XOR in552;

  Logical_Operator_out789_out1 <= Logical_Operator_out277_out1 XOR Logical_Operator_out278_out1;

  Logical_Operator_out790_out1 <= in554 XOR in556;

  Logical_Operator_out791_out1 <= Logical_Operator_out279_out1 XOR Logical_Operator_out280_out1;

  Logical_Operator_out792_out1 <= in558 XOR in560;

  Logical_Operator_out793_out1 <= Logical_Operator_out281_out1 XOR Logical_Operator_out282_out1;

  Logical_Operator_out794_out1 <= in562 XOR in564;

  Logical_Operator_out795_out1 <= Logical_Operator_out283_out1 XOR Logical_Operator_out284_out1;

  Logical_Operator_out796_out1 <= in566 XOR in568;

  Logical_Operator_out797_out1 <= Logical_Operator_out285_out1 XOR Logical_Operator_out286_out1;

  Logical_Operator_out798_out1 <= in570 XOR in572;

  Logical_Operator_out799_out1 <= Logical_Operator_out287_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out800_out1 <= in574 XOR in576;

  Logical_Operator_out801_out1 <= Logical_Operator_out289_out1 XOR Logical_Operator_out290_out1;

  Logical_Operator_out802_out1 <= in578 XOR in580;

  Logical_Operator_out803_out1 <= Logical_Operator_out291_out1 XOR Logical_Operator_out292_out1;

  Logical_Operator_out804_out1 <= in582 XOR in584;

  Logical_Operator_out805_out1 <= Logical_Operator_out293_out1 XOR Logical_Operator_out294_out1;

  Logical_Operator_out806_out1 <= in586 XOR in588;

  Logical_Operator_out807_out1 <= Logical_Operator_out295_out1 XOR Logical_Operator_out296_out1;

  Logical_Operator_out808_out1 <= in590 XOR in592;

  Logical_Operator_out809_out1 <= Logical_Operator_out297_out1 XOR Logical_Operator_out298_out1;

  Logical_Operator_out810_out1 <= in594 XOR in596;

  Logical_Operator_out811_out1 <= Logical_Operator_out299_out1 XOR Logical_Operator_out300_out1;

  Logical_Operator_out812_out1 <= in598 XOR in600;

  Logical_Operator_out813_out1 <= Logical_Operator_out301_out1 XOR Logical_Operator_out302_out1;

  Logical_Operator_out814_out1 <= in602 XOR in604;

  Logical_Operator_out815_out1 <= Logical_Operator_out303_out1 XOR Logical_Operator_out304_out1;

  Logical_Operator_out816_out1 <= in606 XOR in608;

  Logical_Operator_out817_out1 <= Logical_Operator_out305_out1 XOR Logical_Operator_out306_out1;

  Logical_Operator_out818_out1 <= in610 XOR in612;

  Logical_Operator_out819_out1 <= Logical_Operator_out307_out1 XOR Logical_Operator_out308_out1;

  Logical_Operator_out820_out1 <= in614 XOR in616;

  Logical_Operator_out821_out1 <= Logical_Operator_out309_out1 XOR Logical_Operator_out310_out1;

  Logical_Operator_out822_out1 <= in618 XOR in620;

  Logical_Operator_out823_out1 <= Logical_Operator_out311_out1 XOR Logical_Operator_out312_out1;

  Logical_Operator_out824_out1 <= in622 XOR in624;

  Logical_Operator_out825_out1 <= Logical_Operator_out313_out1 XOR Logical_Operator_out314_out1;

  Logical_Operator_out826_out1 <= in626 XOR in628;

  Logical_Operator_out827_out1 <= Logical_Operator_out315_out1 XOR Logical_Operator_out316_out1;

  Logical_Operator_out828_out1 <= in630 XOR in632;

  Logical_Operator_out829_out1 <= Logical_Operator_out317_out1 XOR Logical_Operator_out318_out1;

  Logical_Operator_out830_out1 <= in634 XOR in636;

  Logical_Operator_out831_out1 <= Logical_Operator_out319_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out832_out1 <= in638 XOR in640;

  Logical_Operator_out833_out1 <= Logical_Operator_out321_out1 XOR Logical_Operator_out322_out1;

  Logical_Operator_out834_out1 <= in642 XOR in644;

  Logical_Operator_out835_out1 <= Logical_Operator_out323_out1 XOR Logical_Operator_out324_out1;

  Logical_Operator_out836_out1 <= in646 XOR in648;

  Logical_Operator_out837_out1 <= Logical_Operator_out325_out1 XOR Logical_Operator_out326_out1;

  Logical_Operator_out838_out1 <= in650 XOR in652;

  Logical_Operator_out839_out1 <= Logical_Operator_out327_out1 XOR Logical_Operator_out328_out1;

  Logical_Operator_out840_out1 <= in654 XOR in656;

  Logical_Operator_out841_out1 <= Logical_Operator_out329_out1 XOR Logical_Operator_out330_out1;

  Logical_Operator_out842_out1 <= in658 XOR in660;

  Logical_Operator_out843_out1 <= Logical_Operator_out331_out1 XOR Logical_Operator_out332_out1;

  Logical_Operator_out844_out1 <= in662 XOR in664;

  Logical_Operator_out845_out1 <= Logical_Operator_out333_out1 XOR Logical_Operator_out334_out1;

  Logical_Operator_out846_out1 <= in666 XOR in668;

  Logical_Operator_out847_out1 <= Logical_Operator_out335_out1 XOR Logical_Operator_out336_out1;

  Logical_Operator_out848_out1 <= in670 XOR in672;

  Logical_Operator_out849_out1 <= Logical_Operator_out337_out1 XOR Logical_Operator_out338_out1;

  Logical_Operator_out850_out1 <= in674 XOR in676;

  Logical_Operator_out851_out1 <= Logical_Operator_out339_out1 XOR Logical_Operator_out340_out1;

  Logical_Operator_out852_out1 <= in678 XOR in680;

  Logical_Operator_out853_out1 <= Logical_Operator_out341_out1 XOR Logical_Operator_out342_out1;

  Logical_Operator_out854_out1 <= in682 XOR in684;

  Logical_Operator_out855_out1 <= Logical_Operator_out343_out1 XOR Logical_Operator_out344_out1;

  Logical_Operator_out856_out1 <= in686 XOR in688;

  Logical_Operator_out857_out1 <= Logical_Operator_out345_out1 XOR Logical_Operator_out346_out1;

  Logical_Operator_out858_out1 <= in690 XOR in692;

  Logical_Operator_out859_out1 <= Logical_Operator_out347_out1 XOR Logical_Operator_out348_out1;

  Logical_Operator_out860_out1 <= in694 XOR in696;

  Logical_Operator_out861_out1 <= Logical_Operator_out349_out1 XOR Logical_Operator_out350_out1;

  Logical_Operator_out862_out1 <= in698 XOR in700;

  Logical_Operator_out863_out1 <= Logical_Operator_out351_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out864_out1 <= in702 XOR in704;

  Logical_Operator_out865_out1 <= Logical_Operator_out353_out1 XOR Logical_Operator_out354_out1;

  Logical_Operator_out866_out1 <= in706 XOR in708;

  Logical_Operator_out867_out1 <= Logical_Operator_out355_out1 XOR Logical_Operator_out356_out1;

  Logical_Operator_out868_out1 <= in710 XOR in712;

  Logical_Operator_out869_out1 <= Logical_Operator_out357_out1 XOR Logical_Operator_out358_out1;

  Logical_Operator_out870_out1 <= in714 XOR in716;

  Logical_Operator_out871_out1 <= Logical_Operator_out359_out1 XOR Logical_Operator_out360_out1;

  Logical_Operator_out872_out1 <= in718 XOR in720;

  Logical_Operator_out873_out1 <= Logical_Operator_out361_out1 XOR Logical_Operator_out362_out1;

  Logical_Operator_out874_out1 <= in722 XOR in724;

  Logical_Operator_out875_out1 <= Logical_Operator_out363_out1 XOR Logical_Operator_out364_out1;

  Logical_Operator_out876_out1 <= in726 XOR in728;

  Logical_Operator_out877_out1 <= Logical_Operator_out365_out1 XOR Logical_Operator_out366_out1;

  Logical_Operator_out878_out1 <= in730 XOR in732;

  Logical_Operator_out879_out1 <= Logical_Operator_out367_out1 XOR Logical_Operator_out368_out1;

  Logical_Operator_out880_out1 <= in734 XOR in736;

  Logical_Operator_out881_out1 <= Logical_Operator_out369_out1 XOR Logical_Operator_out370_out1;

  Logical_Operator_out882_out1 <= in738 XOR in740;

  Logical_Operator_out883_out1 <= Logical_Operator_out371_out1 XOR Logical_Operator_out372_out1;

  Logical_Operator_out884_out1 <= in742 XOR in744;

  Logical_Operator_out885_out1 <= Logical_Operator_out373_out1 XOR Logical_Operator_out374_out1;

  Logical_Operator_out886_out1 <= in746 XOR in748;

  Logical_Operator_out887_out1 <= Logical_Operator_out375_out1 XOR Logical_Operator_out376_out1;

  Logical_Operator_out888_out1 <= in750 XOR in752;

  Logical_Operator_out889_out1 <= Logical_Operator_out377_out1 XOR Logical_Operator_out378_out1;

  Logical_Operator_out890_out1 <= in754 XOR in756;

  Logical_Operator_out891_out1 <= Logical_Operator_out379_out1 XOR Logical_Operator_out380_out1;

  Logical_Operator_out892_out1 <= in758 XOR in760;

  Logical_Operator_out893_out1 <= Logical_Operator_out381_out1 XOR Logical_Operator_out382_out1;

  Logical_Operator_out894_out1 <= in762 XOR in764;

  Logical_Operator_out895_out1 <= Logical_Operator_out383_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out896_out1 <= in766 XOR in768;

  Logical_Operator_out897_out1 <= Logical_Operator_out385_out1 XOR Logical_Operator_out386_out1;

  Logical_Operator_out898_out1 <= in770 XOR in772;

  Logical_Operator_out899_out1 <= Logical_Operator_out387_out1 XOR Logical_Operator_out388_out1;

  Logical_Operator_out900_out1 <= in774 XOR in776;

  Logical_Operator_out901_out1 <= Logical_Operator_out389_out1 XOR Logical_Operator_out390_out1;

  Logical_Operator_out902_out1 <= in778 XOR in780;

  Logical_Operator_out903_out1 <= Logical_Operator_out391_out1 XOR Logical_Operator_out392_out1;

  Logical_Operator_out904_out1 <= in782 XOR in784;

  Logical_Operator_out905_out1 <= Logical_Operator_out393_out1 XOR Logical_Operator_out394_out1;

  Logical_Operator_out906_out1 <= in786 XOR in788;

  Logical_Operator_out907_out1 <= Logical_Operator_out395_out1 XOR Logical_Operator_out396_out1;

  Logical_Operator_out908_out1 <= in790 XOR in792;

  Logical_Operator_out909_out1 <= Logical_Operator_out397_out1 XOR Logical_Operator_out398_out1;

  Logical_Operator_out910_out1 <= in794 XOR in796;

  Logical_Operator_out911_out1 <= Logical_Operator_out399_out1 XOR Logical_Operator_out400_out1;

  Logical_Operator_out912_out1 <= in798 XOR in800;

  Logical_Operator_out913_out1 <= Logical_Operator_out401_out1 XOR Logical_Operator_out402_out1;

  Logical_Operator_out914_out1 <= in802 XOR in804;

  Logical_Operator_out915_out1 <= Logical_Operator_out403_out1 XOR Logical_Operator_out404_out1;

  Logical_Operator_out916_out1 <= in806 XOR in808;

  Logical_Operator_out917_out1 <= Logical_Operator_out405_out1 XOR Logical_Operator_out406_out1;

  Logical_Operator_out918_out1 <= in810 XOR in812;

  Logical_Operator_out919_out1 <= Logical_Operator_out407_out1 XOR Logical_Operator_out408_out1;

  Logical_Operator_out920_out1 <= in814 XOR in816;

  Logical_Operator_out921_out1 <= Logical_Operator_out409_out1 XOR Logical_Operator_out410_out1;

  Logical_Operator_out922_out1 <= in818 XOR in820;

  Logical_Operator_out923_out1 <= Logical_Operator_out411_out1 XOR Logical_Operator_out412_out1;

  Logical_Operator_out924_out1 <= in822 XOR in824;

  Logical_Operator_out925_out1 <= Logical_Operator_out413_out1 XOR Logical_Operator_out414_out1;

  Logical_Operator_out926_out1 <= in826 XOR in828;

  Logical_Operator_out927_out1 <= Logical_Operator_out415_out1 XOR Logical_Operator_out416_out1;

  Logical_Operator_out928_out1 <= in830 XOR in832;

  Logical_Operator_out929_out1 <= Logical_Operator_out417_out1 XOR Logical_Operator_out418_out1;

  Logical_Operator_out930_out1 <= in834 XOR in836;

  Logical_Operator_out931_out1 <= Logical_Operator_out419_out1 XOR Logical_Operator_out420_out1;

  Logical_Operator_out932_out1 <= in838 XOR in840;

  Logical_Operator_out933_out1 <= Logical_Operator_out421_out1 XOR Logical_Operator_out422_out1;

  Logical_Operator_out934_out1 <= in842 XOR in844;

  Logical_Operator_out935_out1 <= Logical_Operator_out423_out1 XOR Logical_Operator_out424_out1;

  Logical_Operator_out936_out1 <= in846 XOR in848;

  Logical_Operator_out937_out1 <= Logical_Operator_out425_out1 XOR Logical_Operator_out426_out1;

  Logical_Operator_out938_out1 <= in850 XOR in852;

  Logical_Operator_out939_out1 <= Logical_Operator_out427_out1 XOR Logical_Operator_out428_out1;

  Logical_Operator_out940_out1 <= in854 XOR in856;

  Logical_Operator_out941_out1 <= Logical_Operator_out429_out1 XOR Logical_Operator_out430_out1;

  Logical_Operator_out942_out1 <= in858 XOR in860;

  Logical_Operator_out943_out1 <= Logical_Operator_out431_out1 XOR Logical_Operator_out432_out1;

  Logical_Operator_out944_out1 <= in862 XOR in864;

  Logical_Operator_out945_out1 <= Logical_Operator_out433_out1 XOR Logical_Operator_out434_out1;

  Logical_Operator_out946_out1 <= in866 XOR in868;

  Logical_Operator_out947_out1 <= Logical_Operator_out435_out1 XOR Logical_Operator_out436_out1;

  Logical_Operator_out948_out1 <= in870 XOR in872;

  Logical_Operator_out949_out1 <= Logical_Operator_out437_out1 XOR Logical_Operator_out438_out1;

  Logical_Operator_out950_out1 <= in874 XOR in876;

  Logical_Operator_out951_out1 <= Logical_Operator_out439_out1 XOR Logical_Operator_out440_out1;

  Logical_Operator_out952_out1 <= in878 XOR in880;

  Logical_Operator_out953_out1 <= Logical_Operator_out441_out1 XOR Logical_Operator_out442_out1;

  Logical_Operator_out954_out1 <= in882 XOR in884;

  Logical_Operator_out955_out1 <= Logical_Operator_out443_out1 XOR Logical_Operator_out444_out1;

  Logical_Operator_out956_out1 <= in886 XOR in888;

  Logical_Operator_out957_out1 <= Logical_Operator_out445_out1 XOR Logical_Operator_out446_out1;

  Logical_Operator_out958_out1 <= in890 XOR in892;

  Logical_Operator_out959_out1 <= Logical_Operator_out447_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out960_out1 <= in894 XOR in896;

  Logical_Operator_out961_out1 <= Logical_Operator_out449_out1 XOR Logical_Operator_out450_out1;

  Logical_Operator_out962_out1 <= in898 XOR in900;

  Logical_Operator_out963_out1 <= Logical_Operator_out451_out1 XOR Logical_Operator_out452_out1;

  Logical_Operator_out964_out1 <= in902 XOR in904;

  Logical_Operator_out965_out1 <= Logical_Operator_out453_out1 XOR Logical_Operator_out454_out1;

  Logical_Operator_out966_out1 <= in906 XOR in908;

  Logical_Operator_out967_out1 <= Logical_Operator_out455_out1 XOR Logical_Operator_out456_out1;

  Logical_Operator_out968_out1 <= in910 XOR in912;

  Logical_Operator_out969_out1 <= Logical_Operator_out457_out1 XOR Logical_Operator_out458_out1;

  Logical_Operator_out970_out1 <= in914 XOR in916;

  Logical_Operator_out971_out1 <= Logical_Operator_out459_out1 XOR Logical_Operator_out460_out1;

  Logical_Operator_out972_out1 <= in918 XOR in920;

  Logical_Operator_out973_out1 <= Logical_Operator_out461_out1 XOR Logical_Operator_out462_out1;

  Logical_Operator_out974_out1 <= in922 XOR in924;

  Logical_Operator_out975_out1 <= Logical_Operator_out463_out1 XOR Logical_Operator_out464_out1;

  Logical_Operator_out976_out1 <= in926 XOR in928;

  Logical_Operator_out977_out1 <= Logical_Operator_out465_out1 XOR Logical_Operator_out466_out1;

  Logical_Operator_out978_out1 <= in930 XOR in932;

  Logical_Operator_out979_out1 <= Logical_Operator_out467_out1 XOR Logical_Operator_out468_out1;

  Logical_Operator_out980_out1 <= in934 XOR in936;

  Logical_Operator_out981_out1 <= Logical_Operator_out469_out1 XOR Logical_Operator_out470_out1;

  Logical_Operator_out982_out1 <= in938 XOR in940;

  Logical_Operator_out983_out1 <= Logical_Operator_out471_out1 XOR Logical_Operator_out472_out1;

  Logical_Operator_out984_out1 <= in942 XOR in944;

  Logical_Operator_out985_out1 <= Logical_Operator_out473_out1 XOR Logical_Operator_out474_out1;

  Logical_Operator_out986_out1 <= in946 XOR in948;

  Logical_Operator_out987_out1 <= Logical_Operator_out475_out1 XOR Logical_Operator_out476_out1;

  Logical_Operator_out988_out1 <= in950 XOR in952;

  Logical_Operator_out989_out1 <= Logical_Operator_out477_out1 XOR Logical_Operator_out478_out1;

  Logical_Operator_out990_out1 <= in954 XOR in956;

  Logical_Operator_out991_out1 <= Logical_Operator_out479_out1 XOR Logical_Operator_out480_out1;

  Logical_Operator_out992_out1 <= in958 XOR in960;

  Logical_Operator_out993_out1 <= Logical_Operator_out481_out1 XOR Logical_Operator_out482_out1;

  Logical_Operator_out994_out1 <= in962 XOR in964;

  Logical_Operator_out995_out1 <= Logical_Operator_out483_out1 XOR Logical_Operator_out484_out1;

  Logical_Operator_out996_out1 <= in966 XOR in968;

  Logical_Operator_out997_out1 <= Logical_Operator_out485_out1 XOR Logical_Operator_out486_out1;

  Logical_Operator_out998_out1 <= in970 XOR in972;

  Logical_Operator_out999_out1 <= Logical_Operator_out487_out1 XOR Logical_Operator_out488_out1;

  Logical_Operator_out1000_out1 <= in974 XOR in976;

  Logical_Operator_out1001_out1 <= Logical_Operator_out489_out1 XOR Logical_Operator_out490_out1;

  Logical_Operator_out1002_out1 <= in978 XOR in980;

  Logical_Operator_out1003_out1 <= Logical_Operator_out491_out1 XOR Logical_Operator_out492_out1;

  Logical_Operator_out1004_out1 <= in982 XOR in984;

  Logical_Operator_out1005_out1 <= Logical_Operator_out493_out1 XOR Logical_Operator_out494_out1;

  Logical_Operator_out1006_out1 <= in986 XOR in988;

  Logical_Operator_out1007_out1 <= Logical_Operator_out495_out1 XOR Logical_Operator_out496_out1;

  Logical_Operator_out1008_out1 <= in990 XOR in992;

  Logical_Operator_out1009_out1 <= Logical_Operator_out497_out1 XOR Logical_Operator_out498_out1;

  Logical_Operator_out1010_out1 <= in994 XOR in996;

  Logical_Operator_out1011_out1 <= Logical_Operator_out499_out1 XOR Logical_Operator_out500_out1;

  Logical_Operator_out1012_out1 <= in998 XOR in1000;

  Logical_Operator_out1013_out1 <= Logical_Operator_out501_out1 XOR Logical_Operator_out502_out1;

  Logical_Operator_out1014_out1 <= in1002 XOR in1004;

  Logical_Operator_out1015_out1 <= Logical_Operator_out503_out1 XOR Logical_Operator_out504_out1;

  Logical_Operator_out1016_out1 <= in1006 XOR in1008;

  Logical_Operator_out1017_out1 <= Logical_Operator_out505_out1 XOR Logical_Operator_out506_out1;

  Logical_Operator_out1018_out1 <= in1010 XOR in1012;

  Logical_Operator_out1019_out1 <= Logical_Operator_out507_out1 XOR Logical_Operator_out508_out1;

  Logical_Operator_out1020_out1 <= in1014 XOR in1016;

  Logical_Operator_out1021_out1 <= Logical_Operator_out509_out1 XOR Logical_Operator_out510_out1;

  Logical_Operator_out1022_out1 <= in1018 XOR in1020;

  Logical_Operator_out1023_out1 <= Logical_Operator_out511_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out1024_out1 <= in1022 XOR in1024;

  Logical_Operator_out1025_out1 <= Logical_Operator_out513_out1 XOR Logical_Operator_out515_out1;

  Logical_Operator_out1026_out1 <= Logical_Operator_out514_out1 XOR Logical_Operator_out516_out1;

  Logical_Operator_out1027_out1 <= Logical_Operator_out2_out1 XOR Logical_Operator_out4_out1;

  Logical_Operator_out1028_out1 <= in4 XOR in8;

  Logical_Operator_out1029_out1 <= Logical_Operator_out517_out1 XOR Logical_Operator_out519_out1;

  Logical_Operator_out1030_out1 <= Logical_Operator_out518_out1 XOR Logical_Operator_out520_out1;

  Logical_Operator_out1031_out1 <= Logical_Operator_out6_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out1032_out1 <= in12 XOR in16;

  Logical_Operator_out1033_out1 <= Logical_Operator_out521_out1 XOR Logical_Operator_out523_out1;

  Logical_Operator_out1034_out1 <= Logical_Operator_out522_out1 XOR Logical_Operator_out524_out1;

  Logical_Operator_out1035_out1 <= Logical_Operator_out10_out1 XOR Logical_Operator_out12_out1;

  Logical_Operator_out1036_out1 <= in20 XOR in24;

  Logical_Operator_out1037_out1 <= Logical_Operator_out525_out1 XOR Logical_Operator_out527_out1;

  Logical_Operator_out1038_out1 <= Logical_Operator_out526_out1 XOR Logical_Operator_out528_out1;

  Logical_Operator_out1039_out1 <= Logical_Operator_out14_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out1040_out1 <= in28 XOR in32;

  Logical_Operator_out1041_out1 <= Logical_Operator_out529_out1 XOR Logical_Operator_out531_out1;

  Logical_Operator_out1042_out1 <= Logical_Operator_out530_out1 XOR Logical_Operator_out532_out1;

  Logical_Operator_out1043_out1 <= Logical_Operator_out18_out1 XOR Logical_Operator_out20_out1;

  Logical_Operator_out1044_out1 <= in36 XOR in40;

  Logical_Operator_out1045_out1 <= Logical_Operator_out533_out1 XOR Logical_Operator_out535_out1;

  Logical_Operator_out1046_out1 <= Logical_Operator_out534_out1 XOR Logical_Operator_out536_out1;

  Logical_Operator_out1047_out1 <= Logical_Operator_out22_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out1048_out1 <= in44 XOR in48;

  Logical_Operator_out1049_out1 <= Logical_Operator_out537_out1 XOR Logical_Operator_out539_out1;

  Logical_Operator_out1050_out1 <= Logical_Operator_out538_out1 XOR Logical_Operator_out540_out1;

  Logical_Operator_out1051_out1 <= Logical_Operator_out26_out1 XOR Logical_Operator_out28_out1;

  Logical_Operator_out1052_out1 <= in52 XOR in56;

  Logical_Operator_out1053_out1 <= Logical_Operator_out541_out1 XOR Logical_Operator_out543_out1;

  Logical_Operator_out1054_out1 <= Logical_Operator_out542_out1 XOR Logical_Operator_out544_out1;

  Logical_Operator_out1055_out1 <= Logical_Operator_out30_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out1056_out1 <= in60 XOR in64;

  Logical_Operator_out1057_out1 <= Logical_Operator_out545_out1 XOR Logical_Operator_out547_out1;

  Logical_Operator_out1058_out1 <= Logical_Operator_out546_out1 XOR Logical_Operator_out548_out1;

  Logical_Operator_out1059_out1 <= Logical_Operator_out34_out1 XOR Logical_Operator_out36_out1;

  Logical_Operator_out1060_out1 <= in68 XOR in72;

  Logical_Operator_out1061_out1 <= Logical_Operator_out549_out1 XOR Logical_Operator_out551_out1;

  Logical_Operator_out1062_out1 <= Logical_Operator_out550_out1 XOR Logical_Operator_out552_out1;

  Logical_Operator_out1063_out1 <= Logical_Operator_out38_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out1064_out1 <= in76 XOR in80;

  Logical_Operator_out1065_out1 <= Logical_Operator_out553_out1 XOR Logical_Operator_out555_out1;

  Logical_Operator_out1066_out1 <= Logical_Operator_out554_out1 XOR Logical_Operator_out556_out1;

  Logical_Operator_out1067_out1 <= Logical_Operator_out42_out1 XOR Logical_Operator_out44_out1;

  Logical_Operator_out1068_out1 <= in84 XOR in88;

  Logical_Operator_out1069_out1 <= Logical_Operator_out557_out1 XOR Logical_Operator_out559_out1;

  Logical_Operator_out1070_out1 <= Logical_Operator_out558_out1 XOR Logical_Operator_out560_out1;

  Logical_Operator_out1071_out1 <= Logical_Operator_out46_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out1072_out1 <= in92 XOR in96;

  Logical_Operator_out1073_out1 <= Logical_Operator_out561_out1 XOR Logical_Operator_out563_out1;

  Logical_Operator_out1074_out1 <= Logical_Operator_out562_out1 XOR Logical_Operator_out564_out1;

  Logical_Operator_out1075_out1 <= Logical_Operator_out50_out1 XOR Logical_Operator_out52_out1;

  Logical_Operator_out1076_out1 <= in100 XOR in104;

  Logical_Operator_out1077_out1 <= Logical_Operator_out565_out1 XOR Logical_Operator_out567_out1;

  Logical_Operator_out1078_out1 <= Logical_Operator_out566_out1 XOR Logical_Operator_out568_out1;

  Logical_Operator_out1079_out1 <= Logical_Operator_out54_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out1080_out1 <= in108 XOR in112;

  Logical_Operator_out1081_out1 <= Logical_Operator_out569_out1 XOR Logical_Operator_out571_out1;

  Logical_Operator_out1082_out1 <= Logical_Operator_out570_out1 XOR Logical_Operator_out572_out1;

  Logical_Operator_out1083_out1 <= Logical_Operator_out58_out1 XOR Logical_Operator_out60_out1;

  Logical_Operator_out1084_out1 <= in116 XOR in120;

  Logical_Operator_out1085_out1 <= Logical_Operator_out573_out1 XOR Logical_Operator_out575_out1;

  Logical_Operator_out1086_out1 <= Logical_Operator_out574_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out1087_out1 <= Logical_Operator_out62_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out1088_out1 <= in124 XOR in128;

  Logical_Operator_out1089_out1 <= Logical_Operator_out577_out1 XOR Logical_Operator_out579_out1;

  Logical_Operator_out1090_out1 <= Logical_Operator_out578_out1 XOR Logical_Operator_out580_out1;

  Logical_Operator_out1091_out1 <= Logical_Operator_out66_out1 XOR Logical_Operator_out68_out1;

  Logical_Operator_out1092_out1 <= in132 XOR in136;

  Logical_Operator_out1093_out1 <= Logical_Operator_out581_out1 XOR Logical_Operator_out583_out1;

  Logical_Operator_out1094_out1 <= Logical_Operator_out582_out1 XOR Logical_Operator_out584_out1;

  Logical_Operator_out1095_out1 <= Logical_Operator_out70_out1 XOR Logical_Operator_out72_out1;

  Logical_Operator_out1096_out1 <= in140 XOR in144;

  Logical_Operator_out1097_out1 <= Logical_Operator_out585_out1 XOR Logical_Operator_out587_out1;

  Logical_Operator_out1098_out1 <= Logical_Operator_out586_out1 XOR Logical_Operator_out588_out1;

  Logical_Operator_out1099_out1 <= Logical_Operator_out74_out1 XOR Logical_Operator_out76_out1;

  Logical_Operator_out1100_out1 <= in148 XOR in152;

  Logical_Operator_out1101_out1 <= Logical_Operator_out589_out1 XOR Logical_Operator_out591_out1;

  Logical_Operator_out1102_out1 <= Logical_Operator_out590_out1 XOR Logical_Operator_out592_out1;

  Logical_Operator_out1103_out1 <= Logical_Operator_out78_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out1104_out1 <= in156 XOR in160;

  Logical_Operator_out1105_out1 <= Logical_Operator_out593_out1 XOR Logical_Operator_out595_out1;

  Logical_Operator_out1106_out1 <= Logical_Operator_out594_out1 XOR Logical_Operator_out596_out1;

  Logical_Operator_out1107_out1 <= Logical_Operator_out82_out1 XOR Logical_Operator_out84_out1;

  Logical_Operator_out1108_out1 <= in164 XOR in168;

  Logical_Operator_out1109_out1 <= Logical_Operator_out597_out1 XOR Logical_Operator_out599_out1;

  Logical_Operator_out1110_out1 <= Logical_Operator_out598_out1 XOR Logical_Operator_out600_out1;

  Logical_Operator_out1111_out1 <= Logical_Operator_out86_out1 XOR Logical_Operator_out88_out1;

  Logical_Operator_out1112_out1 <= in172 XOR in176;

  Logical_Operator_out1113_out1 <= Logical_Operator_out601_out1 XOR Logical_Operator_out603_out1;

  Logical_Operator_out1114_out1 <= Logical_Operator_out602_out1 XOR Logical_Operator_out604_out1;

  Logical_Operator_out1115_out1 <= Logical_Operator_out90_out1 XOR Logical_Operator_out92_out1;

  Logical_Operator_out1116_out1 <= in180 XOR in184;

  Logical_Operator_out1117_out1 <= Logical_Operator_out605_out1 XOR Logical_Operator_out607_out1;

  Logical_Operator_out1118_out1 <= Logical_Operator_out606_out1 XOR Logical_Operator_out608_out1;

  Logical_Operator_out1119_out1 <= Logical_Operator_out94_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out1120_out1 <= in188 XOR in192;

  Logical_Operator_out1121_out1 <= Logical_Operator_out609_out1 XOR Logical_Operator_out611_out1;

  Logical_Operator_out1122_out1 <= Logical_Operator_out610_out1 XOR Logical_Operator_out612_out1;

  Logical_Operator_out1123_out1 <= Logical_Operator_out98_out1 XOR Logical_Operator_out100_out1;

  Logical_Operator_out1124_out1 <= in196 XOR in200;

  Logical_Operator_out1125_out1 <= Logical_Operator_out613_out1 XOR Logical_Operator_out615_out1;

  Logical_Operator_out1126_out1 <= Logical_Operator_out614_out1 XOR Logical_Operator_out616_out1;

  Logical_Operator_out1127_out1 <= Logical_Operator_out102_out1 XOR Logical_Operator_out104_out1;

  Logical_Operator_out1128_out1 <= in204 XOR in208;

  Logical_Operator_out1129_out1 <= Logical_Operator_out617_out1 XOR Logical_Operator_out619_out1;

  Logical_Operator_out1130_out1 <= Logical_Operator_out618_out1 XOR Logical_Operator_out620_out1;

  Logical_Operator_out1131_out1 <= Logical_Operator_out106_out1 XOR Logical_Operator_out108_out1;

  Logical_Operator_out1132_out1 <= in212 XOR in216;

  Logical_Operator_out1133_out1 <= Logical_Operator_out621_out1 XOR Logical_Operator_out623_out1;

  Logical_Operator_out1134_out1 <= Logical_Operator_out622_out1 XOR Logical_Operator_out624_out1;

  Logical_Operator_out1135_out1 <= Logical_Operator_out110_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out1136_out1 <= in220 XOR in224;

  Logical_Operator_out1137_out1 <= Logical_Operator_out625_out1 XOR Logical_Operator_out627_out1;

  Logical_Operator_out1138_out1 <= Logical_Operator_out626_out1 XOR Logical_Operator_out628_out1;

  Logical_Operator_out1139_out1 <= Logical_Operator_out114_out1 XOR Logical_Operator_out116_out1;

  Logical_Operator_out1140_out1 <= in228 XOR in232;

  Logical_Operator_out1141_out1 <= Logical_Operator_out629_out1 XOR Logical_Operator_out631_out1;

  Logical_Operator_out1142_out1 <= Logical_Operator_out630_out1 XOR Logical_Operator_out632_out1;

  Logical_Operator_out1143_out1 <= Logical_Operator_out118_out1 XOR Logical_Operator_out120_out1;

  Logical_Operator_out1144_out1 <= in236 XOR in240;

  Logical_Operator_out1145_out1 <= Logical_Operator_out633_out1 XOR Logical_Operator_out635_out1;

  Logical_Operator_out1146_out1 <= Logical_Operator_out634_out1 XOR Logical_Operator_out636_out1;

  Logical_Operator_out1147_out1 <= Logical_Operator_out122_out1 XOR Logical_Operator_out124_out1;

  Logical_Operator_out1148_out1 <= in244 XOR in248;

  Logical_Operator_out1149_out1 <= Logical_Operator_out637_out1 XOR Logical_Operator_out639_out1;

  Logical_Operator_out1150_out1 <= Logical_Operator_out638_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out1151_out1 <= Logical_Operator_out126_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out1152_out1 <= in252 XOR in256;

  Logical_Operator_out1153_out1 <= Logical_Operator_out641_out1 XOR Logical_Operator_out643_out1;

  Logical_Operator_out1154_out1 <= Logical_Operator_out642_out1 XOR Logical_Operator_out644_out1;

  Logical_Operator_out1155_out1 <= Logical_Operator_out130_out1 XOR Logical_Operator_out132_out1;

  Logical_Operator_out1156_out1 <= in260 XOR in264;

  Logical_Operator_out1157_out1 <= Logical_Operator_out645_out1 XOR Logical_Operator_out647_out1;

  Logical_Operator_out1158_out1 <= Logical_Operator_out646_out1 XOR Logical_Operator_out648_out1;

  Logical_Operator_out1159_out1 <= Logical_Operator_out134_out1 XOR Logical_Operator_out136_out1;

  Logical_Operator_out1160_out1 <= in268 XOR in272;

  Logical_Operator_out1161_out1 <= Logical_Operator_out649_out1 XOR Logical_Operator_out651_out1;

  Logical_Operator_out1162_out1 <= Logical_Operator_out650_out1 XOR Logical_Operator_out652_out1;

  Logical_Operator_out1163_out1 <= Logical_Operator_out138_out1 XOR Logical_Operator_out140_out1;

  Logical_Operator_out1164_out1 <= in276 XOR in280;

  Logical_Operator_out1165_out1 <= Logical_Operator_out653_out1 XOR Logical_Operator_out655_out1;

  Logical_Operator_out1166_out1 <= Logical_Operator_out654_out1 XOR Logical_Operator_out656_out1;

  Logical_Operator_out1167_out1 <= Logical_Operator_out142_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out1168_out1 <= in284 XOR in288;

  Logical_Operator_out1169_out1 <= Logical_Operator_out657_out1 XOR Logical_Operator_out659_out1;

  Logical_Operator_out1170_out1 <= Logical_Operator_out658_out1 XOR Logical_Operator_out660_out1;

  Logical_Operator_out1171_out1 <= Logical_Operator_out146_out1 XOR Logical_Operator_out148_out1;

  Logical_Operator_out1172_out1 <= in292 XOR in296;

  Logical_Operator_out1173_out1 <= Logical_Operator_out661_out1 XOR Logical_Operator_out663_out1;

  Logical_Operator_out1174_out1 <= Logical_Operator_out662_out1 XOR Logical_Operator_out664_out1;

  Logical_Operator_out1175_out1 <= Logical_Operator_out150_out1 XOR Logical_Operator_out152_out1;

  Logical_Operator_out1176_out1 <= in300 XOR in304;

  Logical_Operator_out1177_out1 <= Logical_Operator_out665_out1 XOR Logical_Operator_out667_out1;

  Logical_Operator_out1178_out1 <= Logical_Operator_out666_out1 XOR Logical_Operator_out668_out1;

  Logical_Operator_out1179_out1 <= Logical_Operator_out154_out1 XOR Logical_Operator_out156_out1;

  Logical_Operator_out1180_out1 <= in308 XOR in312;

  Logical_Operator_out1181_out1 <= Logical_Operator_out669_out1 XOR Logical_Operator_out671_out1;

  Logical_Operator_out1182_out1 <= Logical_Operator_out670_out1 XOR Logical_Operator_out672_out1;

  Logical_Operator_out1183_out1 <= Logical_Operator_out158_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out1184_out1 <= in316 XOR in320;

  Logical_Operator_out1185_out1 <= Logical_Operator_out673_out1 XOR Logical_Operator_out675_out1;

  Logical_Operator_out1186_out1 <= Logical_Operator_out674_out1 XOR Logical_Operator_out676_out1;

  Logical_Operator_out1187_out1 <= Logical_Operator_out162_out1 XOR Logical_Operator_out164_out1;

  Logical_Operator_out1188_out1 <= in324 XOR in328;

  Logical_Operator_out1189_out1 <= Logical_Operator_out677_out1 XOR Logical_Operator_out679_out1;

  Logical_Operator_out1190_out1 <= Logical_Operator_out678_out1 XOR Logical_Operator_out680_out1;

  Logical_Operator_out1191_out1 <= Logical_Operator_out166_out1 XOR Logical_Operator_out168_out1;

  Logical_Operator_out1192_out1 <= in332 XOR in336;

  Logical_Operator_out1193_out1 <= Logical_Operator_out681_out1 XOR Logical_Operator_out683_out1;

  Logical_Operator_out1194_out1 <= Logical_Operator_out682_out1 XOR Logical_Operator_out684_out1;

  Logical_Operator_out1195_out1 <= Logical_Operator_out170_out1 XOR Logical_Operator_out172_out1;

  Logical_Operator_out1196_out1 <= in340 XOR in344;

  Logical_Operator_out1197_out1 <= Logical_Operator_out685_out1 XOR Logical_Operator_out687_out1;

  Logical_Operator_out1198_out1 <= Logical_Operator_out686_out1 XOR Logical_Operator_out688_out1;

  Logical_Operator_out1199_out1 <= Logical_Operator_out174_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out1200_out1 <= in348 XOR in352;

  Logical_Operator_out1201_out1 <= Logical_Operator_out689_out1 XOR Logical_Operator_out691_out1;

  Logical_Operator_out1202_out1 <= Logical_Operator_out690_out1 XOR Logical_Operator_out692_out1;

  Logical_Operator_out1203_out1 <= Logical_Operator_out178_out1 XOR Logical_Operator_out180_out1;

  Logical_Operator_out1204_out1 <= in356 XOR in360;

  Logical_Operator_out1205_out1 <= Logical_Operator_out693_out1 XOR Logical_Operator_out695_out1;

  Logical_Operator_out1206_out1 <= Logical_Operator_out694_out1 XOR Logical_Operator_out696_out1;

  Logical_Operator_out1207_out1 <= Logical_Operator_out182_out1 XOR Logical_Operator_out184_out1;

  Logical_Operator_out1208_out1 <= in364 XOR in368;

  Logical_Operator_out1209_out1 <= Logical_Operator_out697_out1 XOR Logical_Operator_out699_out1;

  Logical_Operator_out1210_out1 <= Logical_Operator_out698_out1 XOR Logical_Operator_out700_out1;

  Logical_Operator_out1211_out1 <= Logical_Operator_out186_out1 XOR Logical_Operator_out188_out1;

  Logical_Operator_out1212_out1 <= in372 XOR in376;

  Logical_Operator_out1213_out1 <= Logical_Operator_out701_out1 XOR Logical_Operator_out703_out1;

  Logical_Operator_out1214_out1 <= Logical_Operator_out702_out1 XOR Logical_Operator_out704_out1;

  Logical_Operator_out1215_out1 <= Logical_Operator_out190_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out1216_out1 <= in380 XOR in384;

  Logical_Operator_out1217_out1 <= Logical_Operator_out705_out1 XOR Logical_Operator_out707_out1;

  Logical_Operator_out1218_out1 <= Logical_Operator_out706_out1 XOR Logical_Operator_out708_out1;

  Logical_Operator_out1219_out1 <= Logical_Operator_out194_out1 XOR Logical_Operator_out196_out1;

  Logical_Operator_out1220_out1 <= in388 XOR in392;

  Logical_Operator_out1221_out1 <= Logical_Operator_out709_out1 XOR Logical_Operator_out711_out1;

  Logical_Operator_out1222_out1 <= Logical_Operator_out710_out1 XOR Logical_Operator_out712_out1;

  Logical_Operator_out1223_out1 <= Logical_Operator_out198_out1 XOR Logical_Operator_out200_out1;

  Logical_Operator_out1224_out1 <= in396 XOR in400;

  Logical_Operator_out1225_out1 <= Logical_Operator_out713_out1 XOR Logical_Operator_out715_out1;

  Logical_Operator_out1226_out1 <= Logical_Operator_out714_out1 XOR Logical_Operator_out716_out1;

  Logical_Operator_out1227_out1 <= Logical_Operator_out202_out1 XOR Logical_Operator_out204_out1;

  Logical_Operator_out1228_out1 <= in404 XOR in408;

  Logical_Operator_out1229_out1 <= Logical_Operator_out717_out1 XOR Logical_Operator_out719_out1;

  Logical_Operator_out1230_out1 <= Logical_Operator_out718_out1 XOR Logical_Operator_out720_out1;

  Logical_Operator_out1231_out1 <= Logical_Operator_out206_out1 XOR Logical_Operator_out208_out1;

  Logical_Operator_out1232_out1 <= in412 XOR in416;

  Logical_Operator_out1233_out1 <= Logical_Operator_out721_out1 XOR Logical_Operator_out723_out1;

  Logical_Operator_out1234_out1 <= Logical_Operator_out722_out1 XOR Logical_Operator_out724_out1;

  Logical_Operator_out1235_out1 <= Logical_Operator_out210_out1 XOR Logical_Operator_out212_out1;

  Logical_Operator_out1236_out1 <= in420 XOR in424;

  Logical_Operator_out1237_out1 <= Logical_Operator_out725_out1 XOR Logical_Operator_out727_out1;

  Logical_Operator_out1238_out1 <= Logical_Operator_out726_out1 XOR Logical_Operator_out728_out1;

  Logical_Operator_out1239_out1 <= Logical_Operator_out214_out1 XOR Logical_Operator_out216_out1;

  Logical_Operator_out1240_out1 <= in428 XOR in432;

  Logical_Operator_out1241_out1 <= Logical_Operator_out729_out1 XOR Logical_Operator_out731_out1;

  Logical_Operator_out1242_out1 <= Logical_Operator_out730_out1 XOR Logical_Operator_out732_out1;

  Logical_Operator_out1243_out1 <= Logical_Operator_out218_out1 XOR Logical_Operator_out220_out1;

  Logical_Operator_out1244_out1 <= in436 XOR in440;

  Logical_Operator_out1245_out1 <= Logical_Operator_out733_out1 XOR Logical_Operator_out735_out1;

  Logical_Operator_out1246_out1 <= Logical_Operator_out734_out1 XOR Logical_Operator_out736_out1;

  Logical_Operator_out1247_out1 <= Logical_Operator_out222_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out1248_out1 <= in444 XOR in448;

  Logical_Operator_out1249_out1 <= Logical_Operator_out737_out1 XOR Logical_Operator_out739_out1;

  Logical_Operator_out1250_out1 <= Logical_Operator_out738_out1 XOR Logical_Operator_out740_out1;

  Logical_Operator_out1251_out1 <= Logical_Operator_out226_out1 XOR Logical_Operator_out228_out1;

  Logical_Operator_out1252_out1 <= in452 XOR in456;

  Logical_Operator_out1253_out1 <= Logical_Operator_out741_out1 XOR Logical_Operator_out743_out1;

  Logical_Operator_out1254_out1 <= Logical_Operator_out742_out1 XOR Logical_Operator_out744_out1;

  Logical_Operator_out1255_out1 <= Logical_Operator_out230_out1 XOR Logical_Operator_out232_out1;

  Logical_Operator_out1256_out1 <= in460 XOR in464;

  Logical_Operator_out1257_out1 <= Logical_Operator_out745_out1 XOR Logical_Operator_out747_out1;

  Logical_Operator_out1258_out1 <= Logical_Operator_out746_out1 XOR Logical_Operator_out748_out1;

  Logical_Operator_out1259_out1 <= Logical_Operator_out234_out1 XOR Logical_Operator_out236_out1;

  Logical_Operator_out1260_out1 <= in468 XOR in472;

  Logical_Operator_out1261_out1 <= Logical_Operator_out749_out1 XOR Logical_Operator_out751_out1;

  Logical_Operator_out1262_out1 <= Logical_Operator_out750_out1 XOR Logical_Operator_out752_out1;

  Logical_Operator_out1263_out1 <= Logical_Operator_out238_out1 XOR Logical_Operator_out240_out1;

  Logical_Operator_out1264_out1 <= in476 XOR in480;

  Logical_Operator_out1265_out1 <= Logical_Operator_out753_out1 XOR Logical_Operator_out755_out1;

  Logical_Operator_out1266_out1 <= Logical_Operator_out754_out1 XOR Logical_Operator_out756_out1;

  Logical_Operator_out1267_out1 <= Logical_Operator_out242_out1 XOR Logical_Operator_out244_out1;

  Logical_Operator_out1268_out1 <= in484 XOR in488;

  Logical_Operator_out1269_out1 <= Logical_Operator_out757_out1 XOR Logical_Operator_out759_out1;

  Logical_Operator_out1270_out1 <= Logical_Operator_out758_out1 XOR Logical_Operator_out760_out1;

  Logical_Operator_out1271_out1 <= Logical_Operator_out246_out1 XOR Logical_Operator_out248_out1;

  Logical_Operator_out1272_out1 <= in492 XOR in496;

  Logical_Operator_out1273_out1 <= Logical_Operator_out761_out1 XOR Logical_Operator_out763_out1;

  Logical_Operator_out1274_out1 <= Logical_Operator_out762_out1 XOR Logical_Operator_out764_out1;

  Logical_Operator_out1275_out1 <= Logical_Operator_out250_out1 XOR Logical_Operator_out252_out1;

  Logical_Operator_out1276_out1 <= in500 XOR in504;

  Logical_Operator_out1277_out1 <= Logical_Operator_out765_out1 XOR Logical_Operator_out767_out1;

  Logical_Operator_out1278_out1 <= Logical_Operator_out766_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out1279_out1 <= Logical_Operator_out254_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out1280_out1 <= in508 XOR in512;

  Logical_Operator_out1281_out1 <= Logical_Operator_out769_out1 XOR Logical_Operator_out771_out1;

  Logical_Operator_out1282_out1 <= Logical_Operator_out770_out1 XOR Logical_Operator_out772_out1;

  Logical_Operator_out1283_out1 <= Logical_Operator_out258_out1 XOR Logical_Operator_out260_out1;

  Logical_Operator_out1284_out1 <= in516 XOR in520;

  Logical_Operator_out1285_out1 <= Logical_Operator_out773_out1 XOR Logical_Operator_out775_out1;

  Logical_Operator_out1286_out1 <= Logical_Operator_out774_out1 XOR Logical_Operator_out776_out1;

  Logical_Operator_out1287_out1 <= Logical_Operator_out262_out1 XOR Logical_Operator_out264_out1;

  Logical_Operator_out1288_out1 <= in524 XOR in528;

  Logical_Operator_out1289_out1 <= Logical_Operator_out777_out1 XOR Logical_Operator_out779_out1;

  Logical_Operator_out1290_out1 <= Logical_Operator_out778_out1 XOR Logical_Operator_out780_out1;

  Logical_Operator_out1291_out1 <= Logical_Operator_out266_out1 XOR Logical_Operator_out268_out1;

  Logical_Operator_out1292_out1 <= in532 XOR in536;

  Logical_Operator_out1293_out1 <= Logical_Operator_out781_out1 XOR Logical_Operator_out783_out1;

  Logical_Operator_out1294_out1 <= Logical_Operator_out782_out1 XOR Logical_Operator_out784_out1;

  Logical_Operator_out1295_out1 <= Logical_Operator_out270_out1 XOR Logical_Operator_out272_out1;

  Logical_Operator_out1296_out1 <= in540 XOR in544;

  Logical_Operator_out1297_out1 <= Logical_Operator_out785_out1 XOR Logical_Operator_out787_out1;

  Logical_Operator_out1298_out1 <= Logical_Operator_out786_out1 XOR Logical_Operator_out788_out1;

  Logical_Operator_out1299_out1 <= Logical_Operator_out274_out1 XOR Logical_Operator_out276_out1;

  Logical_Operator_out1300_out1 <= in548 XOR in552;

  Logical_Operator_out1301_out1 <= Logical_Operator_out789_out1 XOR Logical_Operator_out791_out1;

  Logical_Operator_out1302_out1 <= Logical_Operator_out790_out1 XOR Logical_Operator_out792_out1;

  Logical_Operator_out1303_out1 <= Logical_Operator_out278_out1 XOR Logical_Operator_out280_out1;

  Logical_Operator_out1304_out1 <= in556 XOR in560;

  Logical_Operator_out1305_out1 <= Logical_Operator_out793_out1 XOR Logical_Operator_out795_out1;

  Logical_Operator_out1306_out1 <= Logical_Operator_out794_out1 XOR Logical_Operator_out796_out1;

  Logical_Operator_out1307_out1 <= Logical_Operator_out282_out1 XOR Logical_Operator_out284_out1;

  Logical_Operator_out1308_out1 <= in564 XOR in568;

  Logical_Operator_out1309_out1 <= Logical_Operator_out797_out1 XOR Logical_Operator_out799_out1;

  Logical_Operator_out1310_out1 <= Logical_Operator_out798_out1 XOR Logical_Operator_out800_out1;

  Logical_Operator_out1311_out1 <= Logical_Operator_out286_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out1312_out1 <= in572 XOR in576;

  Logical_Operator_out1313_out1 <= Logical_Operator_out801_out1 XOR Logical_Operator_out803_out1;

  Logical_Operator_out1314_out1 <= Logical_Operator_out802_out1 XOR Logical_Operator_out804_out1;

  Logical_Operator_out1315_out1 <= Logical_Operator_out290_out1 XOR Logical_Operator_out292_out1;

  Logical_Operator_out1316_out1 <= in580 XOR in584;

  Logical_Operator_out1317_out1 <= Logical_Operator_out805_out1 XOR Logical_Operator_out807_out1;

  Logical_Operator_out1318_out1 <= Logical_Operator_out806_out1 XOR Logical_Operator_out808_out1;

  Logical_Operator_out1319_out1 <= Logical_Operator_out294_out1 XOR Logical_Operator_out296_out1;

  Logical_Operator_out1320_out1 <= in588 XOR in592;

  Logical_Operator_out1321_out1 <= Logical_Operator_out809_out1 XOR Logical_Operator_out811_out1;

  Logical_Operator_out1322_out1 <= Logical_Operator_out810_out1 XOR Logical_Operator_out812_out1;

  Logical_Operator_out1323_out1 <= Logical_Operator_out298_out1 XOR Logical_Operator_out300_out1;

  Logical_Operator_out1324_out1 <= in596 XOR in600;

  Logical_Operator_out1325_out1 <= Logical_Operator_out813_out1 XOR Logical_Operator_out815_out1;

  Logical_Operator_out1326_out1 <= Logical_Operator_out814_out1 XOR Logical_Operator_out816_out1;

  Logical_Operator_out1327_out1 <= Logical_Operator_out302_out1 XOR Logical_Operator_out304_out1;

  Logical_Operator_out1328_out1 <= in604 XOR in608;

  Logical_Operator_out1329_out1 <= Logical_Operator_out817_out1 XOR Logical_Operator_out819_out1;

  Logical_Operator_out1330_out1 <= Logical_Operator_out818_out1 XOR Logical_Operator_out820_out1;

  Logical_Operator_out1331_out1 <= Logical_Operator_out306_out1 XOR Logical_Operator_out308_out1;

  Logical_Operator_out1332_out1 <= in612 XOR in616;

  Logical_Operator_out1333_out1 <= Logical_Operator_out821_out1 XOR Logical_Operator_out823_out1;

  Logical_Operator_out1334_out1 <= Logical_Operator_out822_out1 XOR Logical_Operator_out824_out1;

  Logical_Operator_out1335_out1 <= Logical_Operator_out310_out1 XOR Logical_Operator_out312_out1;

  Logical_Operator_out1336_out1 <= in620 XOR in624;

  Logical_Operator_out1337_out1 <= Logical_Operator_out825_out1 XOR Logical_Operator_out827_out1;

  Logical_Operator_out1338_out1 <= Logical_Operator_out826_out1 XOR Logical_Operator_out828_out1;

  Logical_Operator_out1339_out1 <= Logical_Operator_out314_out1 XOR Logical_Operator_out316_out1;

  Logical_Operator_out1340_out1 <= in628 XOR in632;

  Logical_Operator_out1341_out1 <= Logical_Operator_out829_out1 XOR Logical_Operator_out831_out1;

  Logical_Operator_out1342_out1 <= Logical_Operator_out830_out1 XOR Logical_Operator_out832_out1;

  Logical_Operator_out1343_out1 <= Logical_Operator_out318_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out1344_out1 <= in636 XOR in640;

  Logical_Operator_out1345_out1 <= Logical_Operator_out833_out1 XOR Logical_Operator_out835_out1;

  Logical_Operator_out1346_out1 <= Logical_Operator_out834_out1 XOR Logical_Operator_out836_out1;

  Logical_Operator_out1347_out1 <= Logical_Operator_out322_out1 XOR Logical_Operator_out324_out1;

  Logical_Operator_out1348_out1 <= in644 XOR in648;

  Logical_Operator_out1349_out1 <= Logical_Operator_out837_out1 XOR Logical_Operator_out839_out1;

  Logical_Operator_out1350_out1 <= Logical_Operator_out838_out1 XOR Logical_Operator_out840_out1;

  Logical_Operator_out1351_out1 <= Logical_Operator_out326_out1 XOR Logical_Operator_out328_out1;

  Logical_Operator_out1352_out1 <= in652 XOR in656;

  Logical_Operator_out1353_out1 <= Logical_Operator_out841_out1 XOR Logical_Operator_out843_out1;

  Logical_Operator_out1354_out1 <= Logical_Operator_out842_out1 XOR Logical_Operator_out844_out1;

  Logical_Operator_out1355_out1 <= Logical_Operator_out330_out1 XOR Logical_Operator_out332_out1;

  Logical_Operator_out1356_out1 <= in660 XOR in664;

  Logical_Operator_out1357_out1 <= Logical_Operator_out845_out1 XOR Logical_Operator_out847_out1;

  Logical_Operator_out1358_out1 <= Logical_Operator_out846_out1 XOR Logical_Operator_out848_out1;

  Logical_Operator_out1359_out1 <= Logical_Operator_out334_out1 XOR Logical_Operator_out336_out1;

  Logical_Operator_out1360_out1 <= in668 XOR in672;

  Logical_Operator_out1361_out1 <= Logical_Operator_out849_out1 XOR Logical_Operator_out851_out1;

  Logical_Operator_out1362_out1 <= Logical_Operator_out850_out1 XOR Logical_Operator_out852_out1;

  Logical_Operator_out1363_out1 <= Logical_Operator_out338_out1 XOR Logical_Operator_out340_out1;

  Logical_Operator_out1364_out1 <= in676 XOR in680;

  Logical_Operator_out1365_out1 <= Logical_Operator_out853_out1 XOR Logical_Operator_out855_out1;

  Logical_Operator_out1366_out1 <= Logical_Operator_out854_out1 XOR Logical_Operator_out856_out1;

  Logical_Operator_out1367_out1 <= Logical_Operator_out342_out1 XOR Logical_Operator_out344_out1;

  Logical_Operator_out1368_out1 <= in684 XOR in688;

  Logical_Operator_out1369_out1 <= Logical_Operator_out857_out1 XOR Logical_Operator_out859_out1;

  Logical_Operator_out1370_out1 <= Logical_Operator_out858_out1 XOR Logical_Operator_out860_out1;

  Logical_Operator_out1371_out1 <= Logical_Operator_out346_out1 XOR Logical_Operator_out348_out1;

  Logical_Operator_out1372_out1 <= in692 XOR in696;

  Logical_Operator_out1373_out1 <= Logical_Operator_out861_out1 XOR Logical_Operator_out863_out1;

  Logical_Operator_out1374_out1 <= Logical_Operator_out862_out1 XOR Logical_Operator_out864_out1;

  Logical_Operator_out1375_out1 <= Logical_Operator_out350_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out1376_out1 <= in700 XOR in704;

  Logical_Operator_out1377_out1 <= Logical_Operator_out865_out1 XOR Logical_Operator_out867_out1;

  Logical_Operator_out1378_out1 <= Logical_Operator_out866_out1 XOR Logical_Operator_out868_out1;

  Logical_Operator_out1379_out1 <= Logical_Operator_out354_out1 XOR Logical_Operator_out356_out1;

  Logical_Operator_out1380_out1 <= in708 XOR in712;

  Logical_Operator_out1381_out1 <= Logical_Operator_out869_out1 XOR Logical_Operator_out871_out1;

  Logical_Operator_out1382_out1 <= Logical_Operator_out870_out1 XOR Logical_Operator_out872_out1;

  Logical_Operator_out1383_out1 <= Logical_Operator_out358_out1 XOR Logical_Operator_out360_out1;

  Logical_Operator_out1384_out1 <= in716 XOR in720;

  Logical_Operator_out1385_out1 <= Logical_Operator_out873_out1 XOR Logical_Operator_out875_out1;

  Logical_Operator_out1386_out1 <= Logical_Operator_out874_out1 XOR Logical_Operator_out876_out1;

  Logical_Operator_out1387_out1 <= Logical_Operator_out362_out1 XOR Logical_Operator_out364_out1;

  Logical_Operator_out1388_out1 <= in724 XOR in728;

  Logical_Operator_out1389_out1 <= Logical_Operator_out877_out1 XOR Logical_Operator_out879_out1;

  Logical_Operator_out1390_out1 <= Logical_Operator_out878_out1 XOR Logical_Operator_out880_out1;

  Logical_Operator_out1391_out1 <= Logical_Operator_out366_out1 XOR Logical_Operator_out368_out1;

  Logical_Operator_out1392_out1 <= in732 XOR in736;

  Logical_Operator_out1393_out1 <= Logical_Operator_out881_out1 XOR Logical_Operator_out883_out1;

  Logical_Operator_out1394_out1 <= Logical_Operator_out882_out1 XOR Logical_Operator_out884_out1;

  Logical_Operator_out1395_out1 <= Logical_Operator_out370_out1 XOR Logical_Operator_out372_out1;

  Logical_Operator_out1396_out1 <= in740 XOR in744;

  Logical_Operator_out1397_out1 <= Logical_Operator_out885_out1 XOR Logical_Operator_out887_out1;

  Logical_Operator_out1398_out1 <= Logical_Operator_out886_out1 XOR Logical_Operator_out888_out1;

  Logical_Operator_out1399_out1 <= Logical_Operator_out374_out1 XOR Logical_Operator_out376_out1;

  Logical_Operator_out1400_out1 <= in748 XOR in752;

  Logical_Operator_out1401_out1 <= Logical_Operator_out889_out1 XOR Logical_Operator_out891_out1;

  Logical_Operator_out1402_out1 <= Logical_Operator_out890_out1 XOR Logical_Operator_out892_out1;

  Logical_Operator_out1403_out1 <= Logical_Operator_out378_out1 XOR Logical_Operator_out380_out1;

  Logical_Operator_out1404_out1 <= in756 XOR in760;

  Logical_Operator_out1405_out1 <= Logical_Operator_out893_out1 XOR Logical_Operator_out895_out1;

  Logical_Operator_out1406_out1 <= Logical_Operator_out894_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out1407_out1 <= Logical_Operator_out382_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out1408_out1 <= in764 XOR in768;

  Logical_Operator_out1409_out1 <= Logical_Operator_out897_out1 XOR Logical_Operator_out899_out1;

  Logical_Operator_out1410_out1 <= Logical_Operator_out898_out1 XOR Logical_Operator_out900_out1;

  Logical_Operator_out1411_out1 <= Logical_Operator_out386_out1 XOR Logical_Operator_out388_out1;

  Logical_Operator_out1412_out1 <= in772 XOR in776;

  Logical_Operator_out1413_out1 <= Logical_Operator_out901_out1 XOR Logical_Operator_out903_out1;

  Logical_Operator_out1414_out1 <= Logical_Operator_out902_out1 XOR Logical_Operator_out904_out1;

  Logical_Operator_out1415_out1 <= Logical_Operator_out390_out1 XOR Logical_Operator_out392_out1;

  Logical_Operator_out1416_out1 <= in780 XOR in784;

  Logical_Operator_out1417_out1 <= Logical_Operator_out905_out1 XOR Logical_Operator_out907_out1;

  Logical_Operator_out1418_out1 <= Logical_Operator_out906_out1 XOR Logical_Operator_out908_out1;

  Logical_Operator_out1419_out1 <= Logical_Operator_out394_out1 XOR Logical_Operator_out396_out1;

  Logical_Operator_out1420_out1 <= in788 XOR in792;

  Logical_Operator_out1421_out1 <= Logical_Operator_out909_out1 XOR Logical_Operator_out911_out1;

  Logical_Operator_out1422_out1 <= Logical_Operator_out910_out1 XOR Logical_Operator_out912_out1;

  Logical_Operator_out1423_out1 <= Logical_Operator_out398_out1 XOR Logical_Operator_out400_out1;

  Logical_Operator_out1424_out1 <= in796 XOR in800;

  Logical_Operator_out1425_out1 <= Logical_Operator_out913_out1 XOR Logical_Operator_out915_out1;

  Logical_Operator_out1426_out1 <= Logical_Operator_out914_out1 XOR Logical_Operator_out916_out1;

  Logical_Operator_out1427_out1 <= Logical_Operator_out402_out1 XOR Logical_Operator_out404_out1;

  Logical_Operator_out1428_out1 <= in804 XOR in808;

  Logical_Operator_out1429_out1 <= Logical_Operator_out917_out1 XOR Logical_Operator_out919_out1;

  Logical_Operator_out1430_out1 <= Logical_Operator_out918_out1 XOR Logical_Operator_out920_out1;

  Logical_Operator_out1431_out1 <= Logical_Operator_out406_out1 XOR Logical_Operator_out408_out1;

  Logical_Operator_out1432_out1 <= in812 XOR in816;

  Logical_Operator_out1433_out1 <= Logical_Operator_out921_out1 XOR Logical_Operator_out923_out1;

  Logical_Operator_out1434_out1 <= Logical_Operator_out922_out1 XOR Logical_Operator_out924_out1;

  Logical_Operator_out1435_out1 <= Logical_Operator_out410_out1 XOR Logical_Operator_out412_out1;

  Logical_Operator_out1436_out1 <= in820 XOR in824;

  Logical_Operator_out1437_out1 <= Logical_Operator_out925_out1 XOR Logical_Operator_out927_out1;

  Logical_Operator_out1438_out1 <= Logical_Operator_out926_out1 XOR Logical_Operator_out928_out1;

  Logical_Operator_out1439_out1 <= Logical_Operator_out414_out1 XOR Logical_Operator_out416_out1;

  Logical_Operator_out1440_out1 <= in828 XOR in832;

  Logical_Operator_out1441_out1 <= Logical_Operator_out929_out1 XOR Logical_Operator_out931_out1;

  Logical_Operator_out1442_out1 <= Logical_Operator_out930_out1 XOR Logical_Operator_out932_out1;

  Logical_Operator_out1443_out1 <= Logical_Operator_out418_out1 XOR Logical_Operator_out420_out1;

  Logical_Operator_out1444_out1 <= in836 XOR in840;

  Logical_Operator_out1445_out1 <= Logical_Operator_out933_out1 XOR Logical_Operator_out935_out1;

  Logical_Operator_out1446_out1 <= Logical_Operator_out934_out1 XOR Logical_Operator_out936_out1;

  Logical_Operator_out1447_out1 <= Logical_Operator_out422_out1 XOR Logical_Operator_out424_out1;

  Logical_Operator_out1448_out1 <= in844 XOR in848;

  Logical_Operator_out1449_out1 <= Logical_Operator_out937_out1 XOR Logical_Operator_out939_out1;

  Logical_Operator_out1450_out1 <= Logical_Operator_out938_out1 XOR Logical_Operator_out940_out1;

  Logical_Operator_out1451_out1 <= Logical_Operator_out426_out1 XOR Logical_Operator_out428_out1;

  Logical_Operator_out1452_out1 <= in852 XOR in856;

  Logical_Operator_out1453_out1 <= Logical_Operator_out941_out1 XOR Logical_Operator_out943_out1;

  Logical_Operator_out1454_out1 <= Logical_Operator_out942_out1 XOR Logical_Operator_out944_out1;

  Logical_Operator_out1455_out1 <= Logical_Operator_out430_out1 XOR Logical_Operator_out432_out1;

  Logical_Operator_out1456_out1 <= in860 XOR in864;

  Logical_Operator_out1457_out1 <= Logical_Operator_out945_out1 XOR Logical_Operator_out947_out1;

  Logical_Operator_out1458_out1 <= Logical_Operator_out946_out1 XOR Logical_Operator_out948_out1;

  Logical_Operator_out1459_out1 <= Logical_Operator_out434_out1 XOR Logical_Operator_out436_out1;

  Logical_Operator_out1460_out1 <= in868 XOR in872;

  Logical_Operator_out1461_out1 <= Logical_Operator_out949_out1 XOR Logical_Operator_out951_out1;

  Logical_Operator_out1462_out1 <= Logical_Operator_out950_out1 XOR Logical_Operator_out952_out1;

  Logical_Operator_out1463_out1 <= Logical_Operator_out438_out1 XOR Logical_Operator_out440_out1;

  Logical_Operator_out1464_out1 <= in876 XOR in880;

  Logical_Operator_out1465_out1 <= Logical_Operator_out953_out1 XOR Logical_Operator_out955_out1;

  Logical_Operator_out1466_out1 <= Logical_Operator_out954_out1 XOR Logical_Operator_out956_out1;

  Logical_Operator_out1467_out1 <= Logical_Operator_out442_out1 XOR Logical_Operator_out444_out1;

  Logical_Operator_out1468_out1 <= in884 XOR in888;

  Logical_Operator_out1469_out1 <= Logical_Operator_out957_out1 XOR Logical_Operator_out959_out1;

  Logical_Operator_out1470_out1 <= Logical_Operator_out958_out1 XOR Logical_Operator_out960_out1;

  Logical_Operator_out1471_out1 <= Logical_Operator_out446_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out1472_out1 <= in892 XOR in896;

  Logical_Operator_out1473_out1 <= Logical_Operator_out961_out1 XOR Logical_Operator_out963_out1;

  Logical_Operator_out1474_out1 <= Logical_Operator_out962_out1 XOR Logical_Operator_out964_out1;

  Logical_Operator_out1475_out1 <= Logical_Operator_out450_out1 XOR Logical_Operator_out452_out1;

  Logical_Operator_out1476_out1 <= in900 XOR in904;

  Logical_Operator_out1477_out1 <= Logical_Operator_out965_out1 XOR Logical_Operator_out967_out1;

  Logical_Operator_out1478_out1 <= Logical_Operator_out966_out1 XOR Logical_Operator_out968_out1;

  Logical_Operator_out1479_out1 <= Logical_Operator_out454_out1 XOR Logical_Operator_out456_out1;

  Logical_Operator_out1480_out1 <= in908 XOR in912;

  Logical_Operator_out1481_out1 <= Logical_Operator_out969_out1 XOR Logical_Operator_out971_out1;

  Logical_Operator_out1482_out1 <= Logical_Operator_out970_out1 XOR Logical_Operator_out972_out1;

  Logical_Operator_out1483_out1 <= Logical_Operator_out458_out1 XOR Logical_Operator_out460_out1;

  Logical_Operator_out1484_out1 <= in916 XOR in920;

  Logical_Operator_out1485_out1 <= Logical_Operator_out973_out1 XOR Logical_Operator_out975_out1;

  Logical_Operator_out1486_out1 <= Logical_Operator_out974_out1 XOR Logical_Operator_out976_out1;

  Logical_Operator_out1487_out1 <= Logical_Operator_out462_out1 XOR Logical_Operator_out464_out1;

  Logical_Operator_out1488_out1 <= in924 XOR in928;

  Logical_Operator_out1489_out1 <= Logical_Operator_out977_out1 XOR Logical_Operator_out979_out1;

  Logical_Operator_out1490_out1 <= Logical_Operator_out978_out1 XOR Logical_Operator_out980_out1;

  Logical_Operator_out1491_out1 <= Logical_Operator_out466_out1 XOR Logical_Operator_out468_out1;

  Logical_Operator_out1492_out1 <= in932 XOR in936;

  Logical_Operator_out1493_out1 <= Logical_Operator_out981_out1 XOR Logical_Operator_out983_out1;

  Logical_Operator_out1494_out1 <= Logical_Operator_out982_out1 XOR Logical_Operator_out984_out1;

  Logical_Operator_out1495_out1 <= Logical_Operator_out470_out1 XOR Logical_Operator_out472_out1;

  Logical_Operator_out1496_out1 <= in940 XOR in944;

  Logical_Operator_out1497_out1 <= Logical_Operator_out985_out1 XOR Logical_Operator_out987_out1;

  Logical_Operator_out1498_out1 <= Logical_Operator_out986_out1 XOR Logical_Operator_out988_out1;

  Logical_Operator_out1499_out1 <= Logical_Operator_out474_out1 XOR Logical_Operator_out476_out1;

  Logical_Operator_out1500_out1 <= in948 XOR in952;

  Logical_Operator_out1501_out1 <= Logical_Operator_out989_out1 XOR Logical_Operator_out991_out1;

  Logical_Operator_out1502_out1 <= Logical_Operator_out990_out1 XOR Logical_Operator_out992_out1;

  Logical_Operator_out1503_out1 <= Logical_Operator_out478_out1 XOR Logical_Operator_out480_out1;

  Logical_Operator_out1504_out1 <= in956 XOR in960;

  Logical_Operator_out1505_out1 <= Logical_Operator_out993_out1 XOR Logical_Operator_out995_out1;

  Logical_Operator_out1506_out1 <= Logical_Operator_out994_out1 XOR Logical_Operator_out996_out1;

  Logical_Operator_out1507_out1 <= Logical_Operator_out482_out1 XOR Logical_Operator_out484_out1;

  Logical_Operator_out1508_out1 <= in964 XOR in968;

  Logical_Operator_out1509_out1 <= Logical_Operator_out997_out1 XOR Logical_Operator_out999_out1;

  Logical_Operator_out1510_out1 <= Logical_Operator_out998_out1 XOR Logical_Operator_out1000_out1;

  Logical_Operator_out1511_out1 <= Logical_Operator_out486_out1 XOR Logical_Operator_out488_out1;

  Logical_Operator_out1512_out1 <= in972 XOR in976;

  Logical_Operator_out1513_out1 <= Logical_Operator_out1001_out1 XOR Logical_Operator_out1003_out1;

  Logical_Operator_out1514_out1 <= Logical_Operator_out1002_out1 XOR Logical_Operator_out1004_out1;

  Logical_Operator_out1515_out1 <= Logical_Operator_out490_out1 XOR Logical_Operator_out492_out1;

  Logical_Operator_out1516_out1 <= in980 XOR in984;

  Logical_Operator_out1517_out1 <= Logical_Operator_out1005_out1 XOR Logical_Operator_out1007_out1;

  Logical_Operator_out1518_out1 <= Logical_Operator_out1006_out1 XOR Logical_Operator_out1008_out1;

  Logical_Operator_out1519_out1 <= Logical_Operator_out494_out1 XOR Logical_Operator_out496_out1;

  Logical_Operator_out1520_out1 <= in988 XOR in992;

  Logical_Operator_out1521_out1 <= Logical_Operator_out1009_out1 XOR Logical_Operator_out1011_out1;

  Logical_Operator_out1522_out1 <= Logical_Operator_out1010_out1 XOR Logical_Operator_out1012_out1;

  Logical_Operator_out1523_out1 <= Logical_Operator_out498_out1 XOR Logical_Operator_out500_out1;

  Logical_Operator_out1524_out1 <= in996 XOR in1000;

  Logical_Operator_out1525_out1 <= Logical_Operator_out1013_out1 XOR Logical_Operator_out1015_out1;

  Logical_Operator_out1526_out1 <= Logical_Operator_out1014_out1 XOR Logical_Operator_out1016_out1;

  Logical_Operator_out1527_out1 <= Logical_Operator_out502_out1 XOR Logical_Operator_out504_out1;

  Logical_Operator_out1528_out1 <= in1004 XOR in1008;

  Logical_Operator_out1529_out1 <= Logical_Operator_out1017_out1 XOR Logical_Operator_out1019_out1;

  Logical_Operator_out1530_out1 <= Logical_Operator_out1018_out1 XOR Logical_Operator_out1020_out1;

  Logical_Operator_out1531_out1 <= Logical_Operator_out506_out1 XOR Logical_Operator_out508_out1;

  Logical_Operator_out1532_out1 <= in1012 XOR in1016;

  Logical_Operator_out1533_out1 <= Logical_Operator_out1021_out1 XOR Logical_Operator_out1023_out1;

  Logical_Operator_out1534_out1 <= Logical_Operator_out1022_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out1535_out1 <= Logical_Operator_out510_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out1536_out1 <= in1020 XOR in1024;

  Logical_Operator_out1537_out1 <= Logical_Operator_out1025_out1 XOR Logical_Operator_out1029_out1;

  Logical_Operator_out1538_out1 <= Logical_Operator_out1026_out1 XOR Logical_Operator_out1030_out1;

  Logical_Operator_out1539_out1 <= Logical_Operator_out1027_out1 XOR Logical_Operator_out1031_out1;

  Logical_Operator_out1540_out1 <= Logical_Operator_out1028_out1 XOR Logical_Operator_out1032_out1;

  Logical_Operator_out1541_out1 <= Logical_Operator_out515_out1 XOR Logical_Operator_out519_out1;

  Logical_Operator_out1542_out1 <= Logical_Operator_out516_out1 XOR Logical_Operator_out520_out1;

  Logical_Operator_out1543_out1 <= Logical_Operator_out4_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out1544_out1 <= in8 XOR in16;

  Logical_Operator_out1545_out1 <= Logical_Operator_out1033_out1 XOR Logical_Operator_out1037_out1;

  Logical_Operator_out1546_out1 <= Logical_Operator_out1034_out1 XOR Logical_Operator_out1038_out1;

  Logical_Operator_out1547_out1 <= Logical_Operator_out1035_out1 XOR Logical_Operator_out1039_out1;

  Logical_Operator_out1548_out1 <= Logical_Operator_out1036_out1 XOR Logical_Operator_out1040_out1;

  Logical_Operator_out1549_out1 <= Logical_Operator_out523_out1 XOR Logical_Operator_out527_out1;

  Logical_Operator_out1550_out1 <= Logical_Operator_out524_out1 XOR Logical_Operator_out528_out1;

  Logical_Operator_out1551_out1 <= Logical_Operator_out12_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out1552_out1 <= in24 XOR in32;

  Logical_Operator_out1553_out1 <= Logical_Operator_out1041_out1 XOR Logical_Operator_out1045_out1;

  Logical_Operator_out1554_out1 <= Logical_Operator_out1042_out1 XOR Logical_Operator_out1046_out1;

  Logical_Operator_out1555_out1 <= Logical_Operator_out1043_out1 XOR Logical_Operator_out1047_out1;

  Logical_Operator_out1556_out1 <= Logical_Operator_out1044_out1 XOR Logical_Operator_out1048_out1;

  Logical_Operator_out1557_out1 <= Logical_Operator_out531_out1 XOR Logical_Operator_out535_out1;

  Logical_Operator_out1558_out1 <= Logical_Operator_out532_out1 XOR Logical_Operator_out536_out1;

  Logical_Operator_out1559_out1 <= Logical_Operator_out20_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out1560_out1 <= in40 XOR in48;

  Logical_Operator_out1561_out1 <= Logical_Operator_out1049_out1 XOR Logical_Operator_out1053_out1;

  Logical_Operator_out1562_out1 <= Logical_Operator_out1050_out1 XOR Logical_Operator_out1054_out1;

  Logical_Operator_out1563_out1 <= Logical_Operator_out1051_out1 XOR Logical_Operator_out1055_out1;

  Logical_Operator_out1564_out1 <= Logical_Operator_out1052_out1 XOR Logical_Operator_out1056_out1;

  Logical_Operator_out1565_out1 <= Logical_Operator_out539_out1 XOR Logical_Operator_out543_out1;

  Logical_Operator_out1566_out1 <= Logical_Operator_out540_out1 XOR Logical_Operator_out544_out1;

  Logical_Operator_out1567_out1 <= Logical_Operator_out28_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out1568_out1 <= in56 XOR in64;

  Logical_Operator_out1569_out1 <= Logical_Operator_out1057_out1 XOR Logical_Operator_out1061_out1;

  Logical_Operator_out1570_out1 <= Logical_Operator_out1058_out1 XOR Logical_Operator_out1062_out1;

  Logical_Operator_out1571_out1 <= Logical_Operator_out1059_out1 XOR Logical_Operator_out1063_out1;

  Logical_Operator_out1572_out1 <= Logical_Operator_out1060_out1 XOR Logical_Operator_out1064_out1;

  Logical_Operator_out1573_out1 <= Logical_Operator_out547_out1 XOR Logical_Operator_out551_out1;

  Logical_Operator_out1574_out1 <= Logical_Operator_out548_out1 XOR Logical_Operator_out552_out1;

  Logical_Operator_out1575_out1 <= Logical_Operator_out36_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out1576_out1 <= in72 XOR in80;

  Logical_Operator_out1577_out1 <= Logical_Operator_out1065_out1 XOR Logical_Operator_out1069_out1;

  Logical_Operator_out1578_out1 <= Logical_Operator_out1066_out1 XOR Logical_Operator_out1070_out1;

  Logical_Operator_out1579_out1 <= Logical_Operator_out1067_out1 XOR Logical_Operator_out1071_out1;

  Logical_Operator_out1580_out1 <= Logical_Operator_out1068_out1 XOR Logical_Operator_out1072_out1;

  Logical_Operator_out1581_out1 <= Logical_Operator_out555_out1 XOR Logical_Operator_out559_out1;

  Logical_Operator_out1582_out1 <= Logical_Operator_out556_out1 XOR Logical_Operator_out560_out1;

  Logical_Operator_out1583_out1 <= Logical_Operator_out44_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out1584_out1 <= in88 XOR in96;

  Logical_Operator_out1585_out1 <= Logical_Operator_out1073_out1 XOR Logical_Operator_out1077_out1;

  Logical_Operator_out1586_out1 <= Logical_Operator_out1074_out1 XOR Logical_Operator_out1078_out1;

  Logical_Operator_out1587_out1 <= Logical_Operator_out1075_out1 XOR Logical_Operator_out1079_out1;

  Logical_Operator_out1588_out1 <= Logical_Operator_out1076_out1 XOR Logical_Operator_out1080_out1;

  Logical_Operator_out1589_out1 <= Logical_Operator_out563_out1 XOR Logical_Operator_out567_out1;

  Logical_Operator_out1590_out1 <= Logical_Operator_out564_out1 XOR Logical_Operator_out568_out1;

  Logical_Operator_out1591_out1 <= Logical_Operator_out52_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out1592_out1 <= in104 XOR in112;

  Logical_Operator_out1593_out1 <= Logical_Operator_out1081_out1 XOR Logical_Operator_out1085_out1;

  Logical_Operator_out1594_out1 <= Logical_Operator_out1082_out1 XOR Logical_Operator_out1086_out1;

  Logical_Operator_out1595_out1 <= Logical_Operator_out1083_out1 XOR Logical_Operator_out1087_out1;

  Logical_Operator_out1596_out1 <= Logical_Operator_out1084_out1 XOR Logical_Operator_out1088_out1;

  Logical_Operator_out1597_out1 <= Logical_Operator_out571_out1 XOR Logical_Operator_out575_out1;

  Logical_Operator_out1598_out1 <= Logical_Operator_out572_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out1599_out1 <= Logical_Operator_out60_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out1600_out1 <= in120 XOR in128;

  Logical_Operator_out1601_out1 <= Logical_Operator_out1089_out1 XOR Logical_Operator_out1093_out1;

  Logical_Operator_out1602_out1 <= Logical_Operator_out1090_out1 XOR Logical_Operator_out1094_out1;

  Logical_Operator_out1603_out1 <= Logical_Operator_out1091_out1 XOR Logical_Operator_out1095_out1;

  Logical_Operator_out1604_out1 <= Logical_Operator_out1092_out1 XOR Logical_Operator_out1096_out1;

  Logical_Operator_out1605_out1 <= Logical_Operator_out579_out1 XOR Logical_Operator_out583_out1;

  Logical_Operator_out1606_out1 <= Logical_Operator_out580_out1 XOR Logical_Operator_out584_out1;

  Logical_Operator_out1607_out1 <= Logical_Operator_out68_out1 XOR Logical_Operator_out72_out1;

  Logical_Operator_out1608_out1 <= in136 XOR in144;

  Logical_Operator_out1609_out1 <= Logical_Operator_out1097_out1 XOR Logical_Operator_out1101_out1;

  Logical_Operator_out1610_out1 <= Logical_Operator_out1098_out1 XOR Logical_Operator_out1102_out1;

  Logical_Operator_out1611_out1 <= Logical_Operator_out1099_out1 XOR Logical_Operator_out1103_out1;

  Logical_Operator_out1612_out1 <= Logical_Operator_out1100_out1 XOR Logical_Operator_out1104_out1;

  Logical_Operator_out1613_out1 <= Logical_Operator_out587_out1 XOR Logical_Operator_out591_out1;

  Logical_Operator_out1614_out1 <= Logical_Operator_out588_out1 XOR Logical_Operator_out592_out1;

  Logical_Operator_out1615_out1 <= Logical_Operator_out76_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out1616_out1 <= in152 XOR in160;

  Logical_Operator_out1617_out1 <= Logical_Operator_out1105_out1 XOR Logical_Operator_out1109_out1;

  Logical_Operator_out1618_out1 <= Logical_Operator_out1106_out1 XOR Logical_Operator_out1110_out1;

  Logical_Operator_out1619_out1 <= Logical_Operator_out1107_out1 XOR Logical_Operator_out1111_out1;

  Logical_Operator_out1620_out1 <= Logical_Operator_out1108_out1 XOR Logical_Operator_out1112_out1;

  Logical_Operator_out1621_out1 <= Logical_Operator_out595_out1 XOR Logical_Operator_out599_out1;

  Logical_Operator_out1622_out1 <= Logical_Operator_out596_out1 XOR Logical_Operator_out600_out1;

  Logical_Operator_out1623_out1 <= Logical_Operator_out84_out1 XOR Logical_Operator_out88_out1;

  Logical_Operator_out1624_out1 <= in168 XOR in176;

  Logical_Operator_out1625_out1 <= Logical_Operator_out1113_out1 XOR Logical_Operator_out1117_out1;

  Logical_Operator_out1626_out1 <= Logical_Operator_out1114_out1 XOR Logical_Operator_out1118_out1;

  Logical_Operator_out1627_out1 <= Logical_Operator_out1115_out1 XOR Logical_Operator_out1119_out1;

  Logical_Operator_out1628_out1 <= Logical_Operator_out1116_out1 XOR Logical_Operator_out1120_out1;

  Logical_Operator_out1629_out1 <= Logical_Operator_out603_out1 XOR Logical_Operator_out607_out1;

  Logical_Operator_out1630_out1 <= Logical_Operator_out604_out1 XOR Logical_Operator_out608_out1;

  Logical_Operator_out1631_out1 <= Logical_Operator_out92_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out1632_out1 <= in184 XOR in192;

  Logical_Operator_out1633_out1 <= Logical_Operator_out1121_out1 XOR Logical_Operator_out1125_out1;

  Logical_Operator_out1634_out1 <= Logical_Operator_out1122_out1 XOR Logical_Operator_out1126_out1;

  Logical_Operator_out1635_out1 <= Logical_Operator_out1123_out1 XOR Logical_Operator_out1127_out1;

  Logical_Operator_out1636_out1 <= Logical_Operator_out1124_out1 XOR Logical_Operator_out1128_out1;

  Logical_Operator_out1637_out1 <= Logical_Operator_out611_out1 XOR Logical_Operator_out615_out1;

  Logical_Operator_out1638_out1 <= Logical_Operator_out612_out1 XOR Logical_Operator_out616_out1;

  Logical_Operator_out1639_out1 <= Logical_Operator_out100_out1 XOR Logical_Operator_out104_out1;

  Logical_Operator_out1640_out1 <= in200 XOR in208;

  Logical_Operator_out1641_out1 <= Logical_Operator_out1129_out1 XOR Logical_Operator_out1133_out1;

  Logical_Operator_out1642_out1 <= Logical_Operator_out1130_out1 XOR Logical_Operator_out1134_out1;

  Logical_Operator_out1643_out1 <= Logical_Operator_out1131_out1 XOR Logical_Operator_out1135_out1;

  Logical_Operator_out1644_out1 <= Logical_Operator_out1132_out1 XOR Logical_Operator_out1136_out1;

  Logical_Operator_out1645_out1 <= Logical_Operator_out619_out1 XOR Logical_Operator_out623_out1;

  Logical_Operator_out1646_out1 <= Logical_Operator_out620_out1 XOR Logical_Operator_out624_out1;

  Logical_Operator_out1647_out1 <= Logical_Operator_out108_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out1648_out1 <= in216 XOR in224;

  Logical_Operator_out1649_out1 <= Logical_Operator_out1137_out1 XOR Logical_Operator_out1141_out1;

  Logical_Operator_out1650_out1 <= Logical_Operator_out1138_out1 XOR Logical_Operator_out1142_out1;

  Logical_Operator_out1651_out1 <= Logical_Operator_out1139_out1 XOR Logical_Operator_out1143_out1;

  Logical_Operator_out1652_out1 <= Logical_Operator_out1140_out1 XOR Logical_Operator_out1144_out1;

  Logical_Operator_out1653_out1 <= Logical_Operator_out627_out1 XOR Logical_Operator_out631_out1;

  Logical_Operator_out1654_out1 <= Logical_Operator_out628_out1 XOR Logical_Operator_out632_out1;

  Logical_Operator_out1655_out1 <= Logical_Operator_out116_out1 XOR Logical_Operator_out120_out1;

  Logical_Operator_out1656_out1 <= in232 XOR in240;

  Logical_Operator_out1657_out1 <= Logical_Operator_out1145_out1 XOR Logical_Operator_out1149_out1;

  Logical_Operator_out1658_out1 <= Logical_Operator_out1146_out1 XOR Logical_Operator_out1150_out1;

  Logical_Operator_out1659_out1 <= Logical_Operator_out1147_out1 XOR Logical_Operator_out1151_out1;

  Logical_Operator_out1660_out1 <= Logical_Operator_out1148_out1 XOR Logical_Operator_out1152_out1;

  Logical_Operator_out1661_out1 <= Logical_Operator_out635_out1 XOR Logical_Operator_out639_out1;

  Logical_Operator_out1662_out1 <= Logical_Operator_out636_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out1663_out1 <= Logical_Operator_out124_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out1664_out1 <= in248 XOR in256;

  Logical_Operator_out1665_out1 <= Logical_Operator_out1153_out1 XOR Logical_Operator_out1157_out1;

  Logical_Operator_out1666_out1 <= Logical_Operator_out1154_out1 XOR Logical_Operator_out1158_out1;

  Logical_Operator_out1667_out1 <= Logical_Operator_out1155_out1 XOR Logical_Operator_out1159_out1;

  Logical_Operator_out1668_out1 <= Logical_Operator_out1156_out1 XOR Logical_Operator_out1160_out1;

  Logical_Operator_out1669_out1 <= Logical_Operator_out643_out1 XOR Logical_Operator_out647_out1;

  Logical_Operator_out1670_out1 <= Logical_Operator_out644_out1 XOR Logical_Operator_out648_out1;

  Logical_Operator_out1671_out1 <= Logical_Operator_out132_out1 XOR Logical_Operator_out136_out1;

  Logical_Operator_out1672_out1 <= in264 XOR in272;

  Logical_Operator_out1673_out1 <= Logical_Operator_out1161_out1 XOR Logical_Operator_out1165_out1;

  Logical_Operator_out1674_out1 <= Logical_Operator_out1162_out1 XOR Logical_Operator_out1166_out1;

  Logical_Operator_out1675_out1 <= Logical_Operator_out1163_out1 XOR Logical_Operator_out1167_out1;

  Logical_Operator_out1676_out1 <= Logical_Operator_out1164_out1 XOR Logical_Operator_out1168_out1;

  Logical_Operator_out1677_out1 <= Logical_Operator_out651_out1 XOR Logical_Operator_out655_out1;

  Logical_Operator_out1678_out1 <= Logical_Operator_out652_out1 XOR Logical_Operator_out656_out1;

  Logical_Operator_out1679_out1 <= Logical_Operator_out140_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out1680_out1 <= in280 XOR in288;

  Logical_Operator_out1681_out1 <= Logical_Operator_out1169_out1 XOR Logical_Operator_out1173_out1;

  Logical_Operator_out1682_out1 <= Logical_Operator_out1170_out1 XOR Logical_Operator_out1174_out1;

  Logical_Operator_out1683_out1 <= Logical_Operator_out1171_out1 XOR Logical_Operator_out1175_out1;

  Logical_Operator_out1684_out1 <= Logical_Operator_out1172_out1 XOR Logical_Operator_out1176_out1;

  Logical_Operator_out1685_out1 <= Logical_Operator_out659_out1 XOR Logical_Operator_out663_out1;

  Logical_Operator_out1686_out1 <= Logical_Operator_out660_out1 XOR Logical_Operator_out664_out1;

  Logical_Operator_out1687_out1 <= Logical_Operator_out148_out1 XOR Logical_Operator_out152_out1;

  Logical_Operator_out1688_out1 <= in296 XOR in304;

  Logical_Operator_out1689_out1 <= Logical_Operator_out1177_out1 XOR Logical_Operator_out1181_out1;

  Logical_Operator_out1690_out1 <= Logical_Operator_out1178_out1 XOR Logical_Operator_out1182_out1;

  Logical_Operator_out1691_out1 <= Logical_Operator_out1179_out1 XOR Logical_Operator_out1183_out1;

  Logical_Operator_out1692_out1 <= Logical_Operator_out1180_out1 XOR Logical_Operator_out1184_out1;

  Logical_Operator_out1693_out1 <= Logical_Operator_out667_out1 XOR Logical_Operator_out671_out1;

  Logical_Operator_out1694_out1 <= Logical_Operator_out668_out1 XOR Logical_Operator_out672_out1;

  Logical_Operator_out1695_out1 <= Logical_Operator_out156_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out1696_out1 <= in312 XOR in320;

  Logical_Operator_out1697_out1 <= Logical_Operator_out1185_out1 XOR Logical_Operator_out1189_out1;

  Logical_Operator_out1698_out1 <= Logical_Operator_out1186_out1 XOR Logical_Operator_out1190_out1;

  Logical_Operator_out1699_out1 <= Logical_Operator_out1187_out1 XOR Logical_Operator_out1191_out1;

  Logical_Operator_out1700_out1 <= Logical_Operator_out1188_out1 XOR Logical_Operator_out1192_out1;

  Logical_Operator_out1701_out1 <= Logical_Operator_out675_out1 XOR Logical_Operator_out679_out1;

  Logical_Operator_out1702_out1 <= Logical_Operator_out676_out1 XOR Logical_Operator_out680_out1;

  Logical_Operator_out1703_out1 <= Logical_Operator_out164_out1 XOR Logical_Operator_out168_out1;

  Logical_Operator_out1704_out1 <= in328 XOR in336;

  Logical_Operator_out1705_out1 <= Logical_Operator_out1193_out1 XOR Logical_Operator_out1197_out1;

  Logical_Operator_out1706_out1 <= Logical_Operator_out1194_out1 XOR Logical_Operator_out1198_out1;

  Logical_Operator_out1707_out1 <= Logical_Operator_out1195_out1 XOR Logical_Operator_out1199_out1;

  Logical_Operator_out1708_out1 <= Logical_Operator_out1196_out1 XOR Logical_Operator_out1200_out1;

  Logical_Operator_out1709_out1 <= Logical_Operator_out683_out1 XOR Logical_Operator_out687_out1;

  Logical_Operator_out1710_out1 <= Logical_Operator_out684_out1 XOR Logical_Operator_out688_out1;

  Logical_Operator_out1711_out1 <= Logical_Operator_out172_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out1712_out1 <= in344 XOR in352;

  Logical_Operator_out1713_out1 <= Logical_Operator_out1201_out1 XOR Logical_Operator_out1205_out1;

  Logical_Operator_out1714_out1 <= Logical_Operator_out1202_out1 XOR Logical_Operator_out1206_out1;

  Logical_Operator_out1715_out1 <= Logical_Operator_out1203_out1 XOR Logical_Operator_out1207_out1;

  Logical_Operator_out1716_out1 <= Logical_Operator_out1204_out1 XOR Logical_Operator_out1208_out1;

  Logical_Operator_out1717_out1 <= Logical_Operator_out691_out1 XOR Logical_Operator_out695_out1;

  Logical_Operator_out1718_out1 <= Logical_Operator_out692_out1 XOR Logical_Operator_out696_out1;

  Logical_Operator_out1719_out1 <= Logical_Operator_out180_out1 XOR Logical_Operator_out184_out1;

  Logical_Operator_out1720_out1 <= in360 XOR in368;

  Logical_Operator_out1721_out1 <= Logical_Operator_out1209_out1 XOR Logical_Operator_out1213_out1;

  Logical_Operator_out1722_out1 <= Logical_Operator_out1210_out1 XOR Logical_Operator_out1214_out1;

  Logical_Operator_out1723_out1 <= Logical_Operator_out1211_out1 XOR Logical_Operator_out1215_out1;

  Logical_Operator_out1724_out1 <= Logical_Operator_out1212_out1 XOR Logical_Operator_out1216_out1;

  Logical_Operator_out1725_out1 <= Logical_Operator_out699_out1 XOR Logical_Operator_out703_out1;

  Logical_Operator_out1726_out1 <= Logical_Operator_out700_out1 XOR Logical_Operator_out704_out1;

  Logical_Operator_out1727_out1 <= Logical_Operator_out188_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out1728_out1 <= in376 XOR in384;

  Logical_Operator_out1729_out1 <= Logical_Operator_out1217_out1 XOR Logical_Operator_out1221_out1;

  Logical_Operator_out1730_out1 <= Logical_Operator_out1218_out1 XOR Logical_Operator_out1222_out1;

  Logical_Operator_out1731_out1 <= Logical_Operator_out1219_out1 XOR Logical_Operator_out1223_out1;

  Logical_Operator_out1732_out1 <= Logical_Operator_out1220_out1 XOR Logical_Operator_out1224_out1;

  Logical_Operator_out1733_out1 <= Logical_Operator_out707_out1 XOR Logical_Operator_out711_out1;

  Logical_Operator_out1734_out1 <= Logical_Operator_out708_out1 XOR Logical_Operator_out712_out1;

  Logical_Operator_out1735_out1 <= Logical_Operator_out196_out1 XOR Logical_Operator_out200_out1;

  Logical_Operator_out1736_out1 <= in392 XOR in400;

  Logical_Operator_out1737_out1 <= Logical_Operator_out1225_out1 XOR Logical_Operator_out1229_out1;

  Logical_Operator_out1738_out1 <= Logical_Operator_out1226_out1 XOR Logical_Operator_out1230_out1;

  Logical_Operator_out1739_out1 <= Logical_Operator_out1227_out1 XOR Logical_Operator_out1231_out1;

  Logical_Operator_out1740_out1 <= Logical_Operator_out1228_out1 XOR Logical_Operator_out1232_out1;

  Logical_Operator_out1741_out1 <= Logical_Operator_out715_out1 XOR Logical_Operator_out719_out1;

  Logical_Operator_out1742_out1 <= Logical_Operator_out716_out1 XOR Logical_Operator_out720_out1;

  Logical_Operator_out1743_out1 <= Logical_Operator_out204_out1 XOR Logical_Operator_out208_out1;

  Logical_Operator_out1744_out1 <= in408 XOR in416;

  Logical_Operator_out1745_out1 <= Logical_Operator_out1233_out1 XOR Logical_Operator_out1237_out1;

  Logical_Operator_out1746_out1 <= Logical_Operator_out1234_out1 XOR Logical_Operator_out1238_out1;

  Logical_Operator_out1747_out1 <= Logical_Operator_out1235_out1 XOR Logical_Operator_out1239_out1;

  Logical_Operator_out1748_out1 <= Logical_Operator_out1236_out1 XOR Logical_Operator_out1240_out1;

  Logical_Operator_out1749_out1 <= Logical_Operator_out723_out1 XOR Logical_Operator_out727_out1;

  Logical_Operator_out1750_out1 <= Logical_Operator_out724_out1 XOR Logical_Operator_out728_out1;

  Logical_Operator_out1751_out1 <= Logical_Operator_out212_out1 XOR Logical_Operator_out216_out1;

  Logical_Operator_out1752_out1 <= in424 XOR in432;

  Logical_Operator_out1753_out1 <= Logical_Operator_out1241_out1 XOR Logical_Operator_out1245_out1;

  Logical_Operator_out1754_out1 <= Logical_Operator_out1242_out1 XOR Logical_Operator_out1246_out1;

  Logical_Operator_out1755_out1 <= Logical_Operator_out1243_out1 XOR Logical_Operator_out1247_out1;

  Logical_Operator_out1756_out1 <= Logical_Operator_out1244_out1 XOR Logical_Operator_out1248_out1;

  Logical_Operator_out1757_out1 <= Logical_Operator_out731_out1 XOR Logical_Operator_out735_out1;

  Logical_Operator_out1758_out1 <= Logical_Operator_out732_out1 XOR Logical_Operator_out736_out1;

  Logical_Operator_out1759_out1 <= Logical_Operator_out220_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out1760_out1 <= in440 XOR in448;

  Logical_Operator_out1761_out1 <= Logical_Operator_out1249_out1 XOR Logical_Operator_out1253_out1;

  Logical_Operator_out1762_out1 <= Logical_Operator_out1250_out1 XOR Logical_Operator_out1254_out1;

  Logical_Operator_out1763_out1 <= Logical_Operator_out1251_out1 XOR Logical_Operator_out1255_out1;

  Logical_Operator_out1764_out1 <= Logical_Operator_out1252_out1 XOR Logical_Operator_out1256_out1;

  Logical_Operator_out1765_out1 <= Logical_Operator_out739_out1 XOR Logical_Operator_out743_out1;

  Logical_Operator_out1766_out1 <= Logical_Operator_out740_out1 XOR Logical_Operator_out744_out1;

  Logical_Operator_out1767_out1 <= Logical_Operator_out228_out1 XOR Logical_Operator_out232_out1;

  Logical_Operator_out1768_out1 <= in456 XOR in464;

  Logical_Operator_out1769_out1 <= Logical_Operator_out1257_out1 XOR Logical_Operator_out1261_out1;

  Logical_Operator_out1770_out1 <= Logical_Operator_out1258_out1 XOR Logical_Operator_out1262_out1;

  Logical_Operator_out1771_out1 <= Logical_Operator_out1259_out1 XOR Logical_Operator_out1263_out1;

  Logical_Operator_out1772_out1 <= Logical_Operator_out1260_out1 XOR Logical_Operator_out1264_out1;

  Logical_Operator_out1773_out1 <= Logical_Operator_out747_out1 XOR Logical_Operator_out751_out1;

  Logical_Operator_out1774_out1 <= Logical_Operator_out748_out1 XOR Logical_Operator_out752_out1;

  Logical_Operator_out1775_out1 <= Logical_Operator_out236_out1 XOR Logical_Operator_out240_out1;

  Logical_Operator_out1776_out1 <= in472 XOR in480;

  Logical_Operator_out1777_out1 <= Logical_Operator_out1265_out1 XOR Logical_Operator_out1269_out1;

  Logical_Operator_out1778_out1 <= Logical_Operator_out1266_out1 XOR Logical_Operator_out1270_out1;

  Logical_Operator_out1779_out1 <= Logical_Operator_out1267_out1 XOR Logical_Operator_out1271_out1;

  Logical_Operator_out1780_out1 <= Logical_Operator_out1268_out1 XOR Logical_Operator_out1272_out1;

  Logical_Operator_out1781_out1 <= Logical_Operator_out755_out1 XOR Logical_Operator_out759_out1;

  Logical_Operator_out1782_out1 <= Logical_Operator_out756_out1 XOR Logical_Operator_out760_out1;

  Logical_Operator_out1783_out1 <= Logical_Operator_out244_out1 XOR Logical_Operator_out248_out1;

  Logical_Operator_out1784_out1 <= in488 XOR in496;

  Logical_Operator_out1785_out1 <= Logical_Operator_out1273_out1 XOR Logical_Operator_out1277_out1;

  Logical_Operator_out1786_out1 <= Logical_Operator_out1274_out1 XOR Logical_Operator_out1278_out1;

  Logical_Operator_out1787_out1 <= Logical_Operator_out1275_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out1788_out1 <= Logical_Operator_out1276_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out1789_out1 <= Logical_Operator_out763_out1 XOR Logical_Operator_out767_out1;

  Logical_Operator_out1790_out1 <= Logical_Operator_out764_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out1791_out1 <= Logical_Operator_out252_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out1792_out1 <= in504 XOR in512;

  Logical_Operator_out1793_out1 <= Logical_Operator_out1281_out1 XOR Logical_Operator_out1285_out1;

  Logical_Operator_out1794_out1 <= Logical_Operator_out1282_out1 XOR Logical_Operator_out1286_out1;

  Logical_Operator_out1795_out1 <= Logical_Operator_out1283_out1 XOR Logical_Operator_out1287_out1;

  Logical_Operator_out1796_out1 <= Logical_Operator_out1284_out1 XOR Logical_Operator_out1288_out1;

  Logical_Operator_out1797_out1 <= Logical_Operator_out771_out1 XOR Logical_Operator_out775_out1;

  Logical_Operator_out1798_out1 <= Logical_Operator_out772_out1 XOR Logical_Operator_out776_out1;

  Logical_Operator_out1799_out1 <= Logical_Operator_out260_out1 XOR Logical_Operator_out264_out1;

  Logical_Operator_out1800_out1 <= in520 XOR in528;

  Logical_Operator_out1801_out1 <= Logical_Operator_out1289_out1 XOR Logical_Operator_out1293_out1;

  Logical_Operator_out1802_out1 <= Logical_Operator_out1290_out1 XOR Logical_Operator_out1294_out1;

  Logical_Operator_out1803_out1 <= Logical_Operator_out1291_out1 XOR Logical_Operator_out1295_out1;

  Logical_Operator_out1804_out1 <= Logical_Operator_out1292_out1 XOR Logical_Operator_out1296_out1;

  Logical_Operator_out1805_out1 <= Logical_Operator_out779_out1 XOR Logical_Operator_out783_out1;

  Logical_Operator_out1806_out1 <= Logical_Operator_out780_out1 XOR Logical_Operator_out784_out1;

  Logical_Operator_out1807_out1 <= Logical_Operator_out268_out1 XOR Logical_Operator_out272_out1;

  Logical_Operator_out1808_out1 <= in536 XOR in544;

  Logical_Operator_out1809_out1 <= Logical_Operator_out1297_out1 XOR Logical_Operator_out1301_out1;

  Logical_Operator_out1810_out1 <= Logical_Operator_out1298_out1 XOR Logical_Operator_out1302_out1;

  Logical_Operator_out1811_out1 <= Logical_Operator_out1299_out1 XOR Logical_Operator_out1303_out1;

  Logical_Operator_out1812_out1 <= Logical_Operator_out1300_out1 XOR Logical_Operator_out1304_out1;

  Logical_Operator_out1813_out1 <= Logical_Operator_out787_out1 XOR Logical_Operator_out791_out1;

  Logical_Operator_out1814_out1 <= Logical_Operator_out788_out1 XOR Logical_Operator_out792_out1;

  Logical_Operator_out1815_out1 <= Logical_Operator_out276_out1 XOR Logical_Operator_out280_out1;

  Logical_Operator_out1816_out1 <= in552 XOR in560;

  Logical_Operator_out1817_out1 <= Logical_Operator_out1305_out1 XOR Logical_Operator_out1309_out1;

  Logical_Operator_out1818_out1 <= Logical_Operator_out1306_out1 XOR Logical_Operator_out1310_out1;

  Logical_Operator_out1819_out1 <= Logical_Operator_out1307_out1 XOR Logical_Operator_out1311_out1;

  Logical_Operator_out1820_out1 <= Logical_Operator_out1308_out1 XOR Logical_Operator_out1312_out1;

  Logical_Operator_out1821_out1 <= Logical_Operator_out795_out1 XOR Logical_Operator_out799_out1;

  Logical_Operator_out1822_out1 <= Logical_Operator_out796_out1 XOR Logical_Operator_out800_out1;

  Logical_Operator_out1823_out1 <= Logical_Operator_out284_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out1824_out1 <= in568 XOR in576;

  Logical_Operator_out1825_out1 <= Logical_Operator_out1313_out1 XOR Logical_Operator_out1317_out1;

  Logical_Operator_out1826_out1 <= Logical_Operator_out1314_out1 XOR Logical_Operator_out1318_out1;

  Logical_Operator_out1827_out1 <= Logical_Operator_out1315_out1 XOR Logical_Operator_out1319_out1;

  Logical_Operator_out1828_out1 <= Logical_Operator_out1316_out1 XOR Logical_Operator_out1320_out1;

  Logical_Operator_out1829_out1 <= Logical_Operator_out803_out1 XOR Logical_Operator_out807_out1;

  Logical_Operator_out1830_out1 <= Logical_Operator_out804_out1 XOR Logical_Operator_out808_out1;

  Logical_Operator_out1831_out1 <= Logical_Operator_out292_out1 XOR Logical_Operator_out296_out1;

  Logical_Operator_out1832_out1 <= in584 XOR in592;

  Logical_Operator_out1833_out1 <= Logical_Operator_out1321_out1 XOR Logical_Operator_out1325_out1;

  Logical_Operator_out1834_out1 <= Logical_Operator_out1322_out1 XOR Logical_Operator_out1326_out1;

  Logical_Operator_out1835_out1 <= Logical_Operator_out1323_out1 XOR Logical_Operator_out1327_out1;

  Logical_Operator_out1836_out1 <= Logical_Operator_out1324_out1 XOR Logical_Operator_out1328_out1;

  Logical_Operator_out1837_out1 <= Logical_Operator_out811_out1 XOR Logical_Operator_out815_out1;

  Logical_Operator_out1838_out1 <= Logical_Operator_out812_out1 XOR Logical_Operator_out816_out1;

  Logical_Operator_out1839_out1 <= Logical_Operator_out300_out1 XOR Logical_Operator_out304_out1;

  Logical_Operator_out1840_out1 <= in600 XOR in608;

  Logical_Operator_out1841_out1 <= Logical_Operator_out1329_out1 XOR Logical_Operator_out1333_out1;

  Logical_Operator_out1842_out1 <= Logical_Operator_out1330_out1 XOR Logical_Operator_out1334_out1;

  Logical_Operator_out1843_out1 <= Logical_Operator_out1331_out1 XOR Logical_Operator_out1335_out1;

  Logical_Operator_out1844_out1 <= Logical_Operator_out1332_out1 XOR Logical_Operator_out1336_out1;

  Logical_Operator_out1845_out1 <= Logical_Operator_out819_out1 XOR Logical_Operator_out823_out1;

  Logical_Operator_out1846_out1 <= Logical_Operator_out820_out1 XOR Logical_Operator_out824_out1;

  Logical_Operator_out1847_out1 <= Logical_Operator_out308_out1 XOR Logical_Operator_out312_out1;

  Logical_Operator_out1848_out1 <= in616 XOR in624;

  Logical_Operator_out1849_out1 <= Logical_Operator_out1337_out1 XOR Logical_Operator_out1341_out1;

  Logical_Operator_out1850_out1 <= Logical_Operator_out1338_out1 XOR Logical_Operator_out1342_out1;

  Logical_Operator_out1851_out1 <= Logical_Operator_out1339_out1 XOR Logical_Operator_out1343_out1;

  Logical_Operator_out1852_out1 <= Logical_Operator_out1340_out1 XOR Logical_Operator_out1344_out1;

  Logical_Operator_out1853_out1 <= Logical_Operator_out827_out1 XOR Logical_Operator_out831_out1;

  Logical_Operator_out1854_out1 <= Logical_Operator_out828_out1 XOR Logical_Operator_out832_out1;

  Logical_Operator_out1855_out1 <= Logical_Operator_out316_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out1856_out1 <= in632 XOR in640;

  Logical_Operator_out1857_out1 <= Logical_Operator_out1345_out1 XOR Logical_Operator_out1349_out1;

  Logical_Operator_out1858_out1 <= Logical_Operator_out1346_out1 XOR Logical_Operator_out1350_out1;

  Logical_Operator_out1859_out1 <= Logical_Operator_out1347_out1 XOR Logical_Operator_out1351_out1;

  Logical_Operator_out1860_out1 <= Logical_Operator_out1348_out1 XOR Logical_Operator_out1352_out1;

  Logical_Operator_out1861_out1 <= Logical_Operator_out835_out1 XOR Logical_Operator_out839_out1;

  Logical_Operator_out1862_out1 <= Logical_Operator_out836_out1 XOR Logical_Operator_out840_out1;

  Logical_Operator_out1863_out1 <= Logical_Operator_out324_out1 XOR Logical_Operator_out328_out1;

  Logical_Operator_out1864_out1 <= in648 XOR in656;

  Logical_Operator_out1865_out1 <= Logical_Operator_out1353_out1 XOR Logical_Operator_out1357_out1;

  Logical_Operator_out1866_out1 <= Logical_Operator_out1354_out1 XOR Logical_Operator_out1358_out1;

  Logical_Operator_out1867_out1 <= Logical_Operator_out1355_out1 XOR Logical_Operator_out1359_out1;

  Logical_Operator_out1868_out1 <= Logical_Operator_out1356_out1 XOR Logical_Operator_out1360_out1;

  Logical_Operator_out1869_out1 <= Logical_Operator_out843_out1 XOR Logical_Operator_out847_out1;

  Logical_Operator_out1870_out1 <= Logical_Operator_out844_out1 XOR Logical_Operator_out848_out1;

  Logical_Operator_out1871_out1 <= Logical_Operator_out332_out1 XOR Logical_Operator_out336_out1;

  Logical_Operator_out1872_out1 <= in664 XOR in672;

  Logical_Operator_out1873_out1 <= Logical_Operator_out1361_out1 XOR Logical_Operator_out1365_out1;

  Logical_Operator_out1874_out1 <= Logical_Operator_out1362_out1 XOR Logical_Operator_out1366_out1;

  Logical_Operator_out1875_out1 <= Logical_Operator_out1363_out1 XOR Logical_Operator_out1367_out1;

  Logical_Operator_out1876_out1 <= Logical_Operator_out1364_out1 XOR Logical_Operator_out1368_out1;

  Logical_Operator_out1877_out1 <= Logical_Operator_out851_out1 XOR Logical_Operator_out855_out1;

  Logical_Operator_out1878_out1 <= Logical_Operator_out852_out1 XOR Logical_Operator_out856_out1;

  Logical_Operator_out1879_out1 <= Logical_Operator_out340_out1 XOR Logical_Operator_out344_out1;

  Logical_Operator_out1880_out1 <= in680 XOR in688;

  Logical_Operator_out1881_out1 <= Logical_Operator_out1369_out1 XOR Logical_Operator_out1373_out1;

  Logical_Operator_out1882_out1 <= Logical_Operator_out1370_out1 XOR Logical_Operator_out1374_out1;

  Logical_Operator_out1883_out1 <= Logical_Operator_out1371_out1 XOR Logical_Operator_out1375_out1;

  Logical_Operator_out1884_out1 <= Logical_Operator_out1372_out1 XOR Logical_Operator_out1376_out1;

  Logical_Operator_out1885_out1 <= Logical_Operator_out859_out1 XOR Logical_Operator_out863_out1;

  Logical_Operator_out1886_out1 <= Logical_Operator_out860_out1 XOR Logical_Operator_out864_out1;

  Logical_Operator_out1887_out1 <= Logical_Operator_out348_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out1888_out1 <= in696 XOR in704;

  Logical_Operator_out1889_out1 <= Logical_Operator_out1377_out1 XOR Logical_Operator_out1381_out1;

  Logical_Operator_out1890_out1 <= Logical_Operator_out1378_out1 XOR Logical_Operator_out1382_out1;

  Logical_Operator_out1891_out1 <= Logical_Operator_out1379_out1 XOR Logical_Operator_out1383_out1;

  Logical_Operator_out1892_out1 <= Logical_Operator_out1380_out1 XOR Logical_Operator_out1384_out1;

  Logical_Operator_out1893_out1 <= Logical_Operator_out867_out1 XOR Logical_Operator_out871_out1;

  Logical_Operator_out1894_out1 <= Logical_Operator_out868_out1 XOR Logical_Operator_out872_out1;

  Logical_Operator_out1895_out1 <= Logical_Operator_out356_out1 XOR Logical_Operator_out360_out1;

  Logical_Operator_out1896_out1 <= in712 XOR in720;

  Logical_Operator_out1897_out1 <= Logical_Operator_out1385_out1 XOR Logical_Operator_out1389_out1;

  Logical_Operator_out1898_out1 <= Logical_Operator_out1386_out1 XOR Logical_Operator_out1390_out1;

  Logical_Operator_out1899_out1 <= Logical_Operator_out1387_out1 XOR Logical_Operator_out1391_out1;

  Logical_Operator_out1900_out1 <= Logical_Operator_out1388_out1 XOR Logical_Operator_out1392_out1;

  Logical_Operator_out1901_out1 <= Logical_Operator_out875_out1 XOR Logical_Operator_out879_out1;

  Logical_Operator_out1902_out1 <= Logical_Operator_out876_out1 XOR Logical_Operator_out880_out1;

  Logical_Operator_out1903_out1 <= Logical_Operator_out364_out1 XOR Logical_Operator_out368_out1;

  Logical_Operator_out1904_out1 <= in728 XOR in736;

  Logical_Operator_out1905_out1 <= Logical_Operator_out1393_out1 XOR Logical_Operator_out1397_out1;

  Logical_Operator_out1906_out1 <= Logical_Operator_out1394_out1 XOR Logical_Operator_out1398_out1;

  Logical_Operator_out1907_out1 <= Logical_Operator_out1395_out1 XOR Logical_Operator_out1399_out1;

  Logical_Operator_out1908_out1 <= Logical_Operator_out1396_out1 XOR Logical_Operator_out1400_out1;

  Logical_Operator_out1909_out1 <= Logical_Operator_out883_out1 XOR Logical_Operator_out887_out1;

  Logical_Operator_out1910_out1 <= Logical_Operator_out884_out1 XOR Logical_Operator_out888_out1;

  Logical_Operator_out1911_out1 <= Logical_Operator_out372_out1 XOR Logical_Operator_out376_out1;

  Logical_Operator_out1912_out1 <= in744 XOR in752;

  Logical_Operator_out1913_out1 <= Logical_Operator_out1401_out1 XOR Logical_Operator_out1405_out1;

  Logical_Operator_out1914_out1 <= Logical_Operator_out1402_out1 XOR Logical_Operator_out1406_out1;

  Logical_Operator_out1915_out1 <= Logical_Operator_out1403_out1 XOR Logical_Operator_out1407_out1;

  Logical_Operator_out1916_out1 <= Logical_Operator_out1404_out1 XOR Logical_Operator_out1408_out1;

  Logical_Operator_out1917_out1 <= Logical_Operator_out891_out1 XOR Logical_Operator_out895_out1;

  Logical_Operator_out1918_out1 <= Logical_Operator_out892_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out1919_out1 <= Logical_Operator_out380_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out1920_out1 <= in760 XOR in768;

  Logical_Operator_out1921_out1 <= Logical_Operator_out1409_out1 XOR Logical_Operator_out1413_out1;

  Logical_Operator_out1922_out1 <= Logical_Operator_out1410_out1 XOR Logical_Operator_out1414_out1;

  Logical_Operator_out1923_out1 <= Logical_Operator_out1411_out1 XOR Logical_Operator_out1415_out1;

  Logical_Operator_out1924_out1 <= Logical_Operator_out1412_out1 XOR Logical_Operator_out1416_out1;

  Logical_Operator_out1925_out1 <= Logical_Operator_out899_out1 XOR Logical_Operator_out903_out1;

  Logical_Operator_out1926_out1 <= Logical_Operator_out900_out1 XOR Logical_Operator_out904_out1;

  Logical_Operator_out1927_out1 <= Logical_Operator_out388_out1 XOR Logical_Operator_out392_out1;

  Logical_Operator_out1928_out1 <= in776 XOR in784;

  Logical_Operator_out1929_out1 <= Logical_Operator_out1417_out1 XOR Logical_Operator_out1421_out1;

  Logical_Operator_out1930_out1 <= Logical_Operator_out1418_out1 XOR Logical_Operator_out1422_out1;

  Logical_Operator_out1931_out1 <= Logical_Operator_out1419_out1 XOR Logical_Operator_out1423_out1;

  Logical_Operator_out1932_out1 <= Logical_Operator_out1420_out1 XOR Logical_Operator_out1424_out1;

  Logical_Operator_out1933_out1 <= Logical_Operator_out907_out1 XOR Logical_Operator_out911_out1;

  Logical_Operator_out1934_out1 <= Logical_Operator_out908_out1 XOR Logical_Operator_out912_out1;

  Logical_Operator_out1935_out1 <= Logical_Operator_out396_out1 XOR Logical_Operator_out400_out1;

  Logical_Operator_out1936_out1 <= in792 XOR in800;

  Logical_Operator_out1937_out1 <= Logical_Operator_out1425_out1 XOR Logical_Operator_out1429_out1;

  Logical_Operator_out1938_out1 <= Logical_Operator_out1426_out1 XOR Logical_Operator_out1430_out1;

  Logical_Operator_out1939_out1 <= Logical_Operator_out1427_out1 XOR Logical_Operator_out1431_out1;

  Logical_Operator_out1940_out1 <= Logical_Operator_out1428_out1 XOR Logical_Operator_out1432_out1;

  Logical_Operator_out1941_out1 <= Logical_Operator_out915_out1 XOR Logical_Operator_out919_out1;

  Logical_Operator_out1942_out1 <= Logical_Operator_out916_out1 XOR Logical_Operator_out920_out1;

  Logical_Operator_out1943_out1 <= Logical_Operator_out404_out1 XOR Logical_Operator_out408_out1;

  Logical_Operator_out1944_out1 <= in808 XOR in816;

  Logical_Operator_out1945_out1 <= Logical_Operator_out1433_out1 XOR Logical_Operator_out1437_out1;

  Logical_Operator_out1946_out1 <= Logical_Operator_out1434_out1 XOR Logical_Operator_out1438_out1;

  Logical_Operator_out1947_out1 <= Logical_Operator_out1435_out1 XOR Logical_Operator_out1439_out1;

  Logical_Operator_out1948_out1 <= Logical_Operator_out1436_out1 XOR Logical_Operator_out1440_out1;

  Logical_Operator_out1949_out1 <= Logical_Operator_out923_out1 XOR Logical_Operator_out927_out1;

  Logical_Operator_out1950_out1 <= Logical_Operator_out924_out1 XOR Logical_Operator_out928_out1;

  Logical_Operator_out1951_out1 <= Logical_Operator_out412_out1 XOR Logical_Operator_out416_out1;

  Logical_Operator_out1952_out1 <= in824 XOR in832;

  Logical_Operator_out1953_out1 <= Logical_Operator_out1441_out1 XOR Logical_Operator_out1445_out1;

  Logical_Operator_out1954_out1 <= Logical_Operator_out1442_out1 XOR Logical_Operator_out1446_out1;

  Logical_Operator_out1955_out1 <= Logical_Operator_out1443_out1 XOR Logical_Operator_out1447_out1;

  Logical_Operator_out1956_out1 <= Logical_Operator_out1444_out1 XOR Logical_Operator_out1448_out1;

  Logical_Operator_out1957_out1 <= Logical_Operator_out931_out1 XOR Logical_Operator_out935_out1;

  Logical_Operator_out1958_out1 <= Logical_Operator_out932_out1 XOR Logical_Operator_out936_out1;

  Logical_Operator_out1959_out1 <= Logical_Operator_out420_out1 XOR Logical_Operator_out424_out1;

  Logical_Operator_out1960_out1 <= in840 XOR in848;

  Logical_Operator_out1961_out1 <= Logical_Operator_out1449_out1 XOR Logical_Operator_out1453_out1;

  Logical_Operator_out1962_out1 <= Logical_Operator_out1450_out1 XOR Logical_Operator_out1454_out1;

  Logical_Operator_out1963_out1 <= Logical_Operator_out1451_out1 XOR Logical_Operator_out1455_out1;

  Logical_Operator_out1964_out1 <= Logical_Operator_out1452_out1 XOR Logical_Operator_out1456_out1;

  Logical_Operator_out1965_out1 <= Logical_Operator_out939_out1 XOR Logical_Operator_out943_out1;

  Logical_Operator_out1966_out1 <= Logical_Operator_out940_out1 XOR Logical_Operator_out944_out1;

  Logical_Operator_out1967_out1 <= Logical_Operator_out428_out1 XOR Logical_Operator_out432_out1;

  Logical_Operator_out1968_out1 <= in856 XOR in864;

  Logical_Operator_out1969_out1 <= Logical_Operator_out1457_out1 XOR Logical_Operator_out1461_out1;

  Logical_Operator_out1970_out1 <= Logical_Operator_out1458_out1 XOR Logical_Operator_out1462_out1;

  Logical_Operator_out1971_out1 <= Logical_Operator_out1459_out1 XOR Logical_Operator_out1463_out1;

  Logical_Operator_out1972_out1 <= Logical_Operator_out1460_out1 XOR Logical_Operator_out1464_out1;

  Logical_Operator_out1973_out1 <= Logical_Operator_out947_out1 XOR Logical_Operator_out951_out1;

  Logical_Operator_out1974_out1 <= Logical_Operator_out948_out1 XOR Logical_Operator_out952_out1;

  Logical_Operator_out1975_out1 <= Logical_Operator_out436_out1 XOR Logical_Operator_out440_out1;

  Logical_Operator_out1976_out1 <= in872 XOR in880;

  Logical_Operator_out1977_out1 <= Logical_Operator_out1465_out1 XOR Logical_Operator_out1469_out1;

  Logical_Operator_out1978_out1 <= Logical_Operator_out1466_out1 XOR Logical_Operator_out1470_out1;

  Logical_Operator_out1979_out1 <= Logical_Operator_out1467_out1 XOR Logical_Operator_out1471_out1;

  Logical_Operator_out1980_out1 <= Logical_Operator_out1468_out1 XOR Logical_Operator_out1472_out1;

  Logical_Operator_out1981_out1 <= Logical_Operator_out955_out1 XOR Logical_Operator_out959_out1;

  Logical_Operator_out1982_out1 <= Logical_Operator_out956_out1 XOR Logical_Operator_out960_out1;

  Logical_Operator_out1983_out1 <= Logical_Operator_out444_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out1984_out1 <= in888 XOR in896;

  Logical_Operator_out1985_out1 <= Logical_Operator_out1473_out1 XOR Logical_Operator_out1477_out1;

  Logical_Operator_out1986_out1 <= Logical_Operator_out1474_out1 XOR Logical_Operator_out1478_out1;

  Logical_Operator_out1987_out1 <= Logical_Operator_out1475_out1 XOR Logical_Operator_out1479_out1;

  Logical_Operator_out1988_out1 <= Logical_Operator_out1476_out1 XOR Logical_Operator_out1480_out1;

  Logical_Operator_out1989_out1 <= Logical_Operator_out963_out1 XOR Logical_Operator_out967_out1;

  Logical_Operator_out1990_out1 <= Logical_Operator_out964_out1 XOR Logical_Operator_out968_out1;

  Logical_Operator_out1991_out1 <= Logical_Operator_out452_out1 XOR Logical_Operator_out456_out1;

  Logical_Operator_out1992_out1 <= in904 XOR in912;

  Logical_Operator_out1993_out1 <= Logical_Operator_out1481_out1 XOR Logical_Operator_out1485_out1;

  Logical_Operator_out1994_out1 <= Logical_Operator_out1482_out1 XOR Logical_Operator_out1486_out1;

  Logical_Operator_out1995_out1 <= Logical_Operator_out1483_out1 XOR Logical_Operator_out1487_out1;

  Logical_Operator_out1996_out1 <= Logical_Operator_out1484_out1 XOR Logical_Operator_out1488_out1;

  Logical_Operator_out1997_out1 <= Logical_Operator_out971_out1 XOR Logical_Operator_out975_out1;

  Logical_Operator_out1998_out1 <= Logical_Operator_out972_out1 XOR Logical_Operator_out976_out1;

  Logical_Operator_out1999_out1 <= Logical_Operator_out460_out1 XOR Logical_Operator_out464_out1;

  Logical_Operator_out2000_out1 <= in920 XOR in928;

  Logical_Operator_out2001_out1 <= Logical_Operator_out1489_out1 XOR Logical_Operator_out1493_out1;

  Logical_Operator_out2002_out1 <= Logical_Operator_out1490_out1 XOR Logical_Operator_out1494_out1;

  Logical_Operator_out2003_out1 <= Logical_Operator_out1491_out1 XOR Logical_Operator_out1495_out1;

  Logical_Operator_out2004_out1 <= Logical_Operator_out1492_out1 XOR Logical_Operator_out1496_out1;

  Logical_Operator_out2005_out1 <= Logical_Operator_out979_out1 XOR Logical_Operator_out983_out1;

  Logical_Operator_out2006_out1 <= Logical_Operator_out980_out1 XOR Logical_Operator_out984_out1;

  Logical_Operator_out2007_out1 <= Logical_Operator_out468_out1 XOR Logical_Operator_out472_out1;

  Logical_Operator_out2008_out1 <= in936 XOR in944;

  Logical_Operator_out2009_out1 <= Logical_Operator_out1497_out1 XOR Logical_Operator_out1501_out1;

  Logical_Operator_out2010_out1 <= Logical_Operator_out1498_out1 XOR Logical_Operator_out1502_out1;

  Logical_Operator_out2011_out1 <= Logical_Operator_out1499_out1 XOR Logical_Operator_out1503_out1;

  Logical_Operator_out2012_out1 <= Logical_Operator_out1500_out1 XOR Logical_Operator_out1504_out1;

  Logical_Operator_out2013_out1 <= Logical_Operator_out987_out1 XOR Logical_Operator_out991_out1;

  Logical_Operator_out2014_out1 <= Logical_Operator_out988_out1 XOR Logical_Operator_out992_out1;

  Logical_Operator_out2015_out1 <= Logical_Operator_out476_out1 XOR Logical_Operator_out480_out1;

  Logical_Operator_out2016_out1 <= in952 XOR in960;

  Logical_Operator_out2017_out1 <= Logical_Operator_out1505_out1 XOR Logical_Operator_out1509_out1;

  Logical_Operator_out2018_out1 <= Logical_Operator_out1506_out1 XOR Logical_Operator_out1510_out1;

  Logical_Operator_out2019_out1 <= Logical_Operator_out1507_out1 XOR Logical_Operator_out1511_out1;

  Logical_Operator_out2020_out1 <= Logical_Operator_out1508_out1 XOR Logical_Operator_out1512_out1;

  Logical_Operator_out2021_out1 <= Logical_Operator_out995_out1 XOR Logical_Operator_out999_out1;

  Logical_Operator_out2022_out1 <= Logical_Operator_out996_out1 XOR Logical_Operator_out1000_out1;

  Logical_Operator_out2023_out1 <= Logical_Operator_out484_out1 XOR Logical_Operator_out488_out1;

  Logical_Operator_out2024_out1 <= in968 XOR in976;

  Logical_Operator_out2025_out1 <= Logical_Operator_out1513_out1 XOR Logical_Operator_out1517_out1;

  Logical_Operator_out2026_out1 <= Logical_Operator_out1514_out1 XOR Logical_Operator_out1518_out1;

  Logical_Operator_out2027_out1 <= Logical_Operator_out1515_out1 XOR Logical_Operator_out1519_out1;

  Logical_Operator_out2028_out1 <= Logical_Operator_out1516_out1 XOR Logical_Operator_out1520_out1;

  Logical_Operator_out2029_out1 <= Logical_Operator_out1003_out1 XOR Logical_Operator_out1007_out1;

  Logical_Operator_out2030_out1 <= Logical_Operator_out1004_out1 XOR Logical_Operator_out1008_out1;

  Logical_Operator_out2031_out1 <= Logical_Operator_out492_out1 XOR Logical_Operator_out496_out1;

  Logical_Operator_out2032_out1 <= in984 XOR in992;

  Logical_Operator_out2033_out1 <= Logical_Operator_out1521_out1 XOR Logical_Operator_out1525_out1;

  Logical_Operator_out2034_out1 <= Logical_Operator_out1522_out1 XOR Logical_Operator_out1526_out1;

  Logical_Operator_out2035_out1 <= Logical_Operator_out1523_out1 XOR Logical_Operator_out1527_out1;

  Logical_Operator_out2036_out1 <= Logical_Operator_out1524_out1 XOR Logical_Operator_out1528_out1;

  Logical_Operator_out2037_out1 <= Logical_Operator_out1011_out1 XOR Logical_Operator_out1015_out1;

  Logical_Operator_out2038_out1 <= Logical_Operator_out1012_out1 XOR Logical_Operator_out1016_out1;

  Logical_Operator_out2039_out1 <= Logical_Operator_out500_out1 XOR Logical_Operator_out504_out1;

  Logical_Operator_out2040_out1 <= in1000 XOR in1008;

  Logical_Operator_out2041_out1 <= Logical_Operator_out1529_out1 XOR Logical_Operator_out1533_out1;

  Logical_Operator_out2042_out1 <= Logical_Operator_out1530_out1 XOR Logical_Operator_out1534_out1;

  Logical_Operator_out2043_out1 <= Logical_Operator_out1531_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out2044_out1 <= Logical_Operator_out1532_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out2045_out1 <= Logical_Operator_out1019_out1 XOR Logical_Operator_out1023_out1;

  Logical_Operator_out2046_out1 <= Logical_Operator_out1020_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out2047_out1 <= Logical_Operator_out508_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out2048_out1 <= in1016 XOR in1024;

  Logical_Operator_out2049_out1 <= Logical_Operator_out1537_out1 XOR Logical_Operator_out1545_out1;

  Logical_Operator_out2050_out1 <= Logical_Operator_out1538_out1 XOR Logical_Operator_out1546_out1;

  Logical_Operator_out2051_out1 <= Logical_Operator_out1539_out1 XOR Logical_Operator_out1547_out1;

  Logical_Operator_out2052_out1 <= Logical_Operator_out1540_out1 XOR Logical_Operator_out1548_out1;

  Logical_Operator_out2053_out1 <= Logical_Operator_out1541_out1 XOR Logical_Operator_out1549_out1;

  Logical_Operator_out2054_out1 <= Logical_Operator_out1542_out1 XOR Logical_Operator_out1550_out1;

  Logical_Operator_out2055_out1 <= Logical_Operator_out1543_out1 XOR Logical_Operator_out1551_out1;

  Logical_Operator_out2056_out1 <= Logical_Operator_out1544_out1 XOR Logical_Operator_out1552_out1;

  Logical_Operator_out2057_out1 <= Logical_Operator_out1029_out1 XOR Logical_Operator_out1037_out1;

  Logical_Operator_out2058_out1 <= Logical_Operator_out1030_out1 XOR Logical_Operator_out1038_out1;

  Logical_Operator_out2059_out1 <= Logical_Operator_out1031_out1 XOR Logical_Operator_out1039_out1;

  Logical_Operator_out2060_out1 <= Logical_Operator_out1032_out1 XOR Logical_Operator_out1040_out1;

  Logical_Operator_out2061_out1 <= Logical_Operator_out519_out1 XOR Logical_Operator_out527_out1;

  Logical_Operator_out2062_out1 <= Logical_Operator_out520_out1 XOR Logical_Operator_out528_out1;

  Logical_Operator_out2063_out1 <= Logical_Operator_out8_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out2064_out1 <= in16 XOR in32;

  Logical_Operator_out2065_out1 <= Logical_Operator_out1553_out1 XOR Logical_Operator_out1561_out1;

  Logical_Operator_out2066_out1 <= Logical_Operator_out1554_out1 XOR Logical_Operator_out1562_out1;

  Logical_Operator_out2067_out1 <= Logical_Operator_out1555_out1 XOR Logical_Operator_out1563_out1;

  Logical_Operator_out2068_out1 <= Logical_Operator_out1556_out1 XOR Logical_Operator_out1564_out1;

  Logical_Operator_out2069_out1 <= Logical_Operator_out1557_out1 XOR Logical_Operator_out1565_out1;

  Logical_Operator_out2070_out1 <= Logical_Operator_out1558_out1 XOR Logical_Operator_out1566_out1;

  Logical_Operator_out2071_out1 <= Logical_Operator_out1559_out1 XOR Logical_Operator_out1567_out1;

  Logical_Operator_out2072_out1 <= Logical_Operator_out1560_out1 XOR Logical_Operator_out1568_out1;

  Logical_Operator_out2073_out1 <= Logical_Operator_out1045_out1 XOR Logical_Operator_out1053_out1;

  Logical_Operator_out2074_out1 <= Logical_Operator_out1046_out1 XOR Logical_Operator_out1054_out1;

  Logical_Operator_out2075_out1 <= Logical_Operator_out1047_out1 XOR Logical_Operator_out1055_out1;

  Logical_Operator_out2076_out1 <= Logical_Operator_out1048_out1 XOR Logical_Operator_out1056_out1;

  Logical_Operator_out2077_out1 <= Logical_Operator_out535_out1 XOR Logical_Operator_out543_out1;

  Logical_Operator_out2078_out1 <= Logical_Operator_out536_out1 XOR Logical_Operator_out544_out1;

  Logical_Operator_out2079_out1 <= Logical_Operator_out24_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out2080_out1 <= in48 XOR in64;

  Logical_Operator_out2081_out1 <= Logical_Operator_out1569_out1 XOR Logical_Operator_out1577_out1;

  Logical_Operator_out2082_out1 <= Logical_Operator_out1570_out1 XOR Logical_Operator_out1578_out1;

  Logical_Operator_out2083_out1 <= Logical_Operator_out1571_out1 XOR Logical_Operator_out1579_out1;

  Logical_Operator_out2084_out1 <= Logical_Operator_out1572_out1 XOR Logical_Operator_out1580_out1;

  Logical_Operator_out2085_out1 <= Logical_Operator_out1573_out1 XOR Logical_Operator_out1581_out1;

  Logical_Operator_out2086_out1 <= Logical_Operator_out1574_out1 XOR Logical_Operator_out1582_out1;

  Logical_Operator_out2087_out1 <= Logical_Operator_out1575_out1 XOR Logical_Operator_out1583_out1;

  Logical_Operator_out2088_out1 <= Logical_Operator_out1576_out1 XOR Logical_Operator_out1584_out1;

  Logical_Operator_out2089_out1 <= Logical_Operator_out1061_out1 XOR Logical_Operator_out1069_out1;

  Logical_Operator_out2090_out1 <= Logical_Operator_out1062_out1 XOR Logical_Operator_out1070_out1;

  Logical_Operator_out2091_out1 <= Logical_Operator_out1063_out1 XOR Logical_Operator_out1071_out1;

  Logical_Operator_out2092_out1 <= Logical_Operator_out1064_out1 XOR Logical_Operator_out1072_out1;

  Logical_Operator_out2093_out1 <= Logical_Operator_out551_out1 XOR Logical_Operator_out559_out1;

  Logical_Operator_out2094_out1 <= Logical_Operator_out552_out1 XOR Logical_Operator_out560_out1;

  Logical_Operator_out2095_out1 <= Logical_Operator_out40_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out2096_out1 <= in80 XOR in96;

  Logical_Operator_out2097_out1 <= Logical_Operator_out1585_out1 XOR Logical_Operator_out1593_out1;

  Logical_Operator_out2098_out1 <= Logical_Operator_out1586_out1 XOR Logical_Operator_out1594_out1;

  Logical_Operator_out2099_out1 <= Logical_Operator_out1587_out1 XOR Logical_Operator_out1595_out1;

  Logical_Operator_out2100_out1 <= Logical_Operator_out1588_out1 XOR Logical_Operator_out1596_out1;

  Logical_Operator_out2101_out1 <= Logical_Operator_out1589_out1 XOR Logical_Operator_out1597_out1;

  Logical_Operator_out2102_out1 <= Logical_Operator_out1590_out1 XOR Logical_Operator_out1598_out1;

  Logical_Operator_out2103_out1 <= Logical_Operator_out1591_out1 XOR Logical_Operator_out1599_out1;

  Logical_Operator_out2104_out1 <= Logical_Operator_out1592_out1 XOR Logical_Operator_out1600_out1;

  Logical_Operator_out2105_out1 <= Logical_Operator_out1077_out1 XOR Logical_Operator_out1085_out1;

  Logical_Operator_out2106_out1 <= Logical_Operator_out1078_out1 XOR Logical_Operator_out1086_out1;

  Logical_Operator_out2107_out1 <= Logical_Operator_out1079_out1 XOR Logical_Operator_out1087_out1;

  Logical_Operator_out2108_out1 <= Logical_Operator_out1080_out1 XOR Logical_Operator_out1088_out1;

  Logical_Operator_out2109_out1 <= Logical_Operator_out567_out1 XOR Logical_Operator_out575_out1;

  Logical_Operator_out2110_out1 <= Logical_Operator_out568_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out2111_out1 <= Logical_Operator_out56_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out2112_out1 <= in112 XOR in128;

  Logical_Operator_out2113_out1 <= Logical_Operator_out1601_out1 XOR Logical_Operator_out1609_out1;

  Logical_Operator_out2114_out1 <= Logical_Operator_out1602_out1 XOR Logical_Operator_out1610_out1;

  Logical_Operator_out2115_out1 <= Logical_Operator_out1603_out1 XOR Logical_Operator_out1611_out1;

  Logical_Operator_out2116_out1 <= Logical_Operator_out1604_out1 XOR Logical_Operator_out1612_out1;

  Logical_Operator_out2117_out1 <= Logical_Operator_out1605_out1 XOR Logical_Operator_out1613_out1;

  Logical_Operator_out2118_out1 <= Logical_Operator_out1606_out1 XOR Logical_Operator_out1614_out1;

  Logical_Operator_out2119_out1 <= Logical_Operator_out1607_out1 XOR Logical_Operator_out1615_out1;

  Logical_Operator_out2120_out1 <= Logical_Operator_out1608_out1 XOR Logical_Operator_out1616_out1;

  Logical_Operator_out2121_out1 <= Logical_Operator_out1093_out1 XOR Logical_Operator_out1101_out1;

  Logical_Operator_out2122_out1 <= Logical_Operator_out1094_out1 XOR Logical_Operator_out1102_out1;

  Logical_Operator_out2123_out1 <= Logical_Operator_out1095_out1 XOR Logical_Operator_out1103_out1;

  Logical_Operator_out2124_out1 <= Logical_Operator_out1096_out1 XOR Logical_Operator_out1104_out1;

  Logical_Operator_out2125_out1 <= Logical_Operator_out583_out1 XOR Logical_Operator_out591_out1;

  Logical_Operator_out2126_out1 <= Logical_Operator_out584_out1 XOR Logical_Operator_out592_out1;

  Logical_Operator_out2127_out1 <= Logical_Operator_out72_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out2128_out1 <= in144 XOR in160;

  Logical_Operator_out2129_out1 <= Logical_Operator_out1617_out1 XOR Logical_Operator_out1625_out1;

  Logical_Operator_out2130_out1 <= Logical_Operator_out1618_out1 XOR Logical_Operator_out1626_out1;

  Logical_Operator_out2131_out1 <= Logical_Operator_out1619_out1 XOR Logical_Operator_out1627_out1;

  Logical_Operator_out2132_out1 <= Logical_Operator_out1620_out1 XOR Logical_Operator_out1628_out1;

  Logical_Operator_out2133_out1 <= Logical_Operator_out1621_out1 XOR Logical_Operator_out1629_out1;

  Logical_Operator_out2134_out1 <= Logical_Operator_out1622_out1 XOR Logical_Operator_out1630_out1;

  Logical_Operator_out2135_out1 <= Logical_Operator_out1623_out1 XOR Logical_Operator_out1631_out1;

  Logical_Operator_out2136_out1 <= Logical_Operator_out1624_out1 XOR Logical_Operator_out1632_out1;

  Logical_Operator_out2137_out1 <= Logical_Operator_out1109_out1 XOR Logical_Operator_out1117_out1;

  Logical_Operator_out2138_out1 <= Logical_Operator_out1110_out1 XOR Logical_Operator_out1118_out1;

  Logical_Operator_out2139_out1 <= Logical_Operator_out1111_out1 XOR Logical_Operator_out1119_out1;

  Logical_Operator_out2140_out1 <= Logical_Operator_out1112_out1 XOR Logical_Operator_out1120_out1;

  Logical_Operator_out2141_out1 <= Logical_Operator_out599_out1 XOR Logical_Operator_out607_out1;

  Logical_Operator_out2142_out1 <= Logical_Operator_out600_out1 XOR Logical_Operator_out608_out1;

  Logical_Operator_out2143_out1 <= Logical_Operator_out88_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out2144_out1 <= in176 XOR in192;

  Logical_Operator_out2145_out1 <= Logical_Operator_out1633_out1 XOR Logical_Operator_out1641_out1;

  Logical_Operator_out2146_out1 <= Logical_Operator_out1634_out1 XOR Logical_Operator_out1642_out1;

  Logical_Operator_out2147_out1 <= Logical_Operator_out1635_out1 XOR Logical_Operator_out1643_out1;

  Logical_Operator_out2148_out1 <= Logical_Operator_out1636_out1 XOR Logical_Operator_out1644_out1;

  Logical_Operator_out2149_out1 <= Logical_Operator_out1637_out1 XOR Logical_Operator_out1645_out1;

  Logical_Operator_out2150_out1 <= Logical_Operator_out1638_out1 XOR Logical_Operator_out1646_out1;

  Logical_Operator_out2151_out1 <= Logical_Operator_out1639_out1 XOR Logical_Operator_out1647_out1;

  Logical_Operator_out2152_out1 <= Logical_Operator_out1640_out1 XOR Logical_Operator_out1648_out1;

  Logical_Operator_out2153_out1 <= Logical_Operator_out1125_out1 XOR Logical_Operator_out1133_out1;

  Logical_Operator_out2154_out1 <= Logical_Operator_out1126_out1 XOR Logical_Operator_out1134_out1;

  Logical_Operator_out2155_out1 <= Logical_Operator_out1127_out1 XOR Logical_Operator_out1135_out1;

  Logical_Operator_out2156_out1 <= Logical_Operator_out1128_out1 XOR Logical_Operator_out1136_out1;

  Logical_Operator_out2157_out1 <= Logical_Operator_out615_out1 XOR Logical_Operator_out623_out1;

  Logical_Operator_out2158_out1 <= Logical_Operator_out616_out1 XOR Logical_Operator_out624_out1;

  Logical_Operator_out2159_out1 <= Logical_Operator_out104_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out2160_out1 <= in208 XOR in224;

  Logical_Operator_out2161_out1 <= Logical_Operator_out1649_out1 XOR Logical_Operator_out1657_out1;

  Logical_Operator_out2162_out1 <= Logical_Operator_out1650_out1 XOR Logical_Operator_out1658_out1;

  Logical_Operator_out2163_out1 <= Logical_Operator_out1651_out1 XOR Logical_Operator_out1659_out1;

  Logical_Operator_out2164_out1 <= Logical_Operator_out1652_out1 XOR Logical_Operator_out1660_out1;

  Logical_Operator_out2165_out1 <= Logical_Operator_out1653_out1 XOR Logical_Operator_out1661_out1;

  Logical_Operator_out2166_out1 <= Logical_Operator_out1654_out1 XOR Logical_Operator_out1662_out1;

  Logical_Operator_out2167_out1 <= Logical_Operator_out1655_out1 XOR Logical_Operator_out1663_out1;

  Logical_Operator_out2168_out1 <= Logical_Operator_out1656_out1 XOR Logical_Operator_out1664_out1;

  Logical_Operator_out2169_out1 <= Logical_Operator_out1141_out1 XOR Logical_Operator_out1149_out1;

  Logical_Operator_out2170_out1 <= Logical_Operator_out1142_out1 XOR Logical_Operator_out1150_out1;

  Logical_Operator_out2171_out1 <= Logical_Operator_out1143_out1 XOR Logical_Operator_out1151_out1;

  Logical_Operator_out2172_out1 <= Logical_Operator_out1144_out1 XOR Logical_Operator_out1152_out1;

  Logical_Operator_out2173_out1 <= Logical_Operator_out631_out1 XOR Logical_Operator_out639_out1;

  Logical_Operator_out2174_out1 <= Logical_Operator_out632_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out2175_out1 <= Logical_Operator_out120_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out2176_out1 <= in240 XOR in256;

  Logical_Operator_out2177_out1 <= Logical_Operator_out1665_out1 XOR Logical_Operator_out1673_out1;

  Logical_Operator_out2178_out1 <= Logical_Operator_out1666_out1 XOR Logical_Operator_out1674_out1;

  Logical_Operator_out2179_out1 <= Logical_Operator_out1667_out1 XOR Logical_Operator_out1675_out1;

  Logical_Operator_out2180_out1 <= Logical_Operator_out1668_out1 XOR Logical_Operator_out1676_out1;

  Logical_Operator_out2181_out1 <= Logical_Operator_out1669_out1 XOR Logical_Operator_out1677_out1;

  Logical_Operator_out2182_out1 <= Logical_Operator_out1670_out1 XOR Logical_Operator_out1678_out1;

  Logical_Operator_out2183_out1 <= Logical_Operator_out1671_out1 XOR Logical_Operator_out1679_out1;

  Logical_Operator_out2184_out1 <= Logical_Operator_out1672_out1 XOR Logical_Operator_out1680_out1;

  Logical_Operator_out2185_out1 <= Logical_Operator_out1157_out1 XOR Logical_Operator_out1165_out1;

  Logical_Operator_out2186_out1 <= Logical_Operator_out1158_out1 XOR Logical_Operator_out1166_out1;

  Logical_Operator_out2187_out1 <= Logical_Operator_out1159_out1 XOR Logical_Operator_out1167_out1;

  Logical_Operator_out2188_out1 <= Logical_Operator_out1160_out1 XOR Logical_Operator_out1168_out1;

  Logical_Operator_out2189_out1 <= Logical_Operator_out647_out1 XOR Logical_Operator_out655_out1;

  Logical_Operator_out2190_out1 <= Logical_Operator_out648_out1 XOR Logical_Operator_out656_out1;

  Logical_Operator_out2191_out1 <= Logical_Operator_out136_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out2192_out1 <= in272 XOR in288;

  Logical_Operator_out2193_out1 <= Logical_Operator_out1681_out1 XOR Logical_Operator_out1689_out1;

  Logical_Operator_out2194_out1 <= Logical_Operator_out1682_out1 XOR Logical_Operator_out1690_out1;

  Logical_Operator_out2195_out1 <= Logical_Operator_out1683_out1 XOR Logical_Operator_out1691_out1;

  Logical_Operator_out2196_out1 <= Logical_Operator_out1684_out1 XOR Logical_Operator_out1692_out1;

  Logical_Operator_out2197_out1 <= Logical_Operator_out1685_out1 XOR Logical_Operator_out1693_out1;

  Logical_Operator_out2198_out1 <= Logical_Operator_out1686_out1 XOR Logical_Operator_out1694_out1;

  Logical_Operator_out2199_out1 <= Logical_Operator_out1687_out1 XOR Logical_Operator_out1695_out1;

  Logical_Operator_out2200_out1 <= Logical_Operator_out1688_out1 XOR Logical_Operator_out1696_out1;

  Logical_Operator_out2201_out1 <= Logical_Operator_out1173_out1 XOR Logical_Operator_out1181_out1;

  Logical_Operator_out2202_out1 <= Logical_Operator_out1174_out1 XOR Logical_Operator_out1182_out1;

  Logical_Operator_out2203_out1 <= Logical_Operator_out1175_out1 XOR Logical_Operator_out1183_out1;

  Logical_Operator_out2204_out1 <= Logical_Operator_out1176_out1 XOR Logical_Operator_out1184_out1;

  Logical_Operator_out2205_out1 <= Logical_Operator_out663_out1 XOR Logical_Operator_out671_out1;

  Logical_Operator_out2206_out1 <= Logical_Operator_out664_out1 XOR Logical_Operator_out672_out1;

  Logical_Operator_out2207_out1 <= Logical_Operator_out152_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out2208_out1 <= in304 XOR in320;

  Logical_Operator_out2209_out1 <= Logical_Operator_out1697_out1 XOR Logical_Operator_out1705_out1;

  Logical_Operator_out2210_out1 <= Logical_Operator_out1698_out1 XOR Logical_Operator_out1706_out1;

  Logical_Operator_out2211_out1 <= Logical_Operator_out1699_out1 XOR Logical_Operator_out1707_out1;

  Logical_Operator_out2212_out1 <= Logical_Operator_out1700_out1 XOR Logical_Operator_out1708_out1;

  Logical_Operator_out2213_out1 <= Logical_Operator_out1701_out1 XOR Logical_Operator_out1709_out1;

  Logical_Operator_out2214_out1 <= Logical_Operator_out1702_out1 XOR Logical_Operator_out1710_out1;

  Logical_Operator_out2215_out1 <= Logical_Operator_out1703_out1 XOR Logical_Operator_out1711_out1;

  Logical_Operator_out2216_out1 <= Logical_Operator_out1704_out1 XOR Logical_Operator_out1712_out1;

  Logical_Operator_out2217_out1 <= Logical_Operator_out1189_out1 XOR Logical_Operator_out1197_out1;

  Logical_Operator_out2218_out1 <= Logical_Operator_out1190_out1 XOR Logical_Operator_out1198_out1;

  Logical_Operator_out2219_out1 <= Logical_Operator_out1191_out1 XOR Logical_Operator_out1199_out1;

  Logical_Operator_out2220_out1 <= Logical_Operator_out1192_out1 XOR Logical_Operator_out1200_out1;

  Logical_Operator_out2221_out1 <= Logical_Operator_out679_out1 XOR Logical_Operator_out687_out1;

  Logical_Operator_out2222_out1 <= Logical_Operator_out680_out1 XOR Logical_Operator_out688_out1;

  Logical_Operator_out2223_out1 <= Logical_Operator_out168_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out2224_out1 <= in336 XOR in352;

  Logical_Operator_out2225_out1 <= Logical_Operator_out1713_out1 XOR Logical_Operator_out1721_out1;

  Logical_Operator_out2226_out1 <= Logical_Operator_out1714_out1 XOR Logical_Operator_out1722_out1;

  Logical_Operator_out2227_out1 <= Logical_Operator_out1715_out1 XOR Logical_Operator_out1723_out1;

  Logical_Operator_out2228_out1 <= Logical_Operator_out1716_out1 XOR Logical_Operator_out1724_out1;

  Logical_Operator_out2229_out1 <= Logical_Operator_out1717_out1 XOR Logical_Operator_out1725_out1;

  Logical_Operator_out2230_out1 <= Logical_Operator_out1718_out1 XOR Logical_Operator_out1726_out1;

  Logical_Operator_out2231_out1 <= Logical_Operator_out1719_out1 XOR Logical_Operator_out1727_out1;

  Logical_Operator_out2232_out1 <= Logical_Operator_out1720_out1 XOR Logical_Operator_out1728_out1;

  Logical_Operator_out2233_out1 <= Logical_Operator_out1205_out1 XOR Logical_Operator_out1213_out1;

  Logical_Operator_out2234_out1 <= Logical_Operator_out1206_out1 XOR Logical_Operator_out1214_out1;

  Logical_Operator_out2235_out1 <= Logical_Operator_out1207_out1 XOR Logical_Operator_out1215_out1;

  Logical_Operator_out2236_out1 <= Logical_Operator_out1208_out1 XOR Logical_Operator_out1216_out1;

  Logical_Operator_out2237_out1 <= Logical_Operator_out695_out1 XOR Logical_Operator_out703_out1;

  Logical_Operator_out2238_out1 <= Logical_Operator_out696_out1 XOR Logical_Operator_out704_out1;

  Logical_Operator_out2239_out1 <= Logical_Operator_out184_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out2240_out1 <= in368 XOR in384;

  Logical_Operator_out2241_out1 <= Logical_Operator_out1729_out1 XOR Logical_Operator_out1737_out1;

  Logical_Operator_out2242_out1 <= Logical_Operator_out1730_out1 XOR Logical_Operator_out1738_out1;

  Logical_Operator_out2243_out1 <= Logical_Operator_out1731_out1 XOR Logical_Operator_out1739_out1;

  Logical_Operator_out2244_out1 <= Logical_Operator_out1732_out1 XOR Logical_Operator_out1740_out1;

  Logical_Operator_out2245_out1 <= Logical_Operator_out1733_out1 XOR Logical_Operator_out1741_out1;

  Logical_Operator_out2246_out1 <= Logical_Operator_out1734_out1 XOR Logical_Operator_out1742_out1;

  Logical_Operator_out2247_out1 <= Logical_Operator_out1735_out1 XOR Logical_Operator_out1743_out1;

  Logical_Operator_out2248_out1 <= Logical_Operator_out1736_out1 XOR Logical_Operator_out1744_out1;

  Logical_Operator_out2249_out1 <= Logical_Operator_out1221_out1 XOR Logical_Operator_out1229_out1;

  Logical_Operator_out2250_out1 <= Logical_Operator_out1222_out1 XOR Logical_Operator_out1230_out1;

  Logical_Operator_out2251_out1 <= Logical_Operator_out1223_out1 XOR Logical_Operator_out1231_out1;

  Logical_Operator_out2252_out1 <= Logical_Operator_out1224_out1 XOR Logical_Operator_out1232_out1;

  Logical_Operator_out2253_out1 <= Logical_Operator_out711_out1 XOR Logical_Operator_out719_out1;

  Logical_Operator_out2254_out1 <= Logical_Operator_out712_out1 XOR Logical_Operator_out720_out1;

  Logical_Operator_out2255_out1 <= Logical_Operator_out200_out1 XOR Logical_Operator_out208_out1;

  Logical_Operator_out2256_out1 <= in400 XOR in416;

  Logical_Operator_out2257_out1 <= Logical_Operator_out1745_out1 XOR Logical_Operator_out1753_out1;

  Logical_Operator_out2258_out1 <= Logical_Operator_out1746_out1 XOR Logical_Operator_out1754_out1;

  Logical_Operator_out2259_out1 <= Logical_Operator_out1747_out1 XOR Logical_Operator_out1755_out1;

  Logical_Operator_out2260_out1 <= Logical_Operator_out1748_out1 XOR Logical_Operator_out1756_out1;

  Logical_Operator_out2261_out1 <= Logical_Operator_out1749_out1 XOR Logical_Operator_out1757_out1;

  Logical_Operator_out2262_out1 <= Logical_Operator_out1750_out1 XOR Logical_Operator_out1758_out1;

  Logical_Operator_out2263_out1 <= Logical_Operator_out1751_out1 XOR Logical_Operator_out1759_out1;

  Logical_Operator_out2264_out1 <= Logical_Operator_out1752_out1 XOR Logical_Operator_out1760_out1;

  Logical_Operator_out2265_out1 <= Logical_Operator_out1237_out1 XOR Logical_Operator_out1245_out1;

  Logical_Operator_out2266_out1 <= Logical_Operator_out1238_out1 XOR Logical_Operator_out1246_out1;

  Logical_Operator_out2267_out1 <= Logical_Operator_out1239_out1 XOR Logical_Operator_out1247_out1;

  Logical_Operator_out2268_out1 <= Logical_Operator_out1240_out1 XOR Logical_Operator_out1248_out1;

  Logical_Operator_out2269_out1 <= Logical_Operator_out727_out1 XOR Logical_Operator_out735_out1;

  Logical_Operator_out2270_out1 <= Logical_Operator_out728_out1 XOR Logical_Operator_out736_out1;

  Logical_Operator_out2271_out1 <= Logical_Operator_out216_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out2272_out1 <= in432 XOR in448;

  Logical_Operator_out2273_out1 <= Logical_Operator_out1761_out1 XOR Logical_Operator_out1769_out1;

  Logical_Operator_out2274_out1 <= Logical_Operator_out1762_out1 XOR Logical_Operator_out1770_out1;

  Logical_Operator_out2275_out1 <= Logical_Operator_out1763_out1 XOR Logical_Operator_out1771_out1;

  Logical_Operator_out2276_out1 <= Logical_Operator_out1764_out1 XOR Logical_Operator_out1772_out1;

  Logical_Operator_out2277_out1 <= Logical_Operator_out1765_out1 XOR Logical_Operator_out1773_out1;

  Logical_Operator_out2278_out1 <= Logical_Operator_out1766_out1 XOR Logical_Operator_out1774_out1;

  Logical_Operator_out2279_out1 <= Logical_Operator_out1767_out1 XOR Logical_Operator_out1775_out1;

  Logical_Operator_out2280_out1 <= Logical_Operator_out1768_out1 XOR Logical_Operator_out1776_out1;

  Logical_Operator_out2281_out1 <= Logical_Operator_out1253_out1 XOR Logical_Operator_out1261_out1;

  Logical_Operator_out2282_out1 <= Logical_Operator_out1254_out1 XOR Logical_Operator_out1262_out1;

  Logical_Operator_out2283_out1 <= Logical_Operator_out1255_out1 XOR Logical_Operator_out1263_out1;

  Logical_Operator_out2284_out1 <= Logical_Operator_out1256_out1 XOR Logical_Operator_out1264_out1;

  Logical_Operator_out2285_out1 <= Logical_Operator_out743_out1 XOR Logical_Operator_out751_out1;

  Logical_Operator_out2286_out1 <= Logical_Operator_out744_out1 XOR Logical_Operator_out752_out1;

  Logical_Operator_out2287_out1 <= Logical_Operator_out232_out1 XOR Logical_Operator_out240_out1;

  Logical_Operator_out2288_out1 <= in464 XOR in480;

  Logical_Operator_out2289_out1 <= Logical_Operator_out1777_out1 XOR Logical_Operator_out1785_out1;

  Logical_Operator_out2290_out1 <= Logical_Operator_out1778_out1 XOR Logical_Operator_out1786_out1;

  Logical_Operator_out2291_out1 <= Logical_Operator_out1779_out1 XOR Logical_Operator_out1787_out1;

  Logical_Operator_out2292_out1 <= Logical_Operator_out1780_out1 XOR Logical_Operator_out1788_out1;

  Logical_Operator_out2293_out1 <= Logical_Operator_out1781_out1 XOR Logical_Operator_out1789_out1;

  Logical_Operator_out2294_out1 <= Logical_Operator_out1782_out1 XOR Logical_Operator_out1790_out1;

  Logical_Operator_out2295_out1 <= Logical_Operator_out1783_out1 XOR Logical_Operator_out1791_out1;

  Logical_Operator_out2296_out1 <= Logical_Operator_out1784_out1 XOR Logical_Operator_out1792_out1;

  Logical_Operator_out2297_out1 <= Logical_Operator_out1269_out1 XOR Logical_Operator_out1277_out1;

  Logical_Operator_out2298_out1 <= Logical_Operator_out1270_out1 XOR Logical_Operator_out1278_out1;

  Logical_Operator_out2299_out1 <= Logical_Operator_out1271_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out2300_out1 <= Logical_Operator_out1272_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out2301_out1 <= Logical_Operator_out759_out1 XOR Logical_Operator_out767_out1;

  Logical_Operator_out2302_out1 <= Logical_Operator_out760_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out2303_out1 <= Logical_Operator_out248_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out2304_out1 <= in496 XOR in512;

  Logical_Operator_out2305_out1 <= Logical_Operator_out1793_out1 XOR Logical_Operator_out1801_out1;

  Logical_Operator_out2306_out1 <= Logical_Operator_out1794_out1 XOR Logical_Operator_out1802_out1;

  Logical_Operator_out2307_out1 <= Logical_Operator_out1795_out1 XOR Logical_Operator_out1803_out1;

  Logical_Operator_out2308_out1 <= Logical_Operator_out1796_out1 XOR Logical_Operator_out1804_out1;

  Logical_Operator_out2309_out1 <= Logical_Operator_out1797_out1 XOR Logical_Operator_out1805_out1;

  Logical_Operator_out2310_out1 <= Logical_Operator_out1798_out1 XOR Logical_Operator_out1806_out1;

  Logical_Operator_out2311_out1 <= Logical_Operator_out1799_out1 XOR Logical_Operator_out1807_out1;

  Logical_Operator_out2312_out1 <= Logical_Operator_out1800_out1 XOR Logical_Operator_out1808_out1;

  Logical_Operator_out2313_out1 <= Logical_Operator_out1285_out1 XOR Logical_Operator_out1293_out1;

  Logical_Operator_out2314_out1 <= Logical_Operator_out1286_out1 XOR Logical_Operator_out1294_out1;

  Logical_Operator_out2315_out1 <= Logical_Operator_out1287_out1 XOR Logical_Operator_out1295_out1;

  Logical_Operator_out2316_out1 <= Logical_Operator_out1288_out1 XOR Logical_Operator_out1296_out1;

  Logical_Operator_out2317_out1 <= Logical_Operator_out775_out1 XOR Logical_Operator_out783_out1;

  Logical_Operator_out2318_out1 <= Logical_Operator_out776_out1 XOR Logical_Operator_out784_out1;

  Logical_Operator_out2319_out1 <= Logical_Operator_out264_out1 XOR Logical_Operator_out272_out1;

  Logical_Operator_out2320_out1 <= in528 XOR in544;

  Logical_Operator_out2321_out1 <= Logical_Operator_out1809_out1 XOR Logical_Operator_out1817_out1;

  Logical_Operator_out2322_out1 <= Logical_Operator_out1810_out1 XOR Logical_Operator_out1818_out1;

  Logical_Operator_out2323_out1 <= Logical_Operator_out1811_out1 XOR Logical_Operator_out1819_out1;

  Logical_Operator_out2324_out1 <= Logical_Operator_out1812_out1 XOR Logical_Operator_out1820_out1;

  Logical_Operator_out2325_out1 <= Logical_Operator_out1813_out1 XOR Logical_Operator_out1821_out1;

  Logical_Operator_out2326_out1 <= Logical_Operator_out1814_out1 XOR Logical_Operator_out1822_out1;

  Logical_Operator_out2327_out1 <= Logical_Operator_out1815_out1 XOR Logical_Operator_out1823_out1;

  Logical_Operator_out2328_out1 <= Logical_Operator_out1816_out1 XOR Logical_Operator_out1824_out1;

  Logical_Operator_out2329_out1 <= Logical_Operator_out1301_out1 XOR Logical_Operator_out1309_out1;

  Logical_Operator_out2330_out1 <= Logical_Operator_out1302_out1 XOR Logical_Operator_out1310_out1;

  Logical_Operator_out2331_out1 <= Logical_Operator_out1303_out1 XOR Logical_Operator_out1311_out1;

  Logical_Operator_out2332_out1 <= Logical_Operator_out1304_out1 XOR Logical_Operator_out1312_out1;

  Logical_Operator_out2333_out1 <= Logical_Operator_out791_out1 XOR Logical_Operator_out799_out1;

  Logical_Operator_out2334_out1 <= Logical_Operator_out792_out1 XOR Logical_Operator_out800_out1;

  Logical_Operator_out2335_out1 <= Logical_Operator_out280_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out2336_out1 <= in560 XOR in576;

  Logical_Operator_out2337_out1 <= Logical_Operator_out1825_out1 XOR Logical_Operator_out1833_out1;

  Logical_Operator_out2338_out1 <= Logical_Operator_out1826_out1 XOR Logical_Operator_out1834_out1;

  Logical_Operator_out2339_out1 <= Logical_Operator_out1827_out1 XOR Logical_Operator_out1835_out1;

  Logical_Operator_out2340_out1 <= Logical_Operator_out1828_out1 XOR Logical_Operator_out1836_out1;

  Logical_Operator_out2341_out1 <= Logical_Operator_out1829_out1 XOR Logical_Operator_out1837_out1;

  Logical_Operator_out2342_out1 <= Logical_Operator_out1830_out1 XOR Logical_Operator_out1838_out1;

  Logical_Operator_out2343_out1 <= Logical_Operator_out1831_out1 XOR Logical_Operator_out1839_out1;

  Logical_Operator_out2344_out1 <= Logical_Operator_out1832_out1 XOR Logical_Operator_out1840_out1;

  Logical_Operator_out2345_out1 <= Logical_Operator_out1317_out1 XOR Logical_Operator_out1325_out1;

  Logical_Operator_out2346_out1 <= Logical_Operator_out1318_out1 XOR Logical_Operator_out1326_out1;

  Logical_Operator_out2347_out1 <= Logical_Operator_out1319_out1 XOR Logical_Operator_out1327_out1;

  Logical_Operator_out2348_out1 <= Logical_Operator_out1320_out1 XOR Logical_Operator_out1328_out1;

  Logical_Operator_out2349_out1 <= Logical_Operator_out807_out1 XOR Logical_Operator_out815_out1;

  Logical_Operator_out2350_out1 <= Logical_Operator_out808_out1 XOR Logical_Operator_out816_out1;

  Logical_Operator_out2351_out1 <= Logical_Operator_out296_out1 XOR Logical_Operator_out304_out1;

  Logical_Operator_out2352_out1 <= in592 XOR in608;

  Logical_Operator_out2353_out1 <= Logical_Operator_out1841_out1 XOR Logical_Operator_out1849_out1;

  Logical_Operator_out2354_out1 <= Logical_Operator_out1842_out1 XOR Logical_Operator_out1850_out1;

  Logical_Operator_out2355_out1 <= Logical_Operator_out1843_out1 XOR Logical_Operator_out1851_out1;

  Logical_Operator_out2356_out1 <= Logical_Operator_out1844_out1 XOR Logical_Operator_out1852_out1;

  Logical_Operator_out2357_out1 <= Logical_Operator_out1845_out1 XOR Logical_Operator_out1853_out1;

  Logical_Operator_out2358_out1 <= Logical_Operator_out1846_out1 XOR Logical_Operator_out1854_out1;

  Logical_Operator_out2359_out1 <= Logical_Operator_out1847_out1 XOR Logical_Operator_out1855_out1;

  Logical_Operator_out2360_out1 <= Logical_Operator_out1848_out1 XOR Logical_Operator_out1856_out1;

  Logical_Operator_out2361_out1 <= Logical_Operator_out1333_out1 XOR Logical_Operator_out1341_out1;

  Logical_Operator_out2362_out1 <= Logical_Operator_out1334_out1 XOR Logical_Operator_out1342_out1;

  Logical_Operator_out2363_out1 <= Logical_Operator_out1335_out1 XOR Logical_Operator_out1343_out1;

  Logical_Operator_out2364_out1 <= Logical_Operator_out1336_out1 XOR Logical_Operator_out1344_out1;

  Logical_Operator_out2365_out1 <= Logical_Operator_out823_out1 XOR Logical_Operator_out831_out1;

  Logical_Operator_out2366_out1 <= Logical_Operator_out824_out1 XOR Logical_Operator_out832_out1;

  Logical_Operator_out2367_out1 <= Logical_Operator_out312_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out2368_out1 <= in624 XOR in640;

  Logical_Operator_out2369_out1 <= Logical_Operator_out1857_out1 XOR Logical_Operator_out1865_out1;

  Logical_Operator_out2370_out1 <= Logical_Operator_out1858_out1 XOR Logical_Operator_out1866_out1;

  Logical_Operator_out2371_out1 <= Logical_Operator_out1859_out1 XOR Logical_Operator_out1867_out1;

  Logical_Operator_out2372_out1 <= Logical_Operator_out1860_out1 XOR Logical_Operator_out1868_out1;

  Logical_Operator_out2373_out1 <= Logical_Operator_out1861_out1 XOR Logical_Operator_out1869_out1;

  Logical_Operator_out2374_out1 <= Logical_Operator_out1862_out1 XOR Logical_Operator_out1870_out1;

  Logical_Operator_out2375_out1 <= Logical_Operator_out1863_out1 XOR Logical_Operator_out1871_out1;

  Logical_Operator_out2376_out1 <= Logical_Operator_out1864_out1 XOR Logical_Operator_out1872_out1;

  Logical_Operator_out2377_out1 <= Logical_Operator_out1349_out1 XOR Logical_Operator_out1357_out1;

  Logical_Operator_out2378_out1 <= Logical_Operator_out1350_out1 XOR Logical_Operator_out1358_out1;

  Logical_Operator_out2379_out1 <= Logical_Operator_out1351_out1 XOR Logical_Operator_out1359_out1;

  Logical_Operator_out2380_out1 <= Logical_Operator_out1352_out1 XOR Logical_Operator_out1360_out1;

  Logical_Operator_out2381_out1 <= Logical_Operator_out839_out1 XOR Logical_Operator_out847_out1;

  Logical_Operator_out2382_out1 <= Logical_Operator_out840_out1 XOR Logical_Operator_out848_out1;

  Logical_Operator_out2383_out1 <= Logical_Operator_out328_out1 XOR Logical_Operator_out336_out1;

  Logical_Operator_out2384_out1 <= in656 XOR in672;

  Logical_Operator_out2385_out1 <= Logical_Operator_out1873_out1 XOR Logical_Operator_out1881_out1;

  Logical_Operator_out2386_out1 <= Logical_Operator_out1874_out1 XOR Logical_Operator_out1882_out1;

  Logical_Operator_out2387_out1 <= Logical_Operator_out1875_out1 XOR Logical_Operator_out1883_out1;

  Logical_Operator_out2388_out1 <= Logical_Operator_out1876_out1 XOR Logical_Operator_out1884_out1;

  Logical_Operator_out2389_out1 <= Logical_Operator_out1877_out1 XOR Logical_Operator_out1885_out1;

  Logical_Operator_out2390_out1 <= Logical_Operator_out1878_out1 XOR Logical_Operator_out1886_out1;

  Logical_Operator_out2391_out1 <= Logical_Operator_out1879_out1 XOR Logical_Operator_out1887_out1;

  Logical_Operator_out2392_out1 <= Logical_Operator_out1880_out1 XOR Logical_Operator_out1888_out1;

  Logical_Operator_out2393_out1 <= Logical_Operator_out1365_out1 XOR Logical_Operator_out1373_out1;

  Logical_Operator_out2394_out1 <= Logical_Operator_out1366_out1 XOR Logical_Operator_out1374_out1;

  Logical_Operator_out2395_out1 <= Logical_Operator_out1367_out1 XOR Logical_Operator_out1375_out1;

  Logical_Operator_out2396_out1 <= Logical_Operator_out1368_out1 XOR Logical_Operator_out1376_out1;

  Logical_Operator_out2397_out1 <= Logical_Operator_out855_out1 XOR Logical_Operator_out863_out1;

  Logical_Operator_out2398_out1 <= Logical_Operator_out856_out1 XOR Logical_Operator_out864_out1;

  Logical_Operator_out2399_out1 <= Logical_Operator_out344_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out2400_out1 <= in688 XOR in704;

  Logical_Operator_out2401_out1 <= Logical_Operator_out1889_out1 XOR Logical_Operator_out1897_out1;

  Logical_Operator_out2402_out1 <= Logical_Operator_out1890_out1 XOR Logical_Operator_out1898_out1;

  Logical_Operator_out2403_out1 <= Logical_Operator_out1891_out1 XOR Logical_Operator_out1899_out1;

  Logical_Operator_out2404_out1 <= Logical_Operator_out1892_out1 XOR Logical_Operator_out1900_out1;

  Logical_Operator_out2405_out1 <= Logical_Operator_out1893_out1 XOR Logical_Operator_out1901_out1;

  Logical_Operator_out2406_out1 <= Logical_Operator_out1894_out1 XOR Logical_Operator_out1902_out1;

  Logical_Operator_out2407_out1 <= Logical_Operator_out1895_out1 XOR Logical_Operator_out1903_out1;

  Logical_Operator_out2408_out1 <= Logical_Operator_out1896_out1 XOR Logical_Operator_out1904_out1;

  Logical_Operator_out2409_out1 <= Logical_Operator_out1381_out1 XOR Logical_Operator_out1389_out1;

  Logical_Operator_out2410_out1 <= Logical_Operator_out1382_out1 XOR Logical_Operator_out1390_out1;

  Logical_Operator_out2411_out1 <= Logical_Operator_out1383_out1 XOR Logical_Operator_out1391_out1;

  Logical_Operator_out2412_out1 <= Logical_Operator_out1384_out1 XOR Logical_Operator_out1392_out1;

  Logical_Operator_out2413_out1 <= Logical_Operator_out871_out1 XOR Logical_Operator_out879_out1;

  Logical_Operator_out2414_out1 <= Logical_Operator_out872_out1 XOR Logical_Operator_out880_out1;

  Logical_Operator_out2415_out1 <= Logical_Operator_out360_out1 XOR Logical_Operator_out368_out1;

  Logical_Operator_out2416_out1 <= in720 XOR in736;

  Logical_Operator_out2417_out1 <= Logical_Operator_out1905_out1 XOR Logical_Operator_out1913_out1;

  Logical_Operator_out2418_out1 <= Logical_Operator_out1906_out1 XOR Logical_Operator_out1914_out1;

  Logical_Operator_out2419_out1 <= Logical_Operator_out1907_out1 XOR Logical_Operator_out1915_out1;

  Logical_Operator_out2420_out1 <= Logical_Operator_out1908_out1 XOR Logical_Operator_out1916_out1;

  Logical_Operator_out2421_out1 <= Logical_Operator_out1909_out1 XOR Logical_Operator_out1917_out1;

  Logical_Operator_out2422_out1 <= Logical_Operator_out1910_out1 XOR Logical_Operator_out1918_out1;

  Logical_Operator_out2423_out1 <= Logical_Operator_out1911_out1 XOR Logical_Operator_out1919_out1;

  Logical_Operator_out2424_out1 <= Logical_Operator_out1912_out1 XOR Logical_Operator_out1920_out1;

  Logical_Operator_out2425_out1 <= Logical_Operator_out1397_out1 XOR Logical_Operator_out1405_out1;

  Logical_Operator_out2426_out1 <= Logical_Operator_out1398_out1 XOR Logical_Operator_out1406_out1;

  Logical_Operator_out2427_out1 <= Logical_Operator_out1399_out1 XOR Logical_Operator_out1407_out1;

  Logical_Operator_out2428_out1 <= Logical_Operator_out1400_out1 XOR Logical_Operator_out1408_out1;

  Logical_Operator_out2429_out1 <= Logical_Operator_out887_out1 XOR Logical_Operator_out895_out1;

  Logical_Operator_out2430_out1 <= Logical_Operator_out888_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out2431_out1 <= Logical_Operator_out376_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out2432_out1 <= in752 XOR in768;

  Logical_Operator_out2433_out1 <= Logical_Operator_out1921_out1 XOR Logical_Operator_out1929_out1;

  Logical_Operator_out2434_out1 <= Logical_Operator_out1922_out1 XOR Logical_Operator_out1930_out1;

  Logical_Operator_out2435_out1 <= Logical_Operator_out1923_out1 XOR Logical_Operator_out1931_out1;

  Logical_Operator_out2436_out1 <= Logical_Operator_out1924_out1 XOR Logical_Operator_out1932_out1;

  Logical_Operator_out2437_out1 <= Logical_Operator_out1925_out1 XOR Logical_Operator_out1933_out1;

  Logical_Operator_out2438_out1 <= Logical_Operator_out1926_out1 XOR Logical_Operator_out1934_out1;

  Logical_Operator_out2439_out1 <= Logical_Operator_out1927_out1 XOR Logical_Operator_out1935_out1;

  Logical_Operator_out2440_out1 <= Logical_Operator_out1928_out1 XOR Logical_Operator_out1936_out1;

  Logical_Operator_out2441_out1 <= Logical_Operator_out1413_out1 XOR Logical_Operator_out1421_out1;

  Logical_Operator_out2442_out1 <= Logical_Operator_out1414_out1 XOR Logical_Operator_out1422_out1;

  Logical_Operator_out2443_out1 <= Logical_Operator_out1415_out1 XOR Logical_Operator_out1423_out1;

  Logical_Operator_out2444_out1 <= Logical_Operator_out1416_out1 XOR Logical_Operator_out1424_out1;

  Logical_Operator_out2445_out1 <= Logical_Operator_out903_out1 XOR Logical_Operator_out911_out1;

  Logical_Operator_out2446_out1 <= Logical_Operator_out904_out1 XOR Logical_Operator_out912_out1;

  Logical_Operator_out2447_out1 <= Logical_Operator_out392_out1 XOR Logical_Operator_out400_out1;

  Logical_Operator_out2448_out1 <= in784 XOR in800;

  Logical_Operator_out2449_out1 <= Logical_Operator_out1937_out1 XOR Logical_Operator_out1945_out1;

  Logical_Operator_out2450_out1 <= Logical_Operator_out1938_out1 XOR Logical_Operator_out1946_out1;

  Logical_Operator_out2451_out1 <= Logical_Operator_out1939_out1 XOR Logical_Operator_out1947_out1;

  Logical_Operator_out2452_out1 <= Logical_Operator_out1940_out1 XOR Logical_Operator_out1948_out1;

  Logical_Operator_out2453_out1 <= Logical_Operator_out1941_out1 XOR Logical_Operator_out1949_out1;

  Logical_Operator_out2454_out1 <= Logical_Operator_out1942_out1 XOR Logical_Operator_out1950_out1;

  Logical_Operator_out2455_out1 <= Logical_Operator_out1943_out1 XOR Logical_Operator_out1951_out1;

  Logical_Operator_out2456_out1 <= Logical_Operator_out1944_out1 XOR Logical_Operator_out1952_out1;

  Logical_Operator_out2457_out1 <= Logical_Operator_out1429_out1 XOR Logical_Operator_out1437_out1;

  Logical_Operator_out2458_out1 <= Logical_Operator_out1430_out1 XOR Logical_Operator_out1438_out1;

  Logical_Operator_out2459_out1 <= Logical_Operator_out1431_out1 XOR Logical_Operator_out1439_out1;

  Logical_Operator_out2460_out1 <= Logical_Operator_out1432_out1 XOR Logical_Operator_out1440_out1;

  Logical_Operator_out2461_out1 <= Logical_Operator_out919_out1 XOR Logical_Operator_out927_out1;

  Logical_Operator_out2462_out1 <= Logical_Operator_out920_out1 XOR Logical_Operator_out928_out1;

  Logical_Operator_out2463_out1 <= Logical_Operator_out408_out1 XOR Logical_Operator_out416_out1;

  Logical_Operator_out2464_out1 <= in816 XOR in832;

  Logical_Operator_out2465_out1 <= Logical_Operator_out1953_out1 XOR Logical_Operator_out1961_out1;

  Logical_Operator_out2466_out1 <= Logical_Operator_out1954_out1 XOR Logical_Operator_out1962_out1;

  Logical_Operator_out2467_out1 <= Logical_Operator_out1955_out1 XOR Logical_Operator_out1963_out1;

  Logical_Operator_out2468_out1 <= Logical_Operator_out1956_out1 XOR Logical_Operator_out1964_out1;

  Logical_Operator_out2469_out1 <= Logical_Operator_out1957_out1 XOR Logical_Operator_out1965_out1;

  Logical_Operator_out2470_out1 <= Logical_Operator_out1958_out1 XOR Logical_Operator_out1966_out1;

  Logical_Operator_out2471_out1 <= Logical_Operator_out1959_out1 XOR Logical_Operator_out1967_out1;

  Logical_Operator_out2472_out1 <= Logical_Operator_out1960_out1 XOR Logical_Operator_out1968_out1;

  Logical_Operator_out2473_out1 <= Logical_Operator_out1445_out1 XOR Logical_Operator_out1453_out1;

  Logical_Operator_out2474_out1 <= Logical_Operator_out1446_out1 XOR Logical_Operator_out1454_out1;

  Logical_Operator_out2475_out1 <= Logical_Operator_out1447_out1 XOR Logical_Operator_out1455_out1;

  Logical_Operator_out2476_out1 <= Logical_Operator_out1448_out1 XOR Logical_Operator_out1456_out1;

  Logical_Operator_out2477_out1 <= Logical_Operator_out935_out1 XOR Logical_Operator_out943_out1;

  Logical_Operator_out2478_out1 <= Logical_Operator_out936_out1 XOR Logical_Operator_out944_out1;

  Logical_Operator_out2479_out1 <= Logical_Operator_out424_out1 XOR Logical_Operator_out432_out1;

  Logical_Operator_out2480_out1 <= in848 XOR in864;

  Logical_Operator_out2481_out1 <= Logical_Operator_out1969_out1 XOR Logical_Operator_out1977_out1;

  Logical_Operator_out2482_out1 <= Logical_Operator_out1970_out1 XOR Logical_Operator_out1978_out1;

  Logical_Operator_out2483_out1 <= Logical_Operator_out1971_out1 XOR Logical_Operator_out1979_out1;

  Logical_Operator_out2484_out1 <= Logical_Operator_out1972_out1 XOR Logical_Operator_out1980_out1;

  Logical_Operator_out2485_out1 <= Logical_Operator_out1973_out1 XOR Logical_Operator_out1981_out1;

  Logical_Operator_out2486_out1 <= Logical_Operator_out1974_out1 XOR Logical_Operator_out1982_out1;

  Logical_Operator_out2487_out1 <= Logical_Operator_out1975_out1 XOR Logical_Operator_out1983_out1;

  Logical_Operator_out2488_out1 <= Logical_Operator_out1976_out1 XOR Logical_Operator_out1984_out1;

  Logical_Operator_out2489_out1 <= Logical_Operator_out1461_out1 XOR Logical_Operator_out1469_out1;

  Logical_Operator_out2490_out1 <= Logical_Operator_out1462_out1 XOR Logical_Operator_out1470_out1;

  Logical_Operator_out2491_out1 <= Logical_Operator_out1463_out1 XOR Logical_Operator_out1471_out1;

  Logical_Operator_out2492_out1 <= Logical_Operator_out1464_out1 XOR Logical_Operator_out1472_out1;

  Logical_Operator_out2493_out1 <= Logical_Operator_out951_out1 XOR Logical_Operator_out959_out1;

  Logical_Operator_out2494_out1 <= Logical_Operator_out952_out1 XOR Logical_Operator_out960_out1;

  Logical_Operator_out2495_out1 <= Logical_Operator_out440_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out2496_out1 <= in880 XOR in896;

  Logical_Operator_out2497_out1 <= Logical_Operator_out1985_out1 XOR Logical_Operator_out1993_out1;

  Logical_Operator_out2498_out1 <= Logical_Operator_out1986_out1 XOR Logical_Operator_out1994_out1;

  Logical_Operator_out2499_out1 <= Logical_Operator_out1987_out1 XOR Logical_Operator_out1995_out1;

  Logical_Operator_out2500_out1 <= Logical_Operator_out1988_out1 XOR Logical_Operator_out1996_out1;

  Logical_Operator_out2501_out1 <= Logical_Operator_out1989_out1 XOR Logical_Operator_out1997_out1;

  Logical_Operator_out2502_out1 <= Logical_Operator_out1990_out1 XOR Logical_Operator_out1998_out1;

  Logical_Operator_out2503_out1 <= Logical_Operator_out1991_out1 XOR Logical_Operator_out1999_out1;

  Logical_Operator_out2504_out1 <= Logical_Operator_out1992_out1 XOR Logical_Operator_out2000_out1;

  Logical_Operator_out2505_out1 <= Logical_Operator_out1477_out1 XOR Logical_Operator_out1485_out1;

  Logical_Operator_out2506_out1 <= Logical_Operator_out1478_out1 XOR Logical_Operator_out1486_out1;

  Logical_Operator_out2507_out1 <= Logical_Operator_out1479_out1 XOR Logical_Operator_out1487_out1;

  Logical_Operator_out2508_out1 <= Logical_Operator_out1480_out1 XOR Logical_Operator_out1488_out1;

  Logical_Operator_out2509_out1 <= Logical_Operator_out967_out1 XOR Logical_Operator_out975_out1;

  Logical_Operator_out2510_out1 <= Logical_Operator_out968_out1 XOR Logical_Operator_out976_out1;

  Logical_Operator_out2511_out1 <= Logical_Operator_out456_out1 XOR Logical_Operator_out464_out1;

  Logical_Operator_out2512_out1 <= in912 XOR in928;

  Logical_Operator_out2513_out1 <= Logical_Operator_out2001_out1 XOR Logical_Operator_out2009_out1;

  Logical_Operator_out2514_out1 <= Logical_Operator_out2002_out1 XOR Logical_Operator_out2010_out1;

  Logical_Operator_out2515_out1 <= Logical_Operator_out2003_out1 XOR Logical_Operator_out2011_out1;

  Logical_Operator_out2516_out1 <= Logical_Operator_out2004_out1 XOR Logical_Operator_out2012_out1;

  Logical_Operator_out2517_out1 <= Logical_Operator_out2005_out1 XOR Logical_Operator_out2013_out1;

  Logical_Operator_out2518_out1 <= Logical_Operator_out2006_out1 XOR Logical_Operator_out2014_out1;

  Logical_Operator_out2519_out1 <= Logical_Operator_out2007_out1 XOR Logical_Operator_out2015_out1;

  Logical_Operator_out2520_out1 <= Logical_Operator_out2008_out1 XOR Logical_Operator_out2016_out1;

  Logical_Operator_out2521_out1 <= Logical_Operator_out1493_out1 XOR Logical_Operator_out1501_out1;

  Logical_Operator_out2522_out1 <= Logical_Operator_out1494_out1 XOR Logical_Operator_out1502_out1;

  Logical_Operator_out2523_out1 <= Logical_Operator_out1495_out1 XOR Logical_Operator_out1503_out1;

  Logical_Operator_out2524_out1 <= Logical_Operator_out1496_out1 XOR Logical_Operator_out1504_out1;

  Logical_Operator_out2525_out1 <= Logical_Operator_out983_out1 XOR Logical_Operator_out991_out1;

  Logical_Operator_out2526_out1 <= Logical_Operator_out984_out1 XOR Logical_Operator_out992_out1;

  Logical_Operator_out2527_out1 <= Logical_Operator_out472_out1 XOR Logical_Operator_out480_out1;

  Logical_Operator_out2528_out1 <= in944 XOR in960;

  Logical_Operator_out2529_out1 <= Logical_Operator_out2017_out1 XOR Logical_Operator_out2025_out1;

  Logical_Operator_out2530_out1 <= Logical_Operator_out2018_out1 XOR Logical_Operator_out2026_out1;

  Logical_Operator_out2531_out1 <= Logical_Operator_out2019_out1 XOR Logical_Operator_out2027_out1;

  Logical_Operator_out2532_out1 <= Logical_Operator_out2020_out1 XOR Logical_Operator_out2028_out1;

  Logical_Operator_out2533_out1 <= Logical_Operator_out2021_out1 XOR Logical_Operator_out2029_out1;

  Logical_Operator_out2534_out1 <= Logical_Operator_out2022_out1 XOR Logical_Operator_out2030_out1;

  Logical_Operator_out2535_out1 <= Logical_Operator_out2023_out1 XOR Logical_Operator_out2031_out1;

  Logical_Operator_out2536_out1 <= Logical_Operator_out2024_out1 XOR Logical_Operator_out2032_out1;

  Logical_Operator_out2537_out1 <= Logical_Operator_out1509_out1 XOR Logical_Operator_out1517_out1;

  Logical_Operator_out2538_out1 <= Logical_Operator_out1510_out1 XOR Logical_Operator_out1518_out1;

  Logical_Operator_out2539_out1 <= Logical_Operator_out1511_out1 XOR Logical_Operator_out1519_out1;

  Logical_Operator_out2540_out1 <= Logical_Operator_out1512_out1 XOR Logical_Operator_out1520_out1;

  Logical_Operator_out2541_out1 <= Logical_Operator_out999_out1 XOR Logical_Operator_out1007_out1;

  Logical_Operator_out2542_out1 <= Logical_Operator_out1000_out1 XOR Logical_Operator_out1008_out1;

  Logical_Operator_out2543_out1 <= Logical_Operator_out488_out1 XOR Logical_Operator_out496_out1;

  Logical_Operator_out2544_out1 <= in976 XOR in992;

  Logical_Operator_out2545_out1 <= Logical_Operator_out2033_out1 XOR Logical_Operator_out2041_out1;

  Logical_Operator_out2546_out1 <= Logical_Operator_out2034_out1 XOR Logical_Operator_out2042_out1;

  Logical_Operator_out2547_out1 <= Logical_Operator_out2035_out1 XOR Logical_Operator_out2043_out1;

  Logical_Operator_out2548_out1 <= Logical_Operator_out2036_out1 XOR Logical_Operator_out2044_out1;

  Logical_Operator_out2549_out1 <= Logical_Operator_out2037_out1 XOR Logical_Operator_out2045_out1;

  Logical_Operator_out2550_out1 <= Logical_Operator_out2038_out1 XOR Logical_Operator_out2046_out1;

  Logical_Operator_out2551_out1 <= Logical_Operator_out2039_out1 XOR Logical_Operator_out2047_out1;

  Logical_Operator_out2552_out1 <= Logical_Operator_out2040_out1 XOR Logical_Operator_out2048_out1;

  Logical_Operator_out2553_out1 <= Logical_Operator_out1525_out1 XOR Logical_Operator_out1533_out1;

  Logical_Operator_out2554_out1 <= Logical_Operator_out1526_out1 XOR Logical_Operator_out1534_out1;

  Logical_Operator_out2555_out1 <= Logical_Operator_out1527_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out2556_out1 <= Logical_Operator_out1528_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out2557_out1 <= Logical_Operator_out1015_out1 XOR Logical_Operator_out1023_out1;

  Logical_Operator_out2558_out1 <= Logical_Operator_out1016_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out2559_out1 <= Logical_Operator_out504_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out2560_out1 <= in1008 XOR in1024;

  Logical_Operator_out2561_out1 <= Logical_Operator_out2049_out1 XOR Logical_Operator_out2065_out1;

  Logical_Operator_out2562_out1 <= Logical_Operator_out2050_out1 XOR Logical_Operator_out2066_out1;

  Logical_Operator_out2563_out1 <= Logical_Operator_out2051_out1 XOR Logical_Operator_out2067_out1;

  Logical_Operator_out2564_out1 <= Logical_Operator_out2052_out1 XOR Logical_Operator_out2068_out1;

  Logical_Operator_out2565_out1 <= Logical_Operator_out2053_out1 XOR Logical_Operator_out2069_out1;

  Logical_Operator_out2566_out1 <= Logical_Operator_out2054_out1 XOR Logical_Operator_out2070_out1;

  Logical_Operator_out2567_out1 <= Logical_Operator_out2055_out1 XOR Logical_Operator_out2071_out1;

  Logical_Operator_out2568_out1 <= Logical_Operator_out2056_out1 XOR Logical_Operator_out2072_out1;

  Logical_Operator_out2569_out1 <= Logical_Operator_out2057_out1 XOR Logical_Operator_out2073_out1;

  Logical_Operator_out2570_out1 <= Logical_Operator_out2058_out1 XOR Logical_Operator_out2074_out1;

  Logical_Operator_out2571_out1 <= Logical_Operator_out2059_out1 XOR Logical_Operator_out2075_out1;

  Logical_Operator_out2572_out1 <= Logical_Operator_out2060_out1 XOR Logical_Operator_out2076_out1;

  Logical_Operator_out2573_out1 <= Logical_Operator_out2061_out1 XOR Logical_Operator_out2077_out1;

  Logical_Operator_out2574_out1 <= Logical_Operator_out2062_out1 XOR Logical_Operator_out2078_out1;

  Logical_Operator_out2575_out1 <= Logical_Operator_out2063_out1 XOR Logical_Operator_out2079_out1;

  Logical_Operator_out2576_out1 <= Logical_Operator_out2064_out1 XOR Logical_Operator_out2080_out1;

  Logical_Operator_out2577_out1 <= Logical_Operator_out1545_out1 XOR Logical_Operator_out1561_out1;

  Logical_Operator_out2578_out1 <= Logical_Operator_out1546_out1 XOR Logical_Operator_out1562_out1;

  Logical_Operator_out2579_out1 <= Logical_Operator_out1547_out1 XOR Logical_Operator_out1563_out1;

  Logical_Operator_out2580_out1 <= Logical_Operator_out1548_out1 XOR Logical_Operator_out1564_out1;

  Logical_Operator_out2581_out1 <= Logical_Operator_out1549_out1 XOR Logical_Operator_out1565_out1;

  Logical_Operator_out2582_out1 <= Logical_Operator_out1550_out1 XOR Logical_Operator_out1566_out1;

  Logical_Operator_out2583_out1 <= Logical_Operator_out1551_out1 XOR Logical_Operator_out1567_out1;

  Logical_Operator_out2584_out1 <= Logical_Operator_out1552_out1 XOR Logical_Operator_out1568_out1;

  Logical_Operator_out2585_out1 <= Logical_Operator_out1037_out1 XOR Logical_Operator_out1053_out1;

  Logical_Operator_out2586_out1 <= Logical_Operator_out1038_out1 XOR Logical_Operator_out1054_out1;

  Logical_Operator_out2587_out1 <= Logical_Operator_out1039_out1 XOR Logical_Operator_out1055_out1;

  Logical_Operator_out2588_out1 <= Logical_Operator_out1040_out1 XOR Logical_Operator_out1056_out1;

  Logical_Operator_out2589_out1 <= Logical_Operator_out527_out1 XOR Logical_Operator_out543_out1;

  Logical_Operator_out2590_out1 <= Logical_Operator_out528_out1 XOR Logical_Operator_out544_out1;

  Logical_Operator_out2591_out1 <= Logical_Operator_out16_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out2592_out1 <= in32 XOR in64;

  Logical_Operator_out2593_out1 <= Logical_Operator_out2081_out1 XOR Logical_Operator_out2097_out1;

  Logical_Operator_out2594_out1 <= Logical_Operator_out2082_out1 XOR Logical_Operator_out2098_out1;

  Logical_Operator_out2595_out1 <= Logical_Operator_out2083_out1 XOR Logical_Operator_out2099_out1;

  Logical_Operator_out2596_out1 <= Logical_Operator_out2084_out1 XOR Logical_Operator_out2100_out1;

  Logical_Operator_out2597_out1 <= Logical_Operator_out2085_out1 XOR Logical_Operator_out2101_out1;

  Logical_Operator_out2598_out1 <= Logical_Operator_out2086_out1 XOR Logical_Operator_out2102_out1;

  Logical_Operator_out2599_out1 <= Logical_Operator_out2087_out1 XOR Logical_Operator_out2103_out1;

  Logical_Operator_out2600_out1 <= Logical_Operator_out2088_out1 XOR Logical_Operator_out2104_out1;

  Logical_Operator_out2601_out1 <= Logical_Operator_out2089_out1 XOR Logical_Operator_out2105_out1;

  Logical_Operator_out2602_out1 <= Logical_Operator_out2090_out1 XOR Logical_Operator_out2106_out1;

  Logical_Operator_out2603_out1 <= Logical_Operator_out2091_out1 XOR Logical_Operator_out2107_out1;

  Logical_Operator_out2604_out1 <= Logical_Operator_out2092_out1 XOR Logical_Operator_out2108_out1;

  Logical_Operator_out2605_out1 <= Logical_Operator_out2093_out1 XOR Logical_Operator_out2109_out1;

  Logical_Operator_out2606_out1 <= Logical_Operator_out2094_out1 XOR Logical_Operator_out2110_out1;

  Logical_Operator_out2607_out1 <= Logical_Operator_out2095_out1 XOR Logical_Operator_out2111_out1;

  Logical_Operator_out2608_out1 <= Logical_Operator_out2096_out1 XOR Logical_Operator_out2112_out1;

  Logical_Operator_out2609_out1 <= Logical_Operator_out1577_out1 XOR Logical_Operator_out1593_out1;

  Logical_Operator_out2610_out1 <= Logical_Operator_out1578_out1 XOR Logical_Operator_out1594_out1;

  Logical_Operator_out2611_out1 <= Logical_Operator_out1579_out1 XOR Logical_Operator_out1595_out1;

  Logical_Operator_out2612_out1 <= Logical_Operator_out1580_out1 XOR Logical_Operator_out1596_out1;

  Logical_Operator_out2613_out1 <= Logical_Operator_out1581_out1 XOR Logical_Operator_out1597_out1;

  Logical_Operator_out2614_out1 <= Logical_Operator_out1582_out1 XOR Logical_Operator_out1598_out1;

  Logical_Operator_out2615_out1 <= Logical_Operator_out1583_out1 XOR Logical_Operator_out1599_out1;

  Logical_Operator_out2616_out1 <= Logical_Operator_out1584_out1 XOR Logical_Operator_out1600_out1;

  Logical_Operator_out2617_out1 <= Logical_Operator_out1069_out1 XOR Logical_Operator_out1085_out1;

  Logical_Operator_out2618_out1 <= Logical_Operator_out1070_out1 XOR Logical_Operator_out1086_out1;

  Logical_Operator_out2619_out1 <= Logical_Operator_out1071_out1 XOR Logical_Operator_out1087_out1;

  Logical_Operator_out2620_out1 <= Logical_Operator_out1072_out1 XOR Logical_Operator_out1088_out1;

  Logical_Operator_out2621_out1 <= Logical_Operator_out559_out1 XOR Logical_Operator_out575_out1;

  Logical_Operator_out2622_out1 <= Logical_Operator_out560_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out2623_out1 <= Logical_Operator_out48_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out2624_out1 <= in96 XOR in128;

  Logical_Operator_out2625_out1 <= Logical_Operator_out2113_out1 XOR Logical_Operator_out2129_out1;

  Logical_Operator_out2626_out1 <= Logical_Operator_out2114_out1 XOR Logical_Operator_out2130_out1;

  Logical_Operator_out2627_out1 <= Logical_Operator_out2115_out1 XOR Logical_Operator_out2131_out1;

  Logical_Operator_out2628_out1 <= Logical_Operator_out2116_out1 XOR Logical_Operator_out2132_out1;

  Logical_Operator_out2629_out1 <= Logical_Operator_out2117_out1 XOR Logical_Operator_out2133_out1;

  Logical_Operator_out2630_out1 <= Logical_Operator_out2118_out1 XOR Logical_Operator_out2134_out1;

  Logical_Operator_out2631_out1 <= Logical_Operator_out2119_out1 XOR Logical_Operator_out2135_out1;

  Logical_Operator_out2632_out1 <= Logical_Operator_out2120_out1 XOR Logical_Operator_out2136_out1;

  Logical_Operator_out2633_out1 <= Logical_Operator_out2121_out1 XOR Logical_Operator_out2137_out1;

  Logical_Operator_out2634_out1 <= Logical_Operator_out2122_out1 XOR Logical_Operator_out2138_out1;

  Logical_Operator_out2635_out1 <= Logical_Operator_out2123_out1 XOR Logical_Operator_out2139_out1;

  Logical_Operator_out2636_out1 <= Logical_Operator_out2124_out1 XOR Logical_Operator_out2140_out1;

  Logical_Operator_out2637_out1 <= Logical_Operator_out2125_out1 XOR Logical_Operator_out2141_out1;

  Logical_Operator_out2638_out1 <= Logical_Operator_out2126_out1 XOR Logical_Operator_out2142_out1;

  Logical_Operator_out2639_out1 <= Logical_Operator_out2127_out1 XOR Logical_Operator_out2143_out1;

  Logical_Operator_out2640_out1 <= Logical_Operator_out2128_out1 XOR Logical_Operator_out2144_out1;

  Logical_Operator_out2641_out1 <= Logical_Operator_out1609_out1 XOR Logical_Operator_out1625_out1;

  Logical_Operator_out2642_out1 <= Logical_Operator_out1610_out1 XOR Logical_Operator_out1626_out1;

  Logical_Operator_out2643_out1 <= Logical_Operator_out1611_out1 XOR Logical_Operator_out1627_out1;

  Logical_Operator_out2644_out1 <= Logical_Operator_out1612_out1 XOR Logical_Operator_out1628_out1;

  Logical_Operator_out2645_out1 <= Logical_Operator_out1613_out1 XOR Logical_Operator_out1629_out1;

  Logical_Operator_out2646_out1 <= Logical_Operator_out1614_out1 XOR Logical_Operator_out1630_out1;

  Logical_Operator_out2647_out1 <= Logical_Operator_out1615_out1 XOR Logical_Operator_out1631_out1;

  Logical_Operator_out2648_out1 <= Logical_Operator_out1616_out1 XOR Logical_Operator_out1632_out1;

  Logical_Operator_out2649_out1 <= Logical_Operator_out1101_out1 XOR Logical_Operator_out1117_out1;

  Logical_Operator_out2650_out1 <= Logical_Operator_out1102_out1 XOR Logical_Operator_out1118_out1;

  Logical_Operator_out2651_out1 <= Logical_Operator_out1103_out1 XOR Logical_Operator_out1119_out1;

  Logical_Operator_out2652_out1 <= Logical_Operator_out1104_out1 XOR Logical_Operator_out1120_out1;

  Logical_Operator_out2653_out1 <= Logical_Operator_out591_out1 XOR Logical_Operator_out607_out1;

  Logical_Operator_out2654_out1 <= Logical_Operator_out592_out1 XOR Logical_Operator_out608_out1;

  Logical_Operator_out2655_out1 <= Logical_Operator_out80_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out2656_out1 <= in160 XOR in192;

  Logical_Operator_out2657_out1 <= Logical_Operator_out2145_out1 XOR Logical_Operator_out2161_out1;

  Logical_Operator_out2658_out1 <= Logical_Operator_out2146_out1 XOR Logical_Operator_out2162_out1;

  Logical_Operator_out2659_out1 <= Logical_Operator_out2147_out1 XOR Logical_Operator_out2163_out1;

  Logical_Operator_out2660_out1 <= Logical_Operator_out2148_out1 XOR Logical_Operator_out2164_out1;

  Logical_Operator_out2661_out1 <= Logical_Operator_out2149_out1 XOR Logical_Operator_out2165_out1;

  Logical_Operator_out2662_out1 <= Logical_Operator_out2150_out1 XOR Logical_Operator_out2166_out1;

  Logical_Operator_out2663_out1 <= Logical_Operator_out2151_out1 XOR Logical_Operator_out2167_out1;

  Logical_Operator_out2664_out1 <= Logical_Operator_out2152_out1 XOR Logical_Operator_out2168_out1;

  Logical_Operator_out2665_out1 <= Logical_Operator_out2153_out1 XOR Logical_Operator_out2169_out1;

  Logical_Operator_out2666_out1 <= Logical_Operator_out2154_out1 XOR Logical_Operator_out2170_out1;

  Logical_Operator_out2667_out1 <= Logical_Operator_out2155_out1 XOR Logical_Operator_out2171_out1;

  Logical_Operator_out2668_out1 <= Logical_Operator_out2156_out1 XOR Logical_Operator_out2172_out1;

  Logical_Operator_out2669_out1 <= Logical_Operator_out2157_out1 XOR Logical_Operator_out2173_out1;

  Logical_Operator_out2670_out1 <= Logical_Operator_out2158_out1 XOR Logical_Operator_out2174_out1;

  Logical_Operator_out2671_out1 <= Logical_Operator_out2159_out1 XOR Logical_Operator_out2175_out1;

  Logical_Operator_out2672_out1 <= Logical_Operator_out2160_out1 XOR Logical_Operator_out2176_out1;

  Logical_Operator_out2673_out1 <= Logical_Operator_out1641_out1 XOR Logical_Operator_out1657_out1;

  Logical_Operator_out2674_out1 <= Logical_Operator_out1642_out1 XOR Logical_Operator_out1658_out1;

  Logical_Operator_out2675_out1 <= Logical_Operator_out1643_out1 XOR Logical_Operator_out1659_out1;

  Logical_Operator_out2676_out1 <= Logical_Operator_out1644_out1 XOR Logical_Operator_out1660_out1;

  Logical_Operator_out2677_out1 <= Logical_Operator_out1645_out1 XOR Logical_Operator_out1661_out1;

  Logical_Operator_out2678_out1 <= Logical_Operator_out1646_out1 XOR Logical_Operator_out1662_out1;

  Logical_Operator_out2679_out1 <= Logical_Operator_out1647_out1 XOR Logical_Operator_out1663_out1;

  Logical_Operator_out2680_out1 <= Logical_Operator_out1648_out1 XOR Logical_Operator_out1664_out1;

  Logical_Operator_out2681_out1 <= Logical_Operator_out1133_out1 XOR Logical_Operator_out1149_out1;

  Logical_Operator_out2682_out1 <= Logical_Operator_out1134_out1 XOR Logical_Operator_out1150_out1;

  Logical_Operator_out2683_out1 <= Logical_Operator_out1135_out1 XOR Logical_Operator_out1151_out1;

  Logical_Operator_out2684_out1 <= Logical_Operator_out1136_out1 XOR Logical_Operator_out1152_out1;

  Logical_Operator_out2685_out1 <= Logical_Operator_out623_out1 XOR Logical_Operator_out639_out1;

  Logical_Operator_out2686_out1 <= Logical_Operator_out624_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out2687_out1 <= Logical_Operator_out112_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out2688_out1 <= in224 XOR in256;

  Logical_Operator_out2689_out1 <= Logical_Operator_out2177_out1 XOR Logical_Operator_out2193_out1;

  Logical_Operator_out2690_out1 <= Logical_Operator_out2178_out1 XOR Logical_Operator_out2194_out1;

  Logical_Operator_out2691_out1 <= Logical_Operator_out2179_out1 XOR Logical_Operator_out2195_out1;

  Logical_Operator_out2692_out1 <= Logical_Operator_out2180_out1 XOR Logical_Operator_out2196_out1;

  Logical_Operator_out2693_out1 <= Logical_Operator_out2181_out1 XOR Logical_Operator_out2197_out1;

  Logical_Operator_out2694_out1 <= Logical_Operator_out2182_out1 XOR Logical_Operator_out2198_out1;

  Logical_Operator_out2695_out1 <= Logical_Operator_out2183_out1 XOR Logical_Operator_out2199_out1;

  Logical_Operator_out2696_out1 <= Logical_Operator_out2184_out1 XOR Logical_Operator_out2200_out1;

  Logical_Operator_out2697_out1 <= Logical_Operator_out2185_out1 XOR Logical_Operator_out2201_out1;

  Logical_Operator_out2698_out1 <= Logical_Operator_out2186_out1 XOR Logical_Operator_out2202_out1;

  Logical_Operator_out2699_out1 <= Logical_Operator_out2187_out1 XOR Logical_Operator_out2203_out1;

  Logical_Operator_out2700_out1 <= Logical_Operator_out2188_out1 XOR Logical_Operator_out2204_out1;

  Logical_Operator_out2701_out1 <= Logical_Operator_out2189_out1 XOR Logical_Operator_out2205_out1;

  Logical_Operator_out2702_out1 <= Logical_Operator_out2190_out1 XOR Logical_Operator_out2206_out1;

  Logical_Operator_out2703_out1 <= Logical_Operator_out2191_out1 XOR Logical_Operator_out2207_out1;

  Logical_Operator_out2704_out1 <= Logical_Operator_out2192_out1 XOR Logical_Operator_out2208_out1;

  Logical_Operator_out2705_out1 <= Logical_Operator_out1673_out1 XOR Logical_Operator_out1689_out1;

  Logical_Operator_out2706_out1 <= Logical_Operator_out1674_out1 XOR Logical_Operator_out1690_out1;

  Logical_Operator_out2707_out1 <= Logical_Operator_out1675_out1 XOR Logical_Operator_out1691_out1;

  Logical_Operator_out2708_out1 <= Logical_Operator_out1676_out1 XOR Logical_Operator_out1692_out1;

  Logical_Operator_out2709_out1 <= Logical_Operator_out1677_out1 XOR Logical_Operator_out1693_out1;

  Logical_Operator_out2710_out1 <= Logical_Operator_out1678_out1 XOR Logical_Operator_out1694_out1;

  Logical_Operator_out2711_out1 <= Logical_Operator_out1679_out1 XOR Logical_Operator_out1695_out1;

  Logical_Operator_out2712_out1 <= Logical_Operator_out1680_out1 XOR Logical_Operator_out1696_out1;

  Logical_Operator_out2713_out1 <= Logical_Operator_out1165_out1 XOR Logical_Operator_out1181_out1;

  Logical_Operator_out2714_out1 <= Logical_Operator_out1166_out1 XOR Logical_Operator_out1182_out1;

  Logical_Operator_out2715_out1 <= Logical_Operator_out1167_out1 XOR Logical_Operator_out1183_out1;

  Logical_Operator_out2716_out1 <= Logical_Operator_out1168_out1 XOR Logical_Operator_out1184_out1;

  Logical_Operator_out2717_out1 <= Logical_Operator_out655_out1 XOR Logical_Operator_out671_out1;

  Logical_Operator_out2718_out1 <= Logical_Operator_out656_out1 XOR Logical_Operator_out672_out1;

  Logical_Operator_out2719_out1 <= Logical_Operator_out144_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out2720_out1 <= in288 XOR in320;

  Logical_Operator_out2721_out1 <= Logical_Operator_out2209_out1 XOR Logical_Operator_out2225_out1;

  Logical_Operator_out2722_out1 <= Logical_Operator_out2210_out1 XOR Logical_Operator_out2226_out1;

  Logical_Operator_out2723_out1 <= Logical_Operator_out2211_out1 XOR Logical_Operator_out2227_out1;

  Logical_Operator_out2724_out1 <= Logical_Operator_out2212_out1 XOR Logical_Operator_out2228_out1;

  Logical_Operator_out2725_out1 <= Logical_Operator_out2213_out1 XOR Logical_Operator_out2229_out1;

  Logical_Operator_out2726_out1 <= Logical_Operator_out2214_out1 XOR Logical_Operator_out2230_out1;

  Logical_Operator_out2727_out1 <= Logical_Operator_out2215_out1 XOR Logical_Operator_out2231_out1;

  Logical_Operator_out2728_out1 <= Logical_Operator_out2216_out1 XOR Logical_Operator_out2232_out1;

  Logical_Operator_out2729_out1 <= Logical_Operator_out2217_out1 XOR Logical_Operator_out2233_out1;

  Logical_Operator_out2730_out1 <= Logical_Operator_out2218_out1 XOR Logical_Operator_out2234_out1;

  Logical_Operator_out2731_out1 <= Logical_Operator_out2219_out1 XOR Logical_Operator_out2235_out1;

  Logical_Operator_out2732_out1 <= Logical_Operator_out2220_out1 XOR Logical_Operator_out2236_out1;

  Logical_Operator_out2733_out1 <= Logical_Operator_out2221_out1 XOR Logical_Operator_out2237_out1;

  Logical_Operator_out2734_out1 <= Logical_Operator_out2222_out1 XOR Logical_Operator_out2238_out1;

  Logical_Operator_out2735_out1 <= Logical_Operator_out2223_out1 XOR Logical_Operator_out2239_out1;

  Logical_Operator_out2736_out1 <= Logical_Operator_out2224_out1 XOR Logical_Operator_out2240_out1;

  Logical_Operator_out2737_out1 <= Logical_Operator_out1705_out1 XOR Logical_Operator_out1721_out1;

  Logical_Operator_out2738_out1 <= Logical_Operator_out1706_out1 XOR Logical_Operator_out1722_out1;

  Logical_Operator_out2739_out1 <= Logical_Operator_out1707_out1 XOR Logical_Operator_out1723_out1;

  Logical_Operator_out2740_out1 <= Logical_Operator_out1708_out1 XOR Logical_Operator_out1724_out1;

  Logical_Operator_out2741_out1 <= Logical_Operator_out1709_out1 XOR Logical_Operator_out1725_out1;

  Logical_Operator_out2742_out1 <= Logical_Operator_out1710_out1 XOR Logical_Operator_out1726_out1;

  Logical_Operator_out2743_out1 <= Logical_Operator_out1711_out1 XOR Logical_Operator_out1727_out1;

  Logical_Operator_out2744_out1 <= Logical_Operator_out1712_out1 XOR Logical_Operator_out1728_out1;

  Logical_Operator_out2745_out1 <= Logical_Operator_out1197_out1 XOR Logical_Operator_out1213_out1;

  Logical_Operator_out2746_out1 <= Logical_Operator_out1198_out1 XOR Logical_Operator_out1214_out1;

  Logical_Operator_out2747_out1 <= Logical_Operator_out1199_out1 XOR Logical_Operator_out1215_out1;

  Logical_Operator_out2748_out1 <= Logical_Operator_out1200_out1 XOR Logical_Operator_out1216_out1;

  Logical_Operator_out2749_out1 <= Logical_Operator_out687_out1 XOR Logical_Operator_out703_out1;

  Logical_Operator_out2750_out1 <= Logical_Operator_out688_out1 XOR Logical_Operator_out704_out1;

  Logical_Operator_out2751_out1 <= Logical_Operator_out176_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out2752_out1 <= in352 XOR in384;

  Logical_Operator_out2753_out1 <= Logical_Operator_out2241_out1 XOR Logical_Operator_out2257_out1;

  Logical_Operator_out2754_out1 <= Logical_Operator_out2242_out1 XOR Logical_Operator_out2258_out1;

  Logical_Operator_out2755_out1 <= Logical_Operator_out2243_out1 XOR Logical_Operator_out2259_out1;

  Logical_Operator_out2756_out1 <= Logical_Operator_out2244_out1 XOR Logical_Operator_out2260_out1;

  Logical_Operator_out2757_out1 <= Logical_Operator_out2245_out1 XOR Logical_Operator_out2261_out1;

  Logical_Operator_out2758_out1 <= Logical_Operator_out2246_out1 XOR Logical_Operator_out2262_out1;

  Logical_Operator_out2759_out1 <= Logical_Operator_out2247_out1 XOR Logical_Operator_out2263_out1;

  Logical_Operator_out2760_out1 <= Logical_Operator_out2248_out1 XOR Logical_Operator_out2264_out1;

  Logical_Operator_out2761_out1 <= Logical_Operator_out2249_out1 XOR Logical_Operator_out2265_out1;

  Logical_Operator_out2762_out1 <= Logical_Operator_out2250_out1 XOR Logical_Operator_out2266_out1;

  Logical_Operator_out2763_out1 <= Logical_Operator_out2251_out1 XOR Logical_Operator_out2267_out1;

  Logical_Operator_out2764_out1 <= Logical_Operator_out2252_out1 XOR Logical_Operator_out2268_out1;

  Logical_Operator_out2765_out1 <= Logical_Operator_out2253_out1 XOR Logical_Operator_out2269_out1;

  Logical_Operator_out2766_out1 <= Logical_Operator_out2254_out1 XOR Logical_Operator_out2270_out1;

  Logical_Operator_out2767_out1 <= Logical_Operator_out2255_out1 XOR Logical_Operator_out2271_out1;

  Logical_Operator_out2768_out1 <= Logical_Operator_out2256_out1 XOR Logical_Operator_out2272_out1;

  Logical_Operator_out2769_out1 <= Logical_Operator_out1737_out1 XOR Logical_Operator_out1753_out1;

  Logical_Operator_out2770_out1 <= Logical_Operator_out1738_out1 XOR Logical_Operator_out1754_out1;

  Logical_Operator_out2771_out1 <= Logical_Operator_out1739_out1 XOR Logical_Operator_out1755_out1;

  Logical_Operator_out2772_out1 <= Logical_Operator_out1740_out1 XOR Logical_Operator_out1756_out1;

  Logical_Operator_out2773_out1 <= Logical_Operator_out1741_out1 XOR Logical_Operator_out1757_out1;

  Logical_Operator_out2774_out1 <= Logical_Operator_out1742_out1 XOR Logical_Operator_out1758_out1;

  Logical_Operator_out2775_out1 <= Logical_Operator_out1743_out1 XOR Logical_Operator_out1759_out1;

  Logical_Operator_out2776_out1 <= Logical_Operator_out1744_out1 XOR Logical_Operator_out1760_out1;

  Logical_Operator_out2777_out1 <= Logical_Operator_out1229_out1 XOR Logical_Operator_out1245_out1;

  Logical_Operator_out2778_out1 <= Logical_Operator_out1230_out1 XOR Logical_Operator_out1246_out1;

  Logical_Operator_out2779_out1 <= Logical_Operator_out1231_out1 XOR Logical_Operator_out1247_out1;

  Logical_Operator_out2780_out1 <= Logical_Operator_out1232_out1 XOR Logical_Operator_out1248_out1;

  Logical_Operator_out2781_out1 <= Logical_Operator_out719_out1 XOR Logical_Operator_out735_out1;

  Logical_Operator_out2782_out1 <= Logical_Operator_out720_out1 XOR Logical_Operator_out736_out1;

  Logical_Operator_out2783_out1 <= Logical_Operator_out208_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out2784_out1 <= in416 XOR in448;

  Logical_Operator_out2785_out1 <= Logical_Operator_out2273_out1 XOR Logical_Operator_out2289_out1;

  Logical_Operator_out2786_out1 <= Logical_Operator_out2274_out1 XOR Logical_Operator_out2290_out1;

  Logical_Operator_out2787_out1 <= Logical_Operator_out2275_out1 XOR Logical_Operator_out2291_out1;

  Logical_Operator_out2788_out1 <= Logical_Operator_out2276_out1 XOR Logical_Operator_out2292_out1;

  Logical_Operator_out2789_out1 <= Logical_Operator_out2277_out1 XOR Logical_Operator_out2293_out1;

  Logical_Operator_out2790_out1 <= Logical_Operator_out2278_out1 XOR Logical_Operator_out2294_out1;

  Logical_Operator_out2791_out1 <= Logical_Operator_out2279_out1 XOR Logical_Operator_out2295_out1;

  Logical_Operator_out2792_out1 <= Logical_Operator_out2280_out1 XOR Logical_Operator_out2296_out1;

  Logical_Operator_out2793_out1 <= Logical_Operator_out2281_out1 XOR Logical_Operator_out2297_out1;

  Logical_Operator_out2794_out1 <= Logical_Operator_out2282_out1 XOR Logical_Operator_out2298_out1;

  Logical_Operator_out2795_out1 <= Logical_Operator_out2283_out1 XOR Logical_Operator_out2299_out1;

  Logical_Operator_out2796_out1 <= Logical_Operator_out2284_out1 XOR Logical_Operator_out2300_out1;

  Logical_Operator_out2797_out1 <= Logical_Operator_out2285_out1 XOR Logical_Operator_out2301_out1;

  Logical_Operator_out2798_out1 <= Logical_Operator_out2286_out1 XOR Logical_Operator_out2302_out1;

  Logical_Operator_out2799_out1 <= Logical_Operator_out2287_out1 XOR Logical_Operator_out2303_out1;

  Logical_Operator_out2800_out1 <= Logical_Operator_out2288_out1 XOR Logical_Operator_out2304_out1;

  Logical_Operator_out2801_out1 <= Logical_Operator_out1769_out1 XOR Logical_Operator_out1785_out1;

  Logical_Operator_out2802_out1 <= Logical_Operator_out1770_out1 XOR Logical_Operator_out1786_out1;

  Logical_Operator_out2803_out1 <= Logical_Operator_out1771_out1 XOR Logical_Operator_out1787_out1;

  Logical_Operator_out2804_out1 <= Logical_Operator_out1772_out1 XOR Logical_Operator_out1788_out1;

  Logical_Operator_out2805_out1 <= Logical_Operator_out1773_out1 XOR Logical_Operator_out1789_out1;

  Logical_Operator_out2806_out1 <= Logical_Operator_out1774_out1 XOR Logical_Operator_out1790_out1;

  Logical_Operator_out2807_out1 <= Logical_Operator_out1775_out1 XOR Logical_Operator_out1791_out1;

  Logical_Operator_out2808_out1 <= Logical_Operator_out1776_out1 XOR Logical_Operator_out1792_out1;

  Logical_Operator_out2809_out1 <= Logical_Operator_out1261_out1 XOR Logical_Operator_out1277_out1;

  Logical_Operator_out2810_out1 <= Logical_Operator_out1262_out1 XOR Logical_Operator_out1278_out1;

  Logical_Operator_out2811_out1 <= Logical_Operator_out1263_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out2812_out1 <= Logical_Operator_out1264_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out2813_out1 <= Logical_Operator_out751_out1 XOR Logical_Operator_out767_out1;

  Logical_Operator_out2814_out1 <= Logical_Operator_out752_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out2815_out1 <= Logical_Operator_out240_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out2816_out1 <= in480 XOR in512;

  Logical_Operator_out2817_out1 <= Logical_Operator_out2305_out1 XOR Logical_Operator_out2321_out1;

  Logical_Operator_out2818_out1 <= Logical_Operator_out2306_out1 XOR Logical_Operator_out2322_out1;

  Logical_Operator_out2819_out1 <= Logical_Operator_out2307_out1 XOR Logical_Operator_out2323_out1;

  Logical_Operator_out2820_out1 <= Logical_Operator_out2308_out1 XOR Logical_Operator_out2324_out1;

  Logical_Operator_out2821_out1 <= Logical_Operator_out2309_out1 XOR Logical_Operator_out2325_out1;

  Logical_Operator_out2822_out1 <= Logical_Operator_out2310_out1 XOR Logical_Operator_out2326_out1;

  Logical_Operator_out2823_out1 <= Logical_Operator_out2311_out1 XOR Logical_Operator_out2327_out1;

  Logical_Operator_out2824_out1 <= Logical_Operator_out2312_out1 XOR Logical_Operator_out2328_out1;

  Logical_Operator_out2825_out1 <= Logical_Operator_out2313_out1 XOR Logical_Operator_out2329_out1;

  Logical_Operator_out2826_out1 <= Logical_Operator_out2314_out1 XOR Logical_Operator_out2330_out1;

  Logical_Operator_out2827_out1 <= Logical_Operator_out2315_out1 XOR Logical_Operator_out2331_out1;

  Logical_Operator_out2828_out1 <= Logical_Operator_out2316_out1 XOR Logical_Operator_out2332_out1;

  Logical_Operator_out2829_out1 <= Logical_Operator_out2317_out1 XOR Logical_Operator_out2333_out1;

  Logical_Operator_out2830_out1 <= Logical_Operator_out2318_out1 XOR Logical_Operator_out2334_out1;

  Logical_Operator_out2831_out1 <= Logical_Operator_out2319_out1 XOR Logical_Operator_out2335_out1;

  Logical_Operator_out2832_out1 <= Logical_Operator_out2320_out1 XOR Logical_Operator_out2336_out1;

  Logical_Operator_out2833_out1 <= Logical_Operator_out1801_out1 XOR Logical_Operator_out1817_out1;

  Logical_Operator_out2834_out1 <= Logical_Operator_out1802_out1 XOR Logical_Operator_out1818_out1;

  Logical_Operator_out2835_out1 <= Logical_Operator_out1803_out1 XOR Logical_Operator_out1819_out1;

  Logical_Operator_out2836_out1 <= Logical_Operator_out1804_out1 XOR Logical_Operator_out1820_out1;

  Logical_Operator_out2837_out1 <= Logical_Operator_out1805_out1 XOR Logical_Operator_out1821_out1;

  Logical_Operator_out2838_out1 <= Logical_Operator_out1806_out1 XOR Logical_Operator_out1822_out1;

  Logical_Operator_out2839_out1 <= Logical_Operator_out1807_out1 XOR Logical_Operator_out1823_out1;

  Logical_Operator_out2840_out1 <= Logical_Operator_out1808_out1 XOR Logical_Operator_out1824_out1;

  Logical_Operator_out2841_out1 <= Logical_Operator_out1293_out1 XOR Logical_Operator_out1309_out1;

  Logical_Operator_out2842_out1 <= Logical_Operator_out1294_out1 XOR Logical_Operator_out1310_out1;

  Logical_Operator_out2843_out1 <= Logical_Operator_out1295_out1 XOR Logical_Operator_out1311_out1;

  Logical_Operator_out2844_out1 <= Logical_Operator_out1296_out1 XOR Logical_Operator_out1312_out1;

  Logical_Operator_out2845_out1 <= Logical_Operator_out783_out1 XOR Logical_Operator_out799_out1;

  Logical_Operator_out2846_out1 <= Logical_Operator_out784_out1 XOR Logical_Operator_out800_out1;

  Logical_Operator_out2847_out1 <= Logical_Operator_out272_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out2848_out1 <= in544 XOR in576;

  Logical_Operator_out2849_out1 <= Logical_Operator_out2337_out1 XOR Logical_Operator_out2353_out1;

  Logical_Operator_out2850_out1 <= Logical_Operator_out2338_out1 XOR Logical_Operator_out2354_out1;

  Logical_Operator_out2851_out1 <= Logical_Operator_out2339_out1 XOR Logical_Operator_out2355_out1;

  Logical_Operator_out2852_out1 <= Logical_Operator_out2340_out1 XOR Logical_Operator_out2356_out1;

  Logical_Operator_out2853_out1 <= Logical_Operator_out2341_out1 XOR Logical_Operator_out2357_out1;

  Logical_Operator_out2854_out1 <= Logical_Operator_out2342_out1 XOR Logical_Operator_out2358_out1;

  Logical_Operator_out2855_out1 <= Logical_Operator_out2343_out1 XOR Logical_Operator_out2359_out1;

  Logical_Operator_out2856_out1 <= Logical_Operator_out2344_out1 XOR Logical_Operator_out2360_out1;

  Logical_Operator_out2857_out1 <= Logical_Operator_out2345_out1 XOR Logical_Operator_out2361_out1;

  Logical_Operator_out2858_out1 <= Logical_Operator_out2346_out1 XOR Logical_Operator_out2362_out1;

  Logical_Operator_out2859_out1 <= Logical_Operator_out2347_out1 XOR Logical_Operator_out2363_out1;

  Logical_Operator_out2860_out1 <= Logical_Operator_out2348_out1 XOR Logical_Operator_out2364_out1;

  Logical_Operator_out2861_out1 <= Logical_Operator_out2349_out1 XOR Logical_Operator_out2365_out1;

  Logical_Operator_out2862_out1 <= Logical_Operator_out2350_out1 XOR Logical_Operator_out2366_out1;

  Logical_Operator_out2863_out1 <= Logical_Operator_out2351_out1 XOR Logical_Operator_out2367_out1;

  Logical_Operator_out2864_out1 <= Logical_Operator_out2352_out1 XOR Logical_Operator_out2368_out1;

  Logical_Operator_out2865_out1 <= Logical_Operator_out1833_out1 XOR Logical_Operator_out1849_out1;

  Logical_Operator_out2866_out1 <= Logical_Operator_out1834_out1 XOR Logical_Operator_out1850_out1;

  Logical_Operator_out2867_out1 <= Logical_Operator_out1835_out1 XOR Logical_Operator_out1851_out1;

  Logical_Operator_out2868_out1 <= Logical_Operator_out1836_out1 XOR Logical_Operator_out1852_out1;

  Logical_Operator_out2869_out1 <= Logical_Operator_out1837_out1 XOR Logical_Operator_out1853_out1;

  Logical_Operator_out2870_out1 <= Logical_Operator_out1838_out1 XOR Logical_Operator_out1854_out1;

  Logical_Operator_out2871_out1 <= Logical_Operator_out1839_out1 XOR Logical_Operator_out1855_out1;

  Logical_Operator_out2872_out1 <= Logical_Operator_out1840_out1 XOR Logical_Operator_out1856_out1;

  Logical_Operator_out2873_out1 <= Logical_Operator_out1325_out1 XOR Logical_Operator_out1341_out1;

  Logical_Operator_out2874_out1 <= Logical_Operator_out1326_out1 XOR Logical_Operator_out1342_out1;

  Logical_Operator_out2875_out1 <= Logical_Operator_out1327_out1 XOR Logical_Operator_out1343_out1;

  Logical_Operator_out2876_out1 <= Logical_Operator_out1328_out1 XOR Logical_Operator_out1344_out1;

  Logical_Operator_out2877_out1 <= Logical_Operator_out815_out1 XOR Logical_Operator_out831_out1;

  Logical_Operator_out2878_out1 <= Logical_Operator_out816_out1 XOR Logical_Operator_out832_out1;

  Logical_Operator_out2879_out1 <= Logical_Operator_out304_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out2880_out1 <= in608 XOR in640;

  Logical_Operator_out2881_out1 <= Logical_Operator_out2369_out1 XOR Logical_Operator_out2385_out1;

  Logical_Operator_out2882_out1 <= Logical_Operator_out2370_out1 XOR Logical_Operator_out2386_out1;

  Logical_Operator_out2883_out1 <= Logical_Operator_out2371_out1 XOR Logical_Operator_out2387_out1;

  Logical_Operator_out2884_out1 <= Logical_Operator_out2372_out1 XOR Logical_Operator_out2388_out1;

  Logical_Operator_out2885_out1 <= Logical_Operator_out2373_out1 XOR Logical_Operator_out2389_out1;

  Logical_Operator_out2886_out1 <= Logical_Operator_out2374_out1 XOR Logical_Operator_out2390_out1;

  Logical_Operator_out2887_out1 <= Logical_Operator_out2375_out1 XOR Logical_Operator_out2391_out1;

  Logical_Operator_out2888_out1 <= Logical_Operator_out2376_out1 XOR Logical_Operator_out2392_out1;

  Logical_Operator_out2889_out1 <= Logical_Operator_out2377_out1 XOR Logical_Operator_out2393_out1;

  Logical_Operator_out2890_out1 <= Logical_Operator_out2378_out1 XOR Logical_Operator_out2394_out1;

  Logical_Operator_out2891_out1 <= Logical_Operator_out2379_out1 XOR Logical_Operator_out2395_out1;

  Logical_Operator_out2892_out1 <= Logical_Operator_out2380_out1 XOR Logical_Operator_out2396_out1;

  Logical_Operator_out2893_out1 <= Logical_Operator_out2381_out1 XOR Logical_Operator_out2397_out1;

  Logical_Operator_out2894_out1 <= Logical_Operator_out2382_out1 XOR Logical_Operator_out2398_out1;

  Logical_Operator_out2895_out1 <= Logical_Operator_out2383_out1 XOR Logical_Operator_out2399_out1;

  Logical_Operator_out2896_out1 <= Logical_Operator_out2384_out1 XOR Logical_Operator_out2400_out1;

  Logical_Operator_out2897_out1 <= Logical_Operator_out1865_out1 XOR Logical_Operator_out1881_out1;

  Logical_Operator_out2898_out1 <= Logical_Operator_out1866_out1 XOR Logical_Operator_out1882_out1;

  Logical_Operator_out2899_out1 <= Logical_Operator_out1867_out1 XOR Logical_Operator_out1883_out1;

  Logical_Operator_out2900_out1 <= Logical_Operator_out1868_out1 XOR Logical_Operator_out1884_out1;

  Logical_Operator_out2901_out1 <= Logical_Operator_out1869_out1 XOR Logical_Operator_out1885_out1;

  Logical_Operator_out2902_out1 <= Logical_Operator_out1870_out1 XOR Logical_Operator_out1886_out1;

  Logical_Operator_out2903_out1 <= Logical_Operator_out1871_out1 XOR Logical_Operator_out1887_out1;

  Logical_Operator_out2904_out1 <= Logical_Operator_out1872_out1 XOR Logical_Operator_out1888_out1;

  Logical_Operator_out2905_out1 <= Logical_Operator_out1357_out1 XOR Logical_Operator_out1373_out1;

  Logical_Operator_out2906_out1 <= Logical_Operator_out1358_out1 XOR Logical_Operator_out1374_out1;

  Logical_Operator_out2907_out1 <= Logical_Operator_out1359_out1 XOR Logical_Operator_out1375_out1;

  Logical_Operator_out2908_out1 <= Logical_Operator_out1360_out1 XOR Logical_Operator_out1376_out1;

  Logical_Operator_out2909_out1 <= Logical_Operator_out847_out1 XOR Logical_Operator_out863_out1;

  Logical_Operator_out2910_out1 <= Logical_Operator_out848_out1 XOR Logical_Operator_out864_out1;

  Logical_Operator_out2911_out1 <= Logical_Operator_out336_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out2912_out1 <= in672 XOR in704;

  Logical_Operator_out2913_out1 <= Logical_Operator_out2401_out1 XOR Logical_Operator_out2417_out1;

  Logical_Operator_out2914_out1 <= Logical_Operator_out2402_out1 XOR Logical_Operator_out2418_out1;

  Logical_Operator_out2915_out1 <= Logical_Operator_out2403_out1 XOR Logical_Operator_out2419_out1;

  Logical_Operator_out2916_out1 <= Logical_Operator_out2404_out1 XOR Logical_Operator_out2420_out1;

  Logical_Operator_out2917_out1 <= Logical_Operator_out2405_out1 XOR Logical_Operator_out2421_out1;

  Logical_Operator_out2918_out1 <= Logical_Operator_out2406_out1 XOR Logical_Operator_out2422_out1;

  Logical_Operator_out2919_out1 <= Logical_Operator_out2407_out1 XOR Logical_Operator_out2423_out1;

  Logical_Operator_out2920_out1 <= Logical_Operator_out2408_out1 XOR Logical_Operator_out2424_out1;

  Logical_Operator_out2921_out1 <= Logical_Operator_out2409_out1 XOR Logical_Operator_out2425_out1;

  Logical_Operator_out2922_out1 <= Logical_Operator_out2410_out1 XOR Logical_Operator_out2426_out1;

  Logical_Operator_out2923_out1 <= Logical_Operator_out2411_out1 XOR Logical_Operator_out2427_out1;

  Logical_Operator_out2924_out1 <= Logical_Operator_out2412_out1 XOR Logical_Operator_out2428_out1;

  Logical_Operator_out2925_out1 <= Logical_Operator_out2413_out1 XOR Logical_Operator_out2429_out1;

  Logical_Operator_out2926_out1 <= Logical_Operator_out2414_out1 XOR Logical_Operator_out2430_out1;

  Logical_Operator_out2927_out1 <= Logical_Operator_out2415_out1 XOR Logical_Operator_out2431_out1;

  Logical_Operator_out2928_out1 <= Logical_Operator_out2416_out1 XOR Logical_Operator_out2432_out1;

  Logical_Operator_out2929_out1 <= Logical_Operator_out1897_out1 XOR Logical_Operator_out1913_out1;

  Logical_Operator_out2930_out1 <= Logical_Operator_out1898_out1 XOR Logical_Operator_out1914_out1;

  Logical_Operator_out2931_out1 <= Logical_Operator_out1899_out1 XOR Logical_Operator_out1915_out1;

  Logical_Operator_out2932_out1 <= Logical_Operator_out1900_out1 XOR Logical_Operator_out1916_out1;

  Logical_Operator_out2933_out1 <= Logical_Operator_out1901_out1 XOR Logical_Operator_out1917_out1;

  Logical_Operator_out2934_out1 <= Logical_Operator_out1902_out1 XOR Logical_Operator_out1918_out1;

  Logical_Operator_out2935_out1 <= Logical_Operator_out1903_out1 XOR Logical_Operator_out1919_out1;

  Logical_Operator_out2936_out1 <= Logical_Operator_out1904_out1 XOR Logical_Operator_out1920_out1;

  Logical_Operator_out2937_out1 <= Logical_Operator_out1389_out1 XOR Logical_Operator_out1405_out1;

  Logical_Operator_out2938_out1 <= Logical_Operator_out1390_out1 XOR Logical_Operator_out1406_out1;

  Logical_Operator_out2939_out1 <= Logical_Operator_out1391_out1 XOR Logical_Operator_out1407_out1;

  Logical_Operator_out2940_out1 <= Logical_Operator_out1392_out1 XOR Logical_Operator_out1408_out1;

  Logical_Operator_out2941_out1 <= Logical_Operator_out879_out1 XOR Logical_Operator_out895_out1;

  Logical_Operator_out2942_out1 <= Logical_Operator_out880_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out2943_out1 <= Logical_Operator_out368_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out2944_out1 <= in736 XOR in768;

  Logical_Operator_out2945_out1 <= Logical_Operator_out2433_out1 XOR Logical_Operator_out2449_out1;

  Logical_Operator_out2946_out1 <= Logical_Operator_out2434_out1 XOR Logical_Operator_out2450_out1;

  Logical_Operator_out2947_out1 <= Logical_Operator_out2435_out1 XOR Logical_Operator_out2451_out1;

  Logical_Operator_out2948_out1 <= Logical_Operator_out2436_out1 XOR Logical_Operator_out2452_out1;

  Logical_Operator_out2949_out1 <= Logical_Operator_out2437_out1 XOR Logical_Operator_out2453_out1;

  Logical_Operator_out2950_out1 <= Logical_Operator_out2438_out1 XOR Logical_Operator_out2454_out1;

  Logical_Operator_out2951_out1 <= Logical_Operator_out2439_out1 XOR Logical_Operator_out2455_out1;

  Logical_Operator_out2952_out1 <= Logical_Operator_out2440_out1 XOR Logical_Operator_out2456_out1;

  Logical_Operator_out2953_out1 <= Logical_Operator_out2441_out1 XOR Logical_Operator_out2457_out1;

  Logical_Operator_out2954_out1 <= Logical_Operator_out2442_out1 XOR Logical_Operator_out2458_out1;

  Logical_Operator_out2955_out1 <= Logical_Operator_out2443_out1 XOR Logical_Operator_out2459_out1;

  Logical_Operator_out2956_out1 <= Logical_Operator_out2444_out1 XOR Logical_Operator_out2460_out1;

  Logical_Operator_out2957_out1 <= Logical_Operator_out2445_out1 XOR Logical_Operator_out2461_out1;

  Logical_Operator_out2958_out1 <= Logical_Operator_out2446_out1 XOR Logical_Operator_out2462_out1;

  Logical_Operator_out2959_out1 <= Logical_Operator_out2447_out1 XOR Logical_Operator_out2463_out1;

  Logical_Operator_out2960_out1 <= Logical_Operator_out2448_out1 XOR Logical_Operator_out2464_out1;

  Logical_Operator_out2961_out1 <= Logical_Operator_out1929_out1 XOR Logical_Operator_out1945_out1;

  Logical_Operator_out2962_out1 <= Logical_Operator_out1930_out1 XOR Logical_Operator_out1946_out1;

  Logical_Operator_out2963_out1 <= Logical_Operator_out1931_out1 XOR Logical_Operator_out1947_out1;

  Logical_Operator_out2964_out1 <= Logical_Operator_out1932_out1 XOR Logical_Operator_out1948_out1;

  Logical_Operator_out2965_out1 <= Logical_Operator_out1933_out1 XOR Logical_Operator_out1949_out1;

  Logical_Operator_out2966_out1 <= Logical_Operator_out1934_out1 XOR Logical_Operator_out1950_out1;

  Logical_Operator_out2967_out1 <= Logical_Operator_out1935_out1 XOR Logical_Operator_out1951_out1;

  Logical_Operator_out2968_out1 <= Logical_Operator_out1936_out1 XOR Logical_Operator_out1952_out1;

  Logical_Operator_out2969_out1 <= Logical_Operator_out1421_out1 XOR Logical_Operator_out1437_out1;

  Logical_Operator_out2970_out1 <= Logical_Operator_out1422_out1 XOR Logical_Operator_out1438_out1;

  Logical_Operator_out2971_out1 <= Logical_Operator_out1423_out1 XOR Logical_Operator_out1439_out1;

  Logical_Operator_out2972_out1 <= Logical_Operator_out1424_out1 XOR Logical_Operator_out1440_out1;

  Logical_Operator_out2973_out1 <= Logical_Operator_out911_out1 XOR Logical_Operator_out927_out1;

  Logical_Operator_out2974_out1 <= Logical_Operator_out912_out1 XOR Logical_Operator_out928_out1;

  Logical_Operator_out2975_out1 <= Logical_Operator_out400_out1 XOR Logical_Operator_out416_out1;

  Logical_Operator_out2976_out1 <= in800 XOR in832;

  Logical_Operator_out2977_out1 <= Logical_Operator_out2465_out1 XOR Logical_Operator_out2481_out1;

  Logical_Operator_out2978_out1 <= Logical_Operator_out2466_out1 XOR Logical_Operator_out2482_out1;

  Logical_Operator_out2979_out1 <= Logical_Operator_out2467_out1 XOR Logical_Operator_out2483_out1;

  Logical_Operator_out2980_out1 <= Logical_Operator_out2468_out1 XOR Logical_Operator_out2484_out1;

  Logical_Operator_out2981_out1 <= Logical_Operator_out2469_out1 XOR Logical_Operator_out2485_out1;

  Logical_Operator_out2982_out1 <= Logical_Operator_out2470_out1 XOR Logical_Operator_out2486_out1;

  Logical_Operator_out2983_out1 <= Logical_Operator_out2471_out1 XOR Logical_Operator_out2487_out1;

  Logical_Operator_out2984_out1 <= Logical_Operator_out2472_out1 XOR Logical_Operator_out2488_out1;

  Logical_Operator_out2985_out1 <= Logical_Operator_out2473_out1 XOR Logical_Operator_out2489_out1;

  Logical_Operator_out2986_out1 <= Logical_Operator_out2474_out1 XOR Logical_Operator_out2490_out1;

  Logical_Operator_out2987_out1 <= Logical_Operator_out2475_out1 XOR Logical_Operator_out2491_out1;

  Logical_Operator_out2988_out1 <= Logical_Operator_out2476_out1 XOR Logical_Operator_out2492_out1;

  Logical_Operator_out2989_out1 <= Logical_Operator_out2477_out1 XOR Logical_Operator_out2493_out1;

  Logical_Operator_out2990_out1 <= Logical_Operator_out2478_out1 XOR Logical_Operator_out2494_out1;

  Logical_Operator_out2991_out1 <= Logical_Operator_out2479_out1 XOR Logical_Operator_out2495_out1;

  Logical_Operator_out2992_out1 <= Logical_Operator_out2480_out1 XOR Logical_Operator_out2496_out1;

  Logical_Operator_out2993_out1 <= Logical_Operator_out1961_out1 XOR Logical_Operator_out1977_out1;

  Logical_Operator_out2994_out1 <= Logical_Operator_out1962_out1 XOR Logical_Operator_out1978_out1;

  Logical_Operator_out2995_out1 <= Logical_Operator_out1963_out1 XOR Logical_Operator_out1979_out1;

  Logical_Operator_out2996_out1 <= Logical_Operator_out1964_out1 XOR Logical_Operator_out1980_out1;

  Logical_Operator_out2997_out1 <= Logical_Operator_out1965_out1 XOR Logical_Operator_out1981_out1;

  Logical_Operator_out2998_out1 <= Logical_Operator_out1966_out1 XOR Logical_Operator_out1982_out1;

  Logical_Operator_out2999_out1 <= Logical_Operator_out1967_out1 XOR Logical_Operator_out1983_out1;

  Logical_Operator_out3000_out1 <= Logical_Operator_out1968_out1 XOR Logical_Operator_out1984_out1;

  Logical_Operator_out3001_out1 <= Logical_Operator_out1453_out1 XOR Logical_Operator_out1469_out1;

  Logical_Operator_out3002_out1 <= Logical_Operator_out1454_out1 XOR Logical_Operator_out1470_out1;

  Logical_Operator_out3003_out1 <= Logical_Operator_out1455_out1 XOR Logical_Operator_out1471_out1;

  Logical_Operator_out3004_out1 <= Logical_Operator_out1456_out1 XOR Logical_Operator_out1472_out1;

  Logical_Operator_out3005_out1 <= Logical_Operator_out943_out1 XOR Logical_Operator_out959_out1;

  Logical_Operator_out3006_out1 <= Logical_Operator_out944_out1 XOR Logical_Operator_out960_out1;

  Logical_Operator_out3007_out1 <= Logical_Operator_out432_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out3008_out1 <= in864 XOR in896;

  Logical_Operator_out3009_out1 <= Logical_Operator_out2497_out1 XOR Logical_Operator_out2513_out1;

  Logical_Operator_out3010_out1 <= Logical_Operator_out2498_out1 XOR Logical_Operator_out2514_out1;

  Logical_Operator_out3011_out1 <= Logical_Operator_out2499_out1 XOR Logical_Operator_out2515_out1;

  Logical_Operator_out3012_out1 <= Logical_Operator_out2500_out1 XOR Logical_Operator_out2516_out1;

  Logical_Operator_out3013_out1 <= Logical_Operator_out2501_out1 XOR Logical_Operator_out2517_out1;

  Logical_Operator_out3014_out1 <= Logical_Operator_out2502_out1 XOR Logical_Operator_out2518_out1;

  Logical_Operator_out3015_out1 <= Logical_Operator_out2503_out1 XOR Logical_Operator_out2519_out1;

  Logical_Operator_out3016_out1 <= Logical_Operator_out2504_out1 XOR Logical_Operator_out2520_out1;

  Logical_Operator_out3017_out1 <= Logical_Operator_out2505_out1 XOR Logical_Operator_out2521_out1;

  Logical_Operator_out3018_out1 <= Logical_Operator_out2506_out1 XOR Logical_Operator_out2522_out1;

  Logical_Operator_out3019_out1 <= Logical_Operator_out2507_out1 XOR Logical_Operator_out2523_out1;

  Logical_Operator_out3020_out1 <= Logical_Operator_out2508_out1 XOR Logical_Operator_out2524_out1;

  Logical_Operator_out3021_out1 <= Logical_Operator_out2509_out1 XOR Logical_Operator_out2525_out1;

  Logical_Operator_out3022_out1 <= Logical_Operator_out2510_out1 XOR Logical_Operator_out2526_out1;

  Logical_Operator_out3023_out1 <= Logical_Operator_out2511_out1 XOR Logical_Operator_out2527_out1;

  Logical_Operator_out3024_out1 <= Logical_Operator_out2512_out1 XOR Logical_Operator_out2528_out1;

  Logical_Operator_out3025_out1 <= Logical_Operator_out1993_out1 XOR Logical_Operator_out2009_out1;

  Logical_Operator_out3026_out1 <= Logical_Operator_out1994_out1 XOR Logical_Operator_out2010_out1;

  Logical_Operator_out3027_out1 <= Logical_Operator_out1995_out1 XOR Logical_Operator_out2011_out1;

  Logical_Operator_out3028_out1 <= Logical_Operator_out1996_out1 XOR Logical_Operator_out2012_out1;

  Logical_Operator_out3029_out1 <= Logical_Operator_out1997_out1 XOR Logical_Operator_out2013_out1;

  Logical_Operator_out3030_out1 <= Logical_Operator_out1998_out1 XOR Logical_Operator_out2014_out1;

  Logical_Operator_out3031_out1 <= Logical_Operator_out1999_out1 XOR Logical_Operator_out2015_out1;

  Logical_Operator_out3032_out1 <= Logical_Operator_out2000_out1 XOR Logical_Operator_out2016_out1;

  Logical_Operator_out3033_out1 <= Logical_Operator_out1485_out1 XOR Logical_Operator_out1501_out1;

  Logical_Operator_out3034_out1 <= Logical_Operator_out1486_out1 XOR Logical_Operator_out1502_out1;

  Logical_Operator_out3035_out1 <= Logical_Operator_out1487_out1 XOR Logical_Operator_out1503_out1;

  Logical_Operator_out3036_out1 <= Logical_Operator_out1488_out1 XOR Logical_Operator_out1504_out1;

  Logical_Operator_out3037_out1 <= Logical_Operator_out975_out1 XOR Logical_Operator_out991_out1;

  Logical_Operator_out3038_out1 <= Logical_Operator_out976_out1 XOR Logical_Operator_out992_out1;

  Logical_Operator_out3039_out1 <= Logical_Operator_out464_out1 XOR Logical_Operator_out480_out1;

  Logical_Operator_out3040_out1 <= in928 XOR in960;

  Logical_Operator_out3041_out1 <= Logical_Operator_out2529_out1 XOR Logical_Operator_out2545_out1;

  Logical_Operator_out3042_out1 <= Logical_Operator_out2530_out1 XOR Logical_Operator_out2546_out1;

  Logical_Operator_out3043_out1 <= Logical_Operator_out2531_out1 XOR Logical_Operator_out2547_out1;

  Logical_Operator_out3044_out1 <= Logical_Operator_out2532_out1 XOR Logical_Operator_out2548_out1;

  Logical_Operator_out3045_out1 <= Logical_Operator_out2533_out1 XOR Logical_Operator_out2549_out1;

  Logical_Operator_out3046_out1 <= Logical_Operator_out2534_out1 XOR Logical_Operator_out2550_out1;

  Logical_Operator_out3047_out1 <= Logical_Operator_out2535_out1 XOR Logical_Operator_out2551_out1;

  Logical_Operator_out3048_out1 <= Logical_Operator_out2536_out1 XOR Logical_Operator_out2552_out1;

  Logical_Operator_out3049_out1 <= Logical_Operator_out2537_out1 XOR Logical_Operator_out2553_out1;

  Logical_Operator_out3050_out1 <= Logical_Operator_out2538_out1 XOR Logical_Operator_out2554_out1;

  Logical_Operator_out3051_out1 <= Logical_Operator_out2539_out1 XOR Logical_Operator_out2555_out1;

  Logical_Operator_out3052_out1 <= Logical_Operator_out2540_out1 XOR Logical_Operator_out2556_out1;

  Logical_Operator_out3053_out1 <= Logical_Operator_out2541_out1 XOR Logical_Operator_out2557_out1;

  Logical_Operator_out3054_out1 <= Logical_Operator_out2542_out1 XOR Logical_Operator_out2558_out1;

  Logical_Operator_out3055_out1 <= Logical_Operator_out2543_out1 XOR Logical_Operator_out2559_out1;

  Logical_Operator_out3056_out1 <= Logical_Operator_out2544_out1 XOR Logical_Operator_out2560_out1;

  Logical_Operator_out3057_out1 <= Logical_Operator_out2025_out1 XOR Logical_Operator_out2041_out1;

  Logical_Operator_out3058_out1 <= Logical_Operator_out2026_out1 XOR Logical_Operator_out2042_out1;

  Logical_Operator_out3059_out1 <= Logical_Operator_out2027_out1 XOR Logical_Operator_out2043_out1;

  Logical_Operator_out3060_out1 <= Logical_Operator_out2028_out1 XOR Logical_Operator_out2044_out1;

  Logical_Operator_out3061_out1 <= Logical_Operator_out2029_out1 XOR Logical_Operator_out2045_out1;

  Logical_Operator_out3062_out1 <= Logical_Operator_out2030_out1 XOR Logical_Operator_out2046_out1;

  Logical_Operator_out3063_out1 <= Logical_Operator_out2031_out1 XOR Logical_Operator_out2047_out1;

  Logical_Operator_out3064_out1 <= Logical_Operator_out2032_out1 XOR Logical_Operator_out2048_out1;

  Logical_Operator_out3065_out1 <= Logical_Operator_out1517_out1 XOR Logical_Operator_out1533_out1;

  Logical_Operator_out3066_out1 <= Logical_Operator_out1518_out1 XOR Logical_Operator_out1534_out1;

  Logical_Operator_out3067_out1 <= Logical_Operator_out1519_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out3068_out1 <= Logical_Operator_out1520_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out3069_out1 <= Logical_Operator_out1007_out1 XOR Logical_Operator_out1023_out1;

  Logical_Operator_out3070_out1 <= Logical_Operator_out1008_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out3071_out1 <= Logical_Operator_out496_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out3072_out1 <= in992 XOR in1024;

  Logical_Operator_out3073_out1 <= Logical_Operator_out2561_out1 XOR Logical_Operator_out2593_out1;

  Logical_Operator_out3074_out1 <= Logical_Operator_out2562_out1 XOR Logical_Operator_out2594_out1;

  Logical_Operator_out3075_out1 <= Logical_Operator_out2563_out1 XOR Logical_Operator_out2595_out1;

  Logical_Operator_out3076_out1 <= Logical_Operator_out2564_out1 XOR Logical_Operator_out2596_out1;

  Logical_Operator_out3077_out1 <= Logical_Operator_out2565_out1 XOR Logical_Operator_out2597_out1;

  Logical_Operator_out3078_out1 <= Logical_Operator_out2566_out1 XOR Logical_Operator_out2598_out1;

  Logical_Operator_out3079_out1 <= Logical_Operator_out2567_out1 XOR Logical_Operator_out2599_out1;

  Logical_Operator_out3080_out1 <= Logical_Operator_out2568_out1 XOR Logical_Operator_out2600_out1;

  Logical_Operator_out3081_out1 <= Logical_Operator_out2569_out1 XOR Logical_Operator_out2601_out1;

  Logical_Operator_out3082_out1 <= Logical_Operator_out2570_out1 XOR Logical_Operator_out2602_out1;

  Logical_Operator_out3083_out1 <= Logical_Operator_out2571_out1 XOR Logical_Operator_out2603_out1;

  Logical_Operator_out3084_out1 <= Logical_Operator_out2572_out1 XOR Logical_Operator_out2604_out1;

  Logical_Operator_out3085_out1 <= Logical_Operator_out2573_out1 XOR Logical_Operator_out2605_out1;

  Logical_Operator_out3086_out1 <= Logical_Operator_out2574_out1 XOR Logical_Operator_out2606_out1;

  Logical_Operator_out3087_out1 <= Logical_Operator_out2575_out1 XOR Logical_Operator_out2607_out1;

  Logical_Operator_out3088_out1 <= Logical_Operator_out2576_out1 XOR Logical_Operator_out2608_out1;

  Logical_Operator_out3089_out1 <= Logical_Operator_out2577_out1 XOR Logical_Operator_out2609_out1;

  Logical_Operator_out3090_out1 <= Logical_Operator_out2578_out1 XOR Logical_Operator_out2610_out1;

  Logical_Operator_out3091_out1 <= Logical_Operator_out2579_out1 XOR Logical_Operator_out2611_out1;

  Logical_Operator_out3092_out1 <= Logical_Operator_out2580_out1 XOR Logical_Operator_out2612_out1;

  Logical_Operator_out3093_out1 <= Logical_Operator_out2581_out1 XOR Logical_Operator_out2613_out1;

  Logical_Operator_out3094_out1 <= Logical_Operator_out2582_out1 XOR Logical_Operator_out2614_out1;

  Logical_Operator_out3095_out1 <= Logical_Operator_out2583_out1 XOR Logical_Operator_out2615_out1;

  Logical_Operator_out3096_out1 <= Logical_Operator_out2584_out1 XOR Logical_Operator_out2616_out1;

  Logical_Operator_out3097_out1 <= Logical_Operator_out2585_out1 XOR Logical_Operator_out2617_out1;

  Logical_Operator_out3098_out1 <= Logical_Operator_out2586_out1 XOR Logical_Operator_out2618_out1;

  Logical_Operator_out3099_out1 <= Logical_Operator_out2587_out1 XOR Logical_Operator_out2619_out1;

  Logical_Operator_out3100_out1 <= Logical_Operator_out2588_out1 XOR Logical_Operator_out2620_out1;

  Logical_Operator_out3101_out1 <= Logical_Operator_out2589_out1 XOR Logical_Operator_out2621_out1;

  Logical_Operator_out3102_out1 <= Logical_Operator_out2590_out1 XOR Logical_Operator_out2622_out1;

  Logical_Operator_out3103_out1 <= Logical_Operator_out2591_out1 XOR Logical_Operator_out2623_out1;

  Logical_Operator_out3104_out1 <= Logical_Operator_out2592_out1 XOR Logical_Operator_out2624_out1;

  Logical_Operator_out3105_out1 <= Logical_Operator_out2065_out1 XOR Logical_Operator_out2097_out1;

  Logical_Operator_out3106_out1 <= Logical_Operator_out2066_out1 XOR Logical_Operator_out2098_out1;

  Logical_Operator_out3107_out1 <= Logical_Operator_out2067_out1 XOR Logical_Operator_out2099_out1;

  Logical_Operator_out3108_out1 <= Logical_Operator_out2068_out1 XOR Logical_Operator_out2100_out1;

  Logical_Operator_out3109_out1 <= Logical_Operator_out2069_out1 XOR Logical_Operator_out2101_out1;

  Logical_Operator_out3110_out1 <= Logical_Operator_out2070_out1 XOR Logical_Operator_out2102_out1;

  Logical_Operator_out3111_out1 <= Logical_Operator_out2071_out1 XOR Logical_Operator_out2103_out1;

  Logical_Operator_out3112_out1 <= Logical_Operator_out2072_out1 XOR Logical_Operator_out2104_out1;

  Logical_Operator_out3113_out1 <= Logical_Operator_out2073_out1 XOR Logical_Operator_out2105_out1;

  Logical_Operator_out3114_out1 <= Logical_Operator_out2074_out1 XOR Logical_Operator_out2106_out1;

  Logical_Operator_out3115_out1 <= Logical_Operator_out2075_out1 XOR Logical_Operator_out2107_out1;

  Logical_Operator_out3116_out1 <= Logical_Operator_out2076_out1 XOR Logical_Operator_out2108_out1;

  Logical_Operator_out3117_out1 <= Logical_Operator_out2077_out1 XOR Logical_Operator_out2109_out1;

  Logical_Operator_out3118_out1 <= Logical_Operator_out2078_out1 XOR Logical_Operator_out2110_out1;

  Logical_Operator_out3119_out1 <= Logical_Operator_out2079_out1 XOR Logical_Operator_out2111_out1;

  Logical_Operator_out3120_out1 <= Logical_Operator_out2080_out1 XOR Logical_Operator_out2112_out1;

  Logical_Operator_out3121_out1 <= Logical_Operator_out1561_out1 XOR Logical_Operator_out1593_out1;

  Logical_Operator_out3122_out1 <= Logical_Operator_out1562_out1 XOR Logical_Operator_out1594_out1;

  Logical_Operator_out3123_out1 <= Logical_Operator_out1563_out1 XOR Logical_Operator_out1595_out1;

  Logical_Operator_out3124_out1 <= Logical_Operator_out1564_out1 XOR Logical_Operator_out1596_out1;

  Logical_Operator_out3125_out1 <= Logical_Operator_out1565_out1 XOR Logical_Operator_out1597_out1;

  Logical_Operator_out3126_out1 <= Logical_Operator_out1566_out1 XOR Logical_Operator_out1598_out1;

  Logical_Operator_out3127_out1 <= Logical_Operator_out1567_out1 XOR Logical_Operator_out1599_out1;

  Logical_Operator_out3128_out1 <= Logical_Operator_out1568_out1 XOR Logical_Operator_out1600_out1;

  Logical_Operator_out3129_out1 <= Logical_Operator_out1053_out1 XOR Logical_Operator_out1085_out1;

  Logical_Operator_out3130_out1 <= Logical_Operator_out1054_out1 XOR Logical_Operator_out1086_out1;

  Logical_Operator_out3131_out1 <= Logical_Operator_out1055_out1 XOR Logical_Operator_out1087_out1;

  Logical_Operator_out3132_out1 <= Logical_Operator_out1056_out1 XOR Logical_Operator_out1088_out1;

  Logical_Operator_out3133_out1 <= Logical_Operator_out543_out1 XOR Logical_Operator_out575_out1;

  Logical_Operator_out3134_out1 <= Logical_Operator_out544_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out3135_out1 <= Logical_Operator_out32_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out3136_out1 <= in64 XOR in128;

  Logical_Operator_out3137_out1 <= Logical_Operator_out2625_out1 XOR Logical_Operator_out2657_out1;

  Logical_Operator_out3138_out1 <= Logical_Operator_out2626_out1 XOR Logical_Operator_out2658_out1;

  Logical_Operator_out3139_out1 <= Logical_Operator_out2627_out1 XOR Logical_Operator_out2659_out1;

  Logical_Operator_out3140_out1 <= Logical_Operator_out2628_out1 XOR Logical_Operator_out2660_out1;

  Logical_Operator_out3141_out1 <= Logical_Operator_out2629_out1 XOR Logical_Operator_out2661_out1;

  Logical_Operator_out3142_out1 <= Logical_Operator_out2630_out1 XOR Logical_Operator_out2662_out1;

  Logical_Operator_out3143_out1 <= Logical_Operator_out2631_out1 XOR Logical_Operator_out2663_out1;

  Logical_Operator_out3144_out1 <= Logical_Operator_out2632_out1 XOR Logical_Operator_out2664_out1;

  Logical_Operator_out3145_out1 <= Logical_Operator_out2633_out1 XOR Logical_Operator_out2665_out1;

  Logical_Operator_out3146_out1 <= Logical_Operator_out2634_out1 XOR Logical_Operator_out2666_out1;

  Logical_Operator_out3147_out1 <= Logical_Operator_out2635_out1 XOR Logical_Operator_out2667_out1;

  Logical_Operator_out3148_out1 <= Logical_Operator_out2636_out1 XOR Logical_Operator_out2668_out1;

  Logical_Operator_out3149_out1 <= Logical_Operator_out2637_out1 XOR Logical_Operator_out2669_out1;

  Logical_Operator_out3150_out1 <= Logical_Operator_out2638_out1 XOR Logical_Operator_out2670_out1;

  Logical_Operator_out3151_out1 <= Logical_Operator_out2639_out1 XOR Logical_Operator_out2671_out1;

  Logical_Operator_out3152_out1 <= Logical_Operator_out2640_out1 XOR Logical_Operator_out2672_out1;

  Logical_Operator_out3153_out1 <= Logical_Operator_out2641_out1 XOR Logical_Operator_out2673_out1;

  Logical_Operator_out3154_out1 <= Logical_Operator_out2642_out1 XOR Logical_Operator_out2674_out1;

  Logical_Operator_out3155_out1 <= Logical_Operator_out2643_out1 XOR Logical_Operator_out2675_out1;

  Logical_Operator_out3156_out1 <= Logical_Operator_out2644_out1 XOR Logical_Operator_out2676_out1;

  Logical_Operator_out3157_out1 <= Logical_Operator_out2645_out1 XOR Logical_Operator_out2677_out1;

  Logical_Operator_out3158_out1 <= Logical_Operator_out2646_out1 XOR Logical_Operator_out2678_out1;

  Logical_Operator_out3159_out1 <= Logical_Operator_out2647_out1 XOR Logical_Operator_out2679_out1;

  Logical_Operator_out3160_out1 <= Logical_Operator_out2648_out1 XOR Logical_Operator_out2680_out1;

  Logical_Operator_out3161_out1 <= Logical_Operator_out2649_out1 XOR Logical_Operator_out2681_out1;

  Logical_Operator_out3162_out1 <= Logical_Operator_out2650_out1 XOR Logical_Operator_out2682_out1;

  Logical_Operator_out3163_out1 <= Logical_Operator_out2651_out1 XOR Logical_Operator_out2683_out1;

  Logical_Operator_out3164_out1 <= Logical_Operator_out2652_out1 XOR Logical_Operator_out2684_out1;

  Logical_Operator_out3165_out1 <= Logical_Operator_out2653_out1 XOR Logical_Operator_out2685_out1;

  Logical_Operator_out3166_out1 <= Logical_Operator_out2654_out1 XOR Logical_Operator_out2686_out1;

  Logical_Operator_out3167_out1 <= Logical_Operator_out2655_out1 XOR Logical_Operator_out2687_out1;

  Logical_Operator_out3168_out1 <= Logical_Operator_out2656_out1 XOR Logical_Operator_out2688_out1;

  Logical_Operator_out3169_out1 <= Logical_Operator_out2129_out1 XOR Logical_Operator_out2161_out1;

  Logical_Operator_out3170_out1 <= Logical_Operator_out2130_out1 XOR Logical_Operator_out2162_out1;

  Logical_Operator_out3171_out1 <= Logical_Operator_out2131_out1 XOR Logical_Operator_out2163_out1;

  Logical_Operator_out3172_out1 <= Logical_Operator_out2132_out1 XOR Logical_Operator_out2164_out1;

  Logical_Operator_out3173_out1 <= Logical_Operator_out2133_out1 XOR Logical_Operator_out2165_out1;

  Logical_Operator_out3174_out1 <= Logical_Operator_out2134_out1 XOR Logical_Operator_out2166_out1;

  Logical_Operator_out3175_out1 <= Logical_Operator_out2135_out1 XOR Logical_Operator_out2167_out1;

  Logical_Operator_out3176_out1 <= Logical_Operator_out2136_out1 XOR Logical_Operator_out2168_out1;

  Logical_Operator_out3177_out1 <= Logical_Operator_out2137_out1 XOR Logical_Operator_out2169_out1;

  Logical_Operator_out3178_out1 <= Logical_Operator_out2138_out1 XOR Logical_Operator_out2170_out1;

  Logical_Operator_out3179_out1 <= Logical_Operator_out2139_out1 XOR Logical_Operator_out2171_out1;

  Logical_Operator_out3180_out1 <= Logical_Operator_out2140_out1 XOR Logical_Operator_out2172_out1;

  Logical_Operator_out3181_out1 <= Logical_Operator_out2141_out1 XOR Logical_Operator_out2173_out1;

  Logical_Operator_out3182_out1 <= Logical_Operator_out2142_out1 XOR Logical_Operator_out2174_out1;

  Logical_Operator_out3183_out1 <= Logical_Operator_out2143_out1 XOR Logical_Operator_out2175_out1;

  Logical_Operator_out3184_out1 <= Logical_Operator_out2144_out1 XOR Logical_Operator_out2176_out1;

  Logical_Operator_out3185_out1 <= Logical_Operator_out1625_out1 XOR Logical_Operator_out1657_out1;

  Logical_Operator_out3186_out1 <= Logical_Operator_out1626_out1 XOR Logical_Operator_out1658_out1;

  Logical_Operator_out3187_out1 <= Logical_Operator_out1627_out1 XOR Logical_Operator_out1659_out1;

  Logical_Operator_out3188_out1 <= Logical_Operator_out1628_out1 XOR Logical_Operator_out1660_out1;

  Logical_Operator_out3189_out1 <= Logical_Operator_out1629_out1 XOR Logical_Operator_out1661_out1;

  Logical_Operator_out3190_out1 <= Logical_Operator_out1630_out1 XOR Logical_Operator_out1662_out1;

  Logical_Operator_out3191_out1 <= Logical_Operator_out1631_out1 XOR Logical_Operator_out1663_out1;

  Logical_Operator_out3192_out1 <= Logical_Operator_out1632_out1 XOR Logical_Operator_out1664_out1;

  Logical_Operator_out3193_out1 <= Logical_Operator_out1117_out1 XOR Logical_Operator_out1149_out1;

  Logical_Operator_out3194_out1 <= Logical_Operator_out1118_out1 XOR Logical_Operator_out1150_out1;

  Logical_Operator_out3195_out1 <= Logical_Operator_out1119_out1 XOR Logical_Operator_out1151_out1;

  Logical_Operator_out3196_out1 <= Logical_Operator_out1120_out1 XOR Logical_Operator_out1152_out1;

  Logical_Operator_out3197_out1 <= Logical_Operator_out607_out1 XOR Logical_Operator_out639_out1;

  Logical_Operator_out3198_out1 <= Logical_Operator_out608_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out3199_out1 <= Logical_Operator_out96_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out3200_out1 <= in192 XOR in256;

  Logical_Operator_out3201_out1 <= Logical_Operator_out2689_out1 XOR Logical_Operator_out2721_out1;

  Logical_Operator_out3202_out1 <= Logical_Operator_out2690_out1 XOR Logical_Operator_out2722_out1;

  Logical_Operator_out3203_out1 <= Logical_Operator_out2691_out1 XOR Logical_Operator_out2723_out1;

  Logical_Operator_out3204_out1 <= Logical_Operator_out2692_out1 XOR Logical_Operator_out2724_out1;

  Logical_Operator_out3205_out1 <= Logical_Operator_out2693_out1 XOR Logical_Operator_out2725_out1;

  Logical_Operator_out3206_out1 <= Logical_Operator_out2694_out1 XOR Logical_Operator_out2726_out1;

  Logical_Operator_out3207_out1 <= Logical_Operator_out2695_out1 XOR Logical_Operator_out2727_out1;

  Logical_Operator_out3208_out1 <= Logical_Operator_out2696_out1 XOR Logical_Operator_out2728_out1;

  Logical_Operator_out3209_out1 <= Logical_Operator_out2697_out1 XOR Logical_Operator_out2729_out1;

  Logical_Operator_out3210_out1 <= Logical_Operator_out2698_out1 XOR Logical_Operator_out2730_out1;

  Logical_Operator_out3211_out1 <= Logical_Operator_out2699_out1 XOR Logical_Operator_out2731_out1;

  Logical_Operator_out3212_out1 <= Logical_Operator_out2700_out1 XOR Logical_Operator_out2732_out1;

  Logical_Operator_out3213_out1 <= Logical_Operator_out2701_out1 XOR Logical_Operator_out2733_out1;

  Logical_Operator_out3214_out1 <= Logical_Operator_out2702_out1 XOR Logical_Operator_out2734_out1;

  Logical_Operator_out3215_out1 <= Logical_Operator_out2703_out1 XOR Logical_Operator_out2735_out1;

  Logical_Operator_out3216_out1 <= Logical_Operator_out2704_out1 XOR Logical_Operator_out2736_out1;

  Logical_Operator_out3217_out1 <= Logical_Operator_out2705_out1 XOR Logical_Operator_out2737_out1;

  Logical_Operator_out3218_out1 <= Logical_Operator_out2706_out1 XOR Logical_Operator_out2738_out1;

  Logical_Operator_out3219_out1 <= Logical_Operator_out2707_out1 XOR Logical_Operator_out2739_out1;

  Logical_Operator_out3220_out1 <= Logical_Operator_out2708_out1 XOR Logical_Operator_out2740_out1;

  Logical_Operator_out3221_out1 <= Logical_Operator_out2709_out1 XOR Logical_Operator_out2741_out1;

  Logical_Operator_out3222_out1 <= Logical_Operator_out2710_out1 XOR Logical_Operator_out2742_out1;

  Logical_Operator_out3223_out1 <= Logical_Operator_out2711_out1 XOR Logical_Operator_out2743_out1;

  Logical_Operator_out3224_out1 <= Logical_Operator_out2712_out1 XOR Logical_Operator_out2744_out1;

  Logical_Operator_out3225_out1 <= Logical_Operator_out2713_out1 XOR Logical_Operator_out2745_out1;

  Logical_Operator_out3226_out1 <= Logical_Operator_out2714_out1 XOR Logical_Operator_out2746_out1;

  Logical_Operator_out3227_out1 <= Logical_Operator_out2715_out1 XOR Logical_Operator_out2747_out1;

  Logical_Operator_out3228_out1 <= Logical_Operator_out2716_out1 XOR Logical_Operator_out2748_out1;

  Logical_Operator_out3229_out1 <= Logical_Operator_out2717_out1 XOR Logical_Operator_out2749_out1;

  Logical_Operator_out3230_out1 <= Logical_Operator_out2718_out1 XOR Logical_Operator_out2750_out1;

  Logical_Operator_out3231_out1 <= Logical_Operator_out2719_out1 XOR Logical_Operator_out2751_out1;

  Logical_Operator_out3232_out1 <= Logical_Operator_out2720_out1 XOR Logical_Operator_out2752_out1;

  Logical_Operator_out3233_out1 <= Logical_Operator_out2193_out1 XOR Logical_Operator_out2225_out1;

  Logical_Operator_out3234_out1 <= Logical_Operator_out2194_out1 XOR Logical_Operator_out2226_out1;

  Logical_Operator_out3235_out1 <= Logical_Operator_out2195_out1 XOR Logical_Operator_out2227_out1;

  Logical_Operator_out3236_out1 <= Logical_Operator_out2196_out1 XOR Logical_Operator_out2228_out1;

  Logical_Operator_out3237_out1 <= Logical_Operator_out2197_out1 XOR Logical_Operator_out2229_out1;

  Logical_Operator_out3238_out1 <= Logical_Operator_out2198_out1 XOR Logical_Operator_out2230_out1;

  Logical_Operator_out3239_out1 <= Logical_Operator_out2199_out1 XOR Logical_Operator_out2231_out1;

  Logical_Operator_out3240_out1 <= Logical_Operator_out2200_out1 XOR Logical_Operator_out2232_out1;

  Logical_Operator_out3241_out1 <= Logical_Operator_out2201_out1 XOR Logical_Operator_out2233_out1;

  Logical_Operator_out3242_out1 <= Logical_Operator_out2202_out1 XOR Logical_Operator_out2234_out1;

  Logical_Operator_out3243_out1 <= Logical_Operator_out2203_out1 XOR Logical_Operator_out2235_out1;

  Logical_Operator_out3244_out1 <= Logical_Operator_out2204_out1 XOR Logical_Operator_out2236_out1;

  Logical_Operator_out3245_out1 <= Logical_Operator_out2205_out1 XOR Logical_Operator_out2237_out1;

  Logical_Operator_out3246_out1 <= Logical_Operator_out2206_out1 XOR Logical_Operator_out2238_out1;

  Logical_Operator_out3247_out1 <= Logical_Operator_out2207_out1 XOR Logical_Operator_out2239_out1;

  Logical_Operator_out3248_out1 <= Logical_Operator_out2208_out1 XOR Logical_Operator_out2240_out1;

  Logical_Operator_out3249_out1 <= Logical_Operator_out1689_out1 XOR Logical_Operator_out1721_out1;

  Logical_Operator_out3250_out1 <= Logical_Operator_out1690_out1 XOR Logical_Operator_out1722_out1;

  Logical_Operator_out3251_out1 <= Logical_Operator_out1691_out1 XOR Logical_Operator_out1723_out1;

  Logical_Operator_out3252_out1 <= Logical_Operator_out1692_out1 XOR Logical_Operator_out1724_out1;

  Logical_Operator_out3253_out1 <= Logical_Operator_out1693_out1 XOR Logical_Operator_out1725_out1;

  Logical_Operator_out3254_out1 <= Logical_Operator_out1694_out1 XOR Logical_Operator_out1726_out1;

  Logical_Operator_out3255_out1 <= Logical_Operator_out1695_out1 XOR Logical_Operator_out1727_out1;

  Logical_Operator_out3256_out1 <= Logical_Operator_out1696_out1 XOR Logical_Operator_out1728_out1;

  Logical_Operator_out3257_out1 <= Logical_Operator_out1181_out1 XOR Logical_Operator_out1213_out1;

  Logical_Operator_out3258_out1 <= Logical_Operator_out1182_out1 XOR Logical_Operator_out1214_out1;

  Logical_Operator_out3259_out1 <= Logical_Operator_out1183_out1 XOR Logical_Operator_out1215_out1;

  Logical_Operator_out3260_out1 <= Logical_Operator_out1184_out1 XOR Logical_Operator_out1216_out1;

  Logical_Operator_out3261_out1 <= Logical_Operator_out671_out1 XOR Logical_Operator_out703_out1;

  Logical_Operator_out3262_out1 <= Logical_Operator_out672_out1 XOR Logical_Operator_out704_out1;

  Logical_Operator_out3263_out1 <= Logical_Operator_out160_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out3264_out1 <= in320 XOR in384;

  Logical_Operator_out3265_out1 <= Logical_Operator_out2753_out1 XOR Logical_Operator_out2785_out1;

  Logical_Operator_out3266_out1 <= Logical_Operator_out2754_out1 XOR Logical_Operator_out2786_out1;

  Logical_Operator_out3267_out1 <= Logical_Operator_out2755_out1 XOR Logical_Operator_out2787_out1;

  Logical_Operator_out3268_out1 <= Logical_Operator_out2756_out1 XOR Logical_Operator_out2788_out1;

  Logical_Operator_out3269_out1 <= Logical_Operator_out2757_out1 XOR Logical_Operator_out2789_out1;

  Logical_Operator_out3270_out1 <= Logical_Operator_out2758_out1 XOR Logical_Operator_out2790_out1;

  Logical_Operator_out3271_out1 <= Logical_Operator_out2759_out1 XOR Logical_Operator_out2791_out1;

  Logical_Operator_out3272_out1 <= Logical_Operator_out2760_out1 XOR Logical_Operator_out2792_out1;

  Logical_Operator_out3273_out1 <= Logical_Operator_out2761_out1 XOR Logical_Operator_out2793_out1;

  Logical_Operator_out3274_out1 <= Logical_Operator_out2762_out1 XOR Logical_Operator_out2794_out1;

  Logical_Operator_out3275_out1 <= Logical_Operator_out2763_out1 XOR Logical_Operator_out2795_out1;

  Logical_Operator_out3276_out1 <= Logical_Operator_out2764_out1 XOR Logical_Operator_out2796_out1;

  Logical_Operator_out3277_out1 <= Logical_Operator_out2765_out1 XOR Logical_Operator_out2797_out1;

  Logical_Operator_out3278_out1 <= Logical_Operator_out2766_out1 XOR Logical_Operator_out2798_out1;

  Logical_Operator_out3279_out1 <= Logical_Operator_out2767_out1 XOR Logical_Operator_out2799_out1;

  Logical_Operator_out3280_out1 <= Logical_Operator_out2768_out1 XOR Logical_Operator_out2800_out1;

  Logical_Operator_out3281_out1 <= Logical_Operator_out2769_out1 XOR Logical_Operator_out2801_out1;

  Logical_Operator_out3282_out1 <= Logical_Operator_out2770_out1 XOR Logical_Operator_out2802_out1;

  Logical_Operator_out3283_out1 <= Logical_Operator_out2771_out1 XOR Logical_Operator_out2803_out1;

  Logical_Operator_out3284_out1 <= Logical_Operator_out2772_out1 XOR Logical_Operator_out2804_out1;

  Logical_Operator_out3285_out1 <= Logical_Operator_out2773_out1 XOR Logical_Operator_out2805_out1;

  Logical_Operator_out3286_out1 <= Logical_Operator_out2774_out1 XOR Logical_Operator_out2806_out1;

  Logical_Operator_out3287_out1 <= Logical_Operator_out2775_out1 XOR Logical_Operator_out2807_out1;

  Logical_Operator_out3288_out1 <= Logical_Operator_out2776_out1 XOR Logical_Operator_out2808_out1;

  Logical_Operator_out3289_out1 <= Logical_Operator_out2777_out1 XOR Logical_Operator_out2809_out1;

  Logical_Operator_out3290_out1 <= Logical_Operator_out2778_out1 XOR Logical_Operator_out2810_out1;

  Logical_Operator_out3291_out1 <= Logical_Operator_out2779_out1 XOR Logical_Operator_out2811_out1;

  Logical_Operator_out3292_out1 <= Logical_Operator_out2780_out1 XOR Logical_Operator_out2812_out1;

  Logical_Operator_out3293_out1 <= Logical_Operator_out2781_out1 XOR Logical_Operator_out2813_out1;

  Logical_Operator_out3294_out1 <= Logical_Operator_out2782_out1 XOR Logical_Operator_out2814_out1;

  Logical_Operator_out3295_out1 <= Logical_Operator_out2783_out1 XOR Logical_Operator_out2815_out1;

  Logical_Operator_out3296_out1 <= Logical_Operator_out2784_out1 XOR Logical_Operator_out2816_out1;

  Logical_Operator_out3297_out1 <= Logical_Operator_out2257_out1 XOR Logical_Operator_out2289_out1;

  Logical_Operator_out3298_out1 <= Logical_Operator_out2258_out1 XOR Logical_Operator_out2290_out1;

  Logical_Operator_out3299_out1 <= Logical_Operator_out2259_out1 XOR Logical_Operator_out2291_out1;

  Logical_Operator_out3300_out1 <= Logical_Operator_out2260_out1 XOR Logical_Operator_out2292_out1;

  Logical_Operator_out3301_out1 <= Logical_Operator_out2261_out1 XOR Logical_Operator_out2293_out1;

  Logical_Operator_out3302_out1 <= Logical_Operator_out2262_out1 XOR Logical_Operator_out2294_out1;

  Logical_Operator_out3303_out1 <= Logical_Operator_out2263_out1 XOR Logical_Operator_out2295_out1;

  Logical_Operator_out3304_out1 <= Logical_Operator_out2264_out1 XOR Logical_Operator_out2296_out1;

  Logical_Operator_out3305_out1 <= Logical_Operator_out2265_out1 XOR Logical_Operator_out2297_out1;

  Logical_Operator_out3306_out1 <= Logical_Operator_out2266_out1 XOR Logical_Operator_out2298_out1;

  Logical_Operator_out3307_out1 <= Logical_Operator_out2267_out1 XOR Logical_Operator_out2299_out1;

  Logical_Operator_out3308_out1 <= Logical_Operator_out2268_out1 XOR Logical_Operator_out2300_out1;

  Logical_Operator_out3309_out1 <= Logical_Operator_out2269_out1 XOR Logical_Operator_out2301_out1;

  Logical_Operator_out3310_out1 <= Logical_Operator_out2270_out1 XOR Logical_Operator_out2302_out1;

  Logical_Operator_out3311_out1 <= Logical_Operator_out2271_out1 XOR Logical_Operator_out2303_out1;

  Logical_Operator_out3312_out1 <= Logical_Operator_out2272_out1 XOR Logical_Operator_out2304_out1;

  Logical_Operator_out3313_out1 <= Logical_Operator_out1753_out1 XOR Logical_Operator_out1785_out1;

  Logical_Operator_out3314_out1 <= Logical_Operator_out1754_out1 XOR Logical_Operator_out1786_out1;

  Logical_Operator_out3315_out1 <= Logical_Operator_out1755_out1 XOR Logical_Operator_out1787_out1;

  Logical_Operator_out3316_out1 <= Logical_Operator_out1756_out1 XOR Logical_Operator_out1788_out1;

  Logical_Operator_out3317_out1 <= Logical_Operator_out1757_out1 XOR Logical_Operator_out1789_out1;

  Logical_Operator_out3318_out1 <= Logical_Operator_out1758_out1 XOR Logical_Operator_out1790_out1;

  Logical_Operator_out3319_out1 <= Logical_Operator_out1759_out1 XOR Logical_Operator_out1791_out1;

  Logical_Operator_out3320_out1 <= Logical_Operator_out1760_out1 XOR Logical_Operator_out1792_out1;

  Logical_Operator_out3321_out1 <= Logical_Operator_out1245_out1 XOR Logical_Operator_out1277_out1;

  Logical_Operator_out3322_out1 <= Logical_Operator_out1246_out1 XOR Logical_Operator_out1278_out1;

  Logical_Operator_out3323_out1 <= Logical_Operator_out1247_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out3324_out1 <= Logical_Operator_out1248_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out3325_out1 <= Logical_Operator_out735_out1 XOR Logical_Operator_out767_out1;

  Logical_Operator_out3326_out1 <= Logical_Operator_out736_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out3327_out1 <= Logical_Operator_out224_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out3328_out1 <= in448 XOR in512;

  Logical_Operator_out3329_out1 <= Logical_Operator_out2817_out1 XOR Logical_Operator_out2849_out1;

  Logical_Operator_out3330_out1 <= Logical_Operator_out2818_out1 XOR Logical_Operator_out2850_out1;

  Logical_Operator_out3331_out1 <= Logical_Operator_out2819_out1 XOR Logical_Operator_out2851_out1;

  Logical_Operator_out3332_out1 <= Logical_Operator_out2820_out1 XOR Logical_Operator_out2852_out1;

  Logical_Operator_out3333_out1 <= Logical_Operator_out2821_out1 XOR Logical_Operator_out2853_out1;

  Logical_Operator_out3334_out1 <= Logical_Operator_out2822_out1 XOR Logical_Operator_out2854_out1;

  Logical_Operator_out3335_out1 <= Logical_Operator_out2823_out1 XOR Logical_Operator_out2855_out1;

  Logical_Operator_out3336_out1 <= Logical_Operator_out2824_out1 XOR Logical_Operator_out2856_out1;

  Logical_Operator_out3337_out1 <= Logical_Operator_out2825_out1 XOR Logical_Operator_out2857_out1;

  Logical_Operator_out3338_out1 <= Logical_Operator_out2826_out1 XOR Logical_Operator_out2858_out1;

  Logical_Operator_out3339_out1 <= Logical_Operator_out2827_out1 XOR Logical_Operator_out2859_out1;

  Logical_Operator_out3340_out1 <= Logical_Operator_out2828_out1 XOR Logical_Operator_out2860_out1;

  Logical_Operator_out3341_out1 <= Logical_Operator_out2829_out1 XOR Logical_Operator_out2861_out1;

  Logical_Operator_out3342_out1 <= Logical_Operator_out2830_out1 XOR Logical_Operator_out2862_out1;

  Logical_Operator_out3343_out1 <= Logical_Operator_out2831_out1 XOR Logical_Operator_out2863_out1;

  Logical_Operator_out3344_out1 <= Logical_Operator_out2832_out1 XOR Logical_Operator_out2864_out1;

  Logical_Operator_out3345_out1 <= Logical_Operator_out2833_out1 XOR Logical_Operator_out2865_out1;

  Logical_Operator_out3346_out1 <= Logical_Operator_out2834_out1 XOR Logical_Operator_out2866_out1;

  Logical_Operator_out3347_out1 <= Logical_Operator_out2835_out1 XOR Logical_Operator_out2867_out1;

  Logical_Operator_out3348_out1 <= Logical_Operator_out2836_out1 XOR Logical_Operator_out2868_out1;

  Logical_Operator_out3349_out1 <= Logical_Operator_out2837_out1 XOR Logical_Operator_out2869_out1;

  Logical_Operator_out3350_out1 <= Logical_Operator_out2838_out1 XOR Logical_Operator_out2870_out1;

  Logical_Operator_out3351_out1 <= Logical_Operator_out2839_out1 XOR Logical_Operator_out2871_out1;

  Logical_Operator_out3352_out1 <= Logical_Operator_out2840_out1 XOR Logical_Operator_out2872_out1;

  Logical_Operator_out3353_out1 <= Logical_Operator_out2841_out1 XOR Logical_Operator_out2873_out1;

  Logical_Operator_out3354_out1 <= Logical_Operator_out2842_out1 XOR Logical_Operator_out2874_out1;

  Logical_Operator_out3355_out1 <= Logical_Operator_out2843_out1 XOR Logical_Operator_out2875_out1;

  Logical_Operator_out3356_out1 <= Logical_Operator_out2844_out1 XOR Logical_Operator_out2876_out1;

  Logical_Operator_out3357_out1 <= Logical_Operator_out2845_out1 XOR Logical_Operator_out2877_out1;

  Logical_Operator_out3358_out1 <= Logical_Operator_out2846_out1 XOR Logical_Operator_out2878_out1;

  Logical_Operator_out3359_out1 <= Logical_Operator_out2847_out1 XOR Logical_Operator_out2879_out1;

  Logical_Operator_out3360_out1 <= Logical_Operator_out2848_out1 XOR Logical_Operator_out2880_out1;

  Logical_Operator_out3361_out1 <= Logical_Operator_out2321_out1 XOR Logical_Operator_out2353_out1;

  Logical_Operator_out3362_out1 <= Logical_Operator_out2322_out1 XOR Logical_Operator_out2354_out1;

  Logical_Operator_out3363_out1 <= Logical_Operator_out2323_out1 XOR Logical_Operator_out2355_out1;

  Logical_Operator_out3364_out1 <= Logical_Operator_out2324_out1 XOR Logical_Operator_out2356_out1;

  Logical_Operator_out3365_out1 <= Logical_Operator_out2325_out1 XOR Logical_Operator_out2357_out1;

  Logical_Operator_out3366_out1 <= Logical_Operator_out2326_out1 XOR Logical_Operator_out2358_out1;

  Logical_Operator_out3367_out1 <= Logical_Operator_out2327_out1 XOR Logical_Operator_out2359_out1;

  Logical_Operator_out3368_out1 <= Logical_Operator_out2328_out1 XOR Logical_Operator_out2360_out1;

  Logical_Operator_out3369_out1 <= Logical_Operator_out2329_out1 XOR Logical_Operator_out2361_out1;

  Logical_Operator_out3370_out1 <= Logical_Operator_out2330_out1 XOR Logical_Operator_out2362_out1;

  Logical_Operator_out3371_out1 <= Logical_Operator_out2331_out1 XOR Logical_Operator_out2363_out1;

  Logical_Operator_out3372_out1 <= Logical_Operator_out2332_out1 XOR Logical_Operator_out2364_out1;

  Logical_Operator_out3373_out1 <= Logical_Operator_out2333_out1 XOR Logical_Operator_out2365_out1;

  Logical_Operator_out3374_out1 <= Logical_Operator_out2334_out1 XOR Logical_Operator_out2366_out1;

  Logical_Operator_out3375_out1 <= Logical_Operator_out2335_out1 XOR Logical_Operator_out2367_out1;

  Logical_Operator_out3376_out1 <= Logical_Operator_out2336_out1 XOR Logical_Operator_out2368_out1;

  Logical_Operator_out3377_out1 <= Logical_Operator_out1817_out1 XOR Logical_Operator_out1849_out1;

  Logical_Operator_out3378_out1 <= Logical_Operator_out1818_out1 XOR Logical_Operator_out1850_out1;

  Logical_Operator_out3379_out1 <= Logical_Operator_out1819_out1 XOR Logical_Operator_out1851_out1;

  Logical_Operator_out3380_out1 <= Logical_Operator_out1820_out1 XOR Logical_Operator_out1852_out1;

  Logical_Operator_out3381_out1 <= Logical_Operator_out1821_out1 XOR Logical_Operator_out1853_out1;

  Logical_Operator_out3382_out1 <= Logical_Operator_out1822_out1 XOR Logical_Operator_out1854_out1;

  Logical_Operator_out3383_out1 <= Logical_Operator_out1823_out1 XOR Logical_Operator_out1855_out1;

  Logical_Operator_out3384_out1 <= Logical_Operator_out1824_out1 XOR Logical_Operator_out1856_out1;

  Logical_Operator_out3385_out1 <= Logical_Operator_out1309_out1 XOR Logical_Operator_out1341_out1;

  Logical_Operator_out3386_out1 <= Logical_Operator_out1310_out1 XOR Logical_Operator_out1342_out1;

  Logical_Operator_out3387_out1 <= Logical_Operator_out1311_out1 XOR Logical_Operator_out1343_out1;

  Logical_Operator_out3388_out1 <= Logical_Operator_out1312_out1 XOR Logical_Operator_out1344_out1;

  Logical_Operator_out3389_out1 <= Logical_Operator_out799_out1 XOR Logical_Operator_out831_out1;

  Logical_Operator_out3390_out1 <= Logical_Operator_out800_out1 XOR Logical_Operator_out832_out1;

  Logical_Operator_out3391_out1 <= Logical_Operator_out288_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out3392_out1 <= in576 XOR in640;

  Logical_Operator_out3393_out1 <= Logical_Operator_out2881_out1 XOR Logical_Operator_out2913_out1;

  Logical_Operator_out3394_out1 <= Logical_Operator_out2882_out1 XOR Logical_Operator_out2914_out1;

  Logical_Operator_out3395_out1 <= Logical_Operator_out2883_out1 XOR Logical_Operator_out2915_out1;

  Logical_Operator_out3396_out1 <= Logical_Operator_out2884_out1 XOR Logical_Operator_out2916_out1;

  Logical_Operator_out3397_out1 <= Logical_Operator_out2885_out1 XOR Logical_Operator_out2917_out1;

  Logical_Operator_out3398_out1 <= Logical_Operator_out2886_out1 XOR Logical_Operator_out2918_out1;

  Logical_Operator_out3399_out1 <= Logical_Operator_out2887_out1 XOR Logical_Operator_out2919_out1;

  Logical_Operator_out3400_out1 <= Logical_Operator_out2888_out1 XOR Logical_Operator_out2920_out1;

  Logical_Operator_out3401_out1 <= Logical_Operator_out2889_out1 XOR Logical_Operator_out2921_out1;

  Logical_Operator_out3402_out1 <= Logical_Operator_out2890_out1 XOR Logical_Operator_out2922_out1;

  Logical_Operator_out3403_out1 <= Logical_Operator_out2891_out1 XOR Logical_Operator_out2923_out1;

  Logical_Operator_out3404_out1 <= Logical_Operator_out2892_out1 XOR Logical_Operator_out2924_out1;

  Logical_Operator_out3405_out1 <= Logical_Operator_out2893_out1 XOR Logical_Operator_out2925_out1;

  Logical_Operator_out3406_out1 <= Logical_Operator_out2894_out1 XOR Logical_Operator_out2926_out1;

  Logical_Operator_out3407_out1 <= Logical_Operator_out2895_out1 XOR Logical_Operator_out2927_out1;

  Logical_Operator_out3408_out1 <= Logical_Operator_out2896_out1 XOR Logical_Operator_out2928_out1;

  Logical_Operator_out3409_out1 <= Logical_Operator_out2897_out1 XOR Logical_Operator_out2929_out1;

  Logical_Operator_out3410_out1 <= Logical_Operator_out2898_out1 XOR Logical_Operator_out2930_out1;

  Logical_Operator_out3411_out1 <= Logical_Operator_out2899_out1 XOR Logical_Operator_out2931_out1;

  Logical_Operator_out3412_out1 <= Logical_Operator_out2900_out1 XOR Logical_Operator_out2932_out1;

  Logical_Operator_out3413_out1 <= Logical_Operator_out2901_out1 XOR Logical_Operator_out2933_out1;

  Logical_Operator_out3414_out1 <= Logical_Operator_out2902_out1 XOR Logical_Operator_out2934_out1;

  Logical_Operator_out3415_out1 <= Logical_Operator_out2903_out1 XOR Logical_Operator_out2935_out1;

  Logical_Operator_out3416_out1 <= Logical_Operator_out2904_out1 XOR Logical_Operator_out2936_out1;

  Logical_Operator_out3417_out1 <= Logical_Operator_out2905_out1 XOR Logical_Operator_out2937_out1;

  Logical_Operator_out3418_out1 <= Logical_Operator_out2906_out1 XOR Logical_Operator_out2938_out1;

  Logical_Operator_out3419_out1 <= Logical_Operator_out2907_out1 XOR Logical_Operator_out2939_out1;

  Logical_Operator_out3420_out1 <= Logical_Operator_out2908_out1 XOR Logical_Operator_out2940_out1;

  Logical_Operator_out3421_out1 <= Logical_Operator_out2909_out1 XOR Logical_Operator_out2941_out1;

  Logical_Operator_out3422_out1 <= Logical_Operator_out2910_out1 XOR Logical_Operator_out2942_out1;

  Logical_Operator_out3423_out1 <= Logical_Operator_out2911_out1 XOR Logical_Operator_out2943_out1;

  Logical_Operator_out3424_out1 <= Logical_Operator_out2912_out1 XOR Logical_Operator_out2944_out1;

  Logical_Operator_out3425_out1 <= Logical_Operator_out2385_out1 XOR Logical_Operator_out2417_out1;

  Logical_Operator_out3426_out1 <= Logical_Operator_out2386_out1 XOR Logical_Operator_out2418_out1;

  Logical_Operator_out3427_out1 <= Logical_Operator_out2387_out1 XOR Logical_Operator_out2419_out1;

  Logical_Operator_out3428_out1 <= Logical_Operator_out2388_out1 XOR Logical_Operator_out2420_out1;

  Logical_Operator_out3429_out1 <= Logical_Operator_out2389_out1 XOR Logical_Operator_out2421_out1;

  Logical_Operator_out3430_out1 <= Logical_Operator_out2390_out1 XOR Logical_Operator_out2422_out1;

  Logical_Operator_out3431_out1 <= Logical_Operator_out2391_out1 XOR Logical_Operator_out2423_out1;

  Logical_Operator_out3432_out1 <= Logical_Operator_out2392_out1 XOR Logical_Operator_out2424_out1;

  Logical_Operator_out3433_out1 <= Logical_Operator_out2393_out1 XOR Logical_Operator_out2425_out1;

  Logical_Operator_out3434_out1 <= Logical_Operator_out2394_out1 XOR Logical_Operator_out2426_out1;

  Logical_Operator_out3435_out1 <= Logical_Operator_out2395_out1 XOR Logical_Operator_out2427_out1;

  Logical_Operator_out3436_out1 <= Logical_Operator_out2396_out1 XOR Logical_Operator_out2428_out1;

  Logical_Operator_out3437_out1 <= Logical_Operator_out2397_out1 XOR Logical_Operator_out2429_out1;

  Logical_Operator_out3438_out1 <= Logical_Operator_out2398_out1 XOR Logical_Operator_out2430_out1;

  Logical_Operator_out3439_out1 <= Logical_Operator_out2399_out1 XOR Logical_Operator_out2431_out1;

  Logical_Operator_out3440_out1 <= Logical_Operator_out2400_out1 XOR Logical_Operator_out2432_out1;

  Logical_Operator_out3441_out1 <= Logical_Operator_out1881_out1 XOR Logical_Operator_out1913_out1;

  Logical_Operator_out3442_out1 <= Logical_Operator_out1882_out1 XOR Logical_Operator_out1914_out1;

  Logical_Operator_out3443_out1 <= Logical_Operator_out1883_out1 XOR Logical_Operator_out1915_out1;

  Logical_Operator_out3444_out1 <= Logical_Operator_out1884_out1 XOR Logical_Operator_out1916_out1;

  Logical_Operator_out3445_out1 <= Logical_Operator_out1885_out1 XOR Logical_Operator_out1917_out1;

  Logical_Operator_out3446_out1 <= Logical_Operator_out1886_out1 XOR Logical_Operator_out1918_out1;

  Logical_Operator_out3447_out1 <= Logical_Operator_out1887_out1 XOR Logical_Operator_out1919_out1;

  Logical_Operator_out3448_out1 <= Logical_Operator_out1888_out1 XOR Logical_Operator_out1920_out1;

  Logical_Operator_out3449_out1 <= Logical_Operator_out1373_out1 XOR Logical_Operator_out1405_out1;

  Logical_Operator_out3450_out1 <= Logical_Operator_out1374_out1 XOR Logical_Operator_out1406_out1;

  Logical_Operator_out3451_out1 <= Logical_Operator_out1375_out1 XOR Logical_Operator_out1407_out1;

  Logical_Operator_out3452_out1 <= Logical_Operator_out1376_out1 XOR Logical_Operator_out1408_out1;

  Logical_Operator_out3453_out1 <= Logical_Operator_out863_out1 XOR Logical_Operator_out895_out1;

  Logical_Operator_out3454_out1 <= Logical_Operator_out864_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out3455_out1 <= Logical_Operator_out352_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out3456_out1 <= in704 XOR in768;

  Logical_Operator_out3457_out1 <= Logical_Operator_out2945_out1 XOR Logical_Operator_out2977_out1;

  Logical_Operator_out3458_out1 <= Logical_Operator_out2946_out1 XOR Logical_Operator_out2978_out1;

  Logical_Operator_out3459_out1 <= Logical_Operator_out2947_out1 XOR Logical_Operator_out2979_out1;

  Logical_Operator_out3460_out1 <= Logical_Operator_out2948_out1 XOR Logical_Operator_out2980_out1;

  Logical_Operator_out3461_out1 <= Logical_Operator_out2949_out1 XOR Logical_Operator_out2981_out1;

  Logical_Operator_out3462_out1 <= Logical_Operator_out2950_out1 XOR Logical_Operator_out2982_out1;

  Logical_Operator_out3463_out1 <= Logical_Operator_out2951_out1 XOR Logical_Operator_out2983_out1;

  Logical_Operator_out3464_out1 <= Logical_Operator_out2952_out1 XOR Logical_Operator_out2984_out1;

  Logical_Operator_out3465_out1 <= Logical_Operator_out2953_out1 XOR Logical_Operator_out2985_out1;

  Logical_Operator_out3466_out1 <= Logical_Operator_out2954_out1 XOR Logical_Operator_out2986_out1;

  Logical_Operator_out3467_out1 <= Logical_Operator_out2955_out1 XOR Logical_Operator_out2987_out1;

  Logical_Operator_out3468_out1 <= Logical_Operator_out2956_out1 XOR Logical_Operator_out2988_out1;

  Logical_Operator_out3469_out1 <= Logical_Operator_out2957_out1 XOR Logical_Operator_out2989_out1;

  Logical_Operator_out3470_out1 <= Logical_Operator_out2958_out1 XOR Logical_Operator_out2990_out1;

  Logical_Operator_out3471_out1 <= Logical_Operator_out2959_out1 XOR Logical_Operator_out2991_out1;

  Logical_Operator_out3472_out1 <= Logical_Operator_out2960_out1 XOR Logical_Operator_out2992_out1;

  Logical_Operator_out3473_out1 <= Logical_Operator_out2961_out1 XOR Logical_Operator_out2993_out1;

  Logical_Operator_out3474_out1 <= Logical_Operator_out2962_out1 XOR Logical_Operator_out2994_out1;

  Logical_Operator_out3475_out1 <= Logical_Operator_out2963_out1 XOR Logical_Operator_out2995_out1;

  Logical_Operator_out3476_out1 <= Logical_Operator_out2964_out1 XOR Logical_Operator_out2996_out1;

  Logical_Operator_out3477_out1 <= Logical_Operator_out2965_out1 XOR Logical_Operator_out2997_out1;

  Logical_Operator_out3478_out1 <= Logical_Operator_out2966_out1 XOR Logical_Operator_out2998_out1;

  Logical_Operator_out3479_out1 <= Logical_Operator_out2967_out1 XOR Logical_Operator_out2999_out1;

  Logical_Operator_out3480_out1 <= Logical_Operator_out2968_out1 XOR Logical_Operator_out3000_out1;

  Logical_Operator_out3481_out1 <= Logical_Operator_out2969_out1 XOR Logical_Operator_out3001_out1;

  Logical_Operator_out3482_out1 <= Logical_Operator_out2970_out1 XOR Logical_Operator_out3002_out1;

  Logical_Operator_out3483_out1 <= Logical_Operator_out2971_out1 XOR Logical_Operator_out3003_out1;

  Logical_Operator_out3484_out1 <= Logical_Operator_out2972_out1 XOR Logical_Operator_out3004_out1;

  Logical_Operator_out3485_out1 <= Logical_Operator_out2973_out1 XOR Logical_Operator_out3005_out1;

  Logical_Operator_out3486_out1 <= Logical_Operator_out2974_out1 XOR Logical_Operator_out3006_out1;

  Logical_Operator_out3487_out1 <= Logical_Operator_out2975_out1 XOR Logical_Operator_out3007_out1;

  Logical_Operator_out3488_out1 <= Logical_Operator_out2976_out1 XOR Logical_Operator_out3008_out1;

  Logical_Operator_out3489_out1 <= Logical_Operator_out2449_out1 XOR Logical_Operator_out2481_out1;

  Logical_Operator_out3490_out1 <= Logical_Operator_out2450_out1 XOR Logical_Operator_out2482_out1;

  Logical_Operator_out3491_out1 <= Logical_Operator_out2451_out1 XOR Logical_Operator_out2483_out1;

  Logical_Operator_out3492_out1 <= Logical_Operator_out2452_out1 XOR Logical_Operator_out2484_out1;

  Logical_Operator_out3493_out1 <= Logical_Operator_out2453_out1 XOR Logical_Operator_out2485_out1;

  Logical_Operator_out3494_out1 <= Logical_Operator_out2454_out1 XOR Logical_Operator_out2486_out1;

  Logical_Operator_out3495_out1 <= Logical_Operator_out2455_out1 XOR Logical_Operator_out2487_out1;

  Logical_Operator_out3496_out1 <= Logical_Operator_out2456_out1 XOR Logical_Operator_out2488_out1;

  Logical_Operator_out3497_out1 <= Logical_Operator_out2457_out1 XOR Logical_Operator_out2489_out1;

  Logical_Operator_out3498_out1 <= Logical_Operator_out2458_out1 XOR Logical_Operator_out2490_out1;

  Logical_Operator_out3499_out1 <= Logical_Operator_out2459_out1 XOR Logical_Operator_out2491_out1;

  Logical_Operator_out3500_out1 <= Logical_Operator_out2460_out1 XOR Logical_Operator_out2492_out1;

  Logical_Operator_out3501_out1 <= Logical_Operator_out2461_out1 XOR Logical_Operator_out2493_out1;

  Logical_Operator_out3502_out1 <= Logical_Operator_out2462_out1 XOR Logical_Operator_out2494_out1;

  Logical_Operator_out3503_out1 <= Logical_Operator_out2463_out1 XOR Logical_Operator_out2495_out1;

  Logical_Operator_out3504_out1 <= Logical_Operator_out2464_out1 XOR Logical_Operator_out2496_out1;

  Logical_Operator_out3505_out1 <= Logical_Operator_out1945_out1 XOR Logical_Operator_out1977_out1;

  Logical_Operator_out3506_out1 <= Logical_Operator_out1946_out1 XOR Logical_Operator_out1978_out1;

  Logical_Operator_out3507_out1 <= Logical_Operator_out1947_out1 XOR Logical_Operator_out1979_out1;

  Logical_Operator_out3508_out1 <= Logical_Operator_out1948_out1 XOR Logical_Operator_out1980_out1;

  Logical_Operator_out3509_out1 <= Logical_Operator_out1949_out1 XOR Logical_Operator_out1981_out1;

  Logical_Operator_out3510_out1 <= Logical_Operator_out1950_out1 XOR Logical_Operator_out1982_out1;

  Logical_Operator_out3511_out1 <= Logical_Operator_out1951_out1 XOR Logical_Operator_out1983_out1;

  Logical_Operator_out3512_out1 <= Logical_Operator_out1952_out1 XOR Logical_Operator_out1984_out1;

  Logical_Operator_out3513_out1 <= Logical_Operator_out1437_out1 XOR Logical_Operator_out1469_out1;

  Logical_Operator_out3514_out1 <= Logical_Operator_out1438_out1 XOR Logical_Operator_out1470_out1;

  Logical_Operator_out3515_out1 <= Logical_Operator_out1439_out1 XOR Logical_Operator_out1471_out1;

  Logical_Operator_out3516_out1 <= Logical_Operator_out1440_out1 XOR Logical_Operator_out1472_out1;

  Logical_Operator_out3517_out1 <= Logical_Operator_out927_out1 XOR Logical_Operator_out959_out1;

  Logical_Operator_out3518_out1 <= Logical_Operator_out928_out1 XOR Logical_Operator_out960_out1;

  Logical_Operator_out3519_out1 <= Logical_Operator_out416_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out3520_out1 <= in832 XOR in896;

  Logical_Operator_out3521_out1 <= Logical_Operator_out3009_out1 XOR Logical_Operator_out3041_out1;

  Logical_Operator_out3522_out1 <= Logical_Operator_out3010_out1 XOR Logical_Operator_out3042_out1;

  Logical_Operator_out3523_out1 <= Logical_Operator_out3011_out1 XOR Logical_Operator_out3043_out1;

  Logical_Operator_out3524_out1 <= Logical_Operator_out3012_out1 XOR Logical_Operator_out3044_out1;

  Logical_Operator_out3525_out1 <= Logical_Operator_out3013_out1 XOR Logical_Operator_out3045_out1;

  Logical_Operator_out3526_out1 <= Logical_Operator_out3014_out1 XOR Logical_Operator_out3046_out1;

  Logical_Operator_out3527_out1 <= Logical_Operator_out3015_out1 XOR Logical_Operator_out3047_out1;

  Logical_Operator_out3528_out1 <= Logical_Operator_out3016_out1 XOR Logical_Operator_out3048_out1;

  Logical_Operator_out3529_out1 <= Logical_Operator_out3017_out1 XOR Logical_Operator_out3049_out1;

  Logical_Operator_out3530_out1 <= Logical_Operator_out3018_out1 XOR Logical_Operator_out3050_out1;

  Logical_Operator_out3531_out1 <= Logical_Operator_out3019_out1 XOR Logical_Operator_out3051_out1;

  Logical_Operator_out3532_out1 <= Logical_Operator_out3020_out1 XOR Logical_Operator_out3052_out1;

  Logical_Operator_out3533_out1 <= Logical_Operator_out3021_out1 XOR Logical_Operator_out3053_out1;

  Logical_Operator_out3534_out1 <= Logical_Operator_out3022_out1 XOR Logical_Operator_out3054_out1;

  Logical_Operator_out3535_out1 <= Logical_Operator_out3023_out1 XOR Logical_Operator_out3055_out1;

  Logical_Operator_out3536_out1 <= Logical_Operator_out3024_out1 XOR Logical_Operator_out3056_out1;

  Logical_Operator_out3537_out1 <= Logical_Operator_out3025_out1 XOR Logical_Operator_out3057_out1;

  Logical_Operator_out3538_out1 <= Logical_Operator_out3026_out1 XOR Logical_Operator_out3058_out1;

  Logical_Operator_out3539_out1 <= Logical_Operator_out3027_out1 XOR Logical_Operator_out3059_out1;

  Logical_Operator_out3540_out1 <= Logical_Operator_out3028_out1 XOR Logical_Operator_out3060_out1;

  Logical_Operator_out3541_out1 <= Logical_Operator_out3029_out1 XOR Logical_Operator_out3061_out1;

  Logical_Operator_out3542_out1 <= Logical_Operator_out3030_out1 XOR Logical_Operator_out3062_out1;

  Logical_Operator_out3543_out1 <= Logical_Operator_out3031_out1 XOR Logical_Operator_out3063_out1;

  Logical_Operator_out3544_out1 <= Logical_Operator_out3032_out1 XOR Logical_Operator_out3064_out1;

  Logical_Operator_out3545_out1 <= Logical_Operator_out3033_out1 XOR Logical_Operator_out3065_out1;

  Logical_Operator_out3546_out1 <= Logical_Operator_out3034_out1 XOR Logical_Operator_out3066_out1;

  Logical_Operator_out3547_out1 <= Logical_Operator_out3035_out1 XOR Logical_Operator_out3067_out1;

  Logical_Operator_out3548_out1 <= Logical_Operator_out3036_out1 XOR Logical_Operator_out3068_out1;

  Logical_Operator_out3549_out1 <= Logical_Operator_out3037_out1 XOR Logical_Operator_out3069_out1;

  Logical_Operator_out3550_out1 <= Logical_Operator_out3038_out1 XOR Logical_Operator_out3070_out1;

  Logical_Operator_out3551_out1 <= Logical_Operator_out3039_out1 XOR Logical_Operator_out3071_out1;

  Logical_Operator_out3552_out1 <= Logical_Operator_out3040_out1 XOR Logical_Operator_out3072_out1;

  Logical_Operator_out3553_out1 <= Logical_Operator_out2513_out1 XOR Logical_Operator_out2545_out1;

  Logical_Operator_out3554_out1 <= Logical_Operator_out2514_out1 XOR Logical_Operator_out2546_out1;

  Logical_Operator_out3555_out1 <= Logical_Operator_out2515_out1 XOR Logical_Operator_out2547_out1;

  Logical_Operator_out3556_out1 <= Logical_Operator_out2516_out1 XOR Logical_Operator_out2548_out1;

  Logical_Operator_out3557_out1 <= Logical_Operator_out2517_out1 XOR Logical_Operator_out2549_out1;

  Logical_Operator_out3558_out1 <= Logical_Operator_out2518_out1 XOR Logical_Operator_out2550_out1;

  Logical_Operator_out3559_out1 <= Logical_Operator_out2519_out1 XOR Logical_Operator_out2551_out1;

  Logical_Operator_out3560_out1 <= Logical_Operator_out2520_out1 XOR Logical_Operator_out2552_out1;

  Logical_Operator_out3561_out1 <= Logical_Operator_out2521_out1 XOR Logical_Operator_out2553_out1;

  Logical_Operator_out3562_out1 <= Logical_Operator_out2522_out1 XOR Logical_Operator_out2554_out1;

  Logical_Operator_out3563_out1 <= Logical_Operator_out2523_out1 XOR Logical_Operator_out2555_out1;

  Logical_Operator_out3564_out1 <= Logical_Operator_out2524_out1 XOR Logical_Operator_out2556_out1;

  Logical_Operator_out3565_out1 <= Logical_Operator_out2525_out1 XOR Logical_Operator_out2557_out1;

  Logical_Operator_out3566_out1 <= Logical_Operator_out2526_out1 XOR Logical_Operator_out2558_out1;

  Logical_Operator_out3567_out1 <= Logical_Operator_out2527_out1 XOR Logical_Operator_out2559_out1;

  Logical_Operator_out3568_out1 <= Logical_Operator_out2528_out1 XOR Logical_Operator_out2560_out1;

  Logical_Operator_out3569_out1 <= Logical_Operator_out2009_out1 XOR Logical_Operator_out2041_out1;

  Logical_Operator_out3570_out1 <= Logical_Operator_out2010_out1 XOR Logical_Operator_out2042_out1;

  Logical_Operator_out3571_out1 <= Logical_Operator_out2011_out1 XOR Logical_Operator_out2043_out1;

  Logical_Operator_out3572_out1 <= Logical_Operator_out2012_out1 XOR Logical_Operator_out2044_out1;

  Logical_Operator_out3573_out1 <= Logical_Operator_out2013_out1 XOR Logical_Operator_out2045_out1;

  Logical_Operator_out3574_out1 <= Logical_Operator_out2014_out1 XOR Logical_Operator_out2046_out1;

  Logical_Operator_out3575_out1 <= Logical_Operator_out2015_out1 XOR Logical_Operator_out2047_out1;

  Logical_Operator_out3576_out1 <= Logical_Operator_out2016_out1 XOR Logical_Operator_out2048_out1;

  Logical_Operator_out3577_out1 <= Logical_Operator_out1501_out1 XOR Logical_Operator_out1533_out1;

  Logical_Operator_out3578_out1 <= Logical_Operator_out1502_out1 XOR Logical_Operator_out1534_out1;

  Logical_Operator_out3579_out1 <= Logical_Operator_out1503_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out3580_out1 <= Logical_Operator_out1504_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out3581_out1 <= Logical_Operator_out991_out1 XOR Logical_Operator_out1023_out1;

  Logical_Operator_out3582_out1 <= Logical_Operator_out992_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out3583_out1 <= Logical_Operator_out480_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out3584_out1 <= in960 XOR in1024;

  Logical_Operator_out3585_out1 <= Logical_Operator_out3073_out1 XOR Logical_Operator_out3137_out1;

  Logical_Operator_out3586_out1 <= Logical_Operator_out3074_out1 XOR Logical_Operator_out3138_out1;

  Logical_Operator_out3587_out1 <= Logical_Operator_out3075_out1 XOR Logical_Operator_out3139_out1;

  Logical_Operator_out3588_out1 <= Logical_Operator_out3076_out1 XOR Logical_Operator_out3140_out1;

  Logical_Operator_out3589_out1 <= Logical_Operator_out3077_out1 XOR Logical_Operator_out3141_out1;

  Logical_Operator_out3590_out1 <= Logical_Operator_out3078_out1 XOR Logical_Operator_out3142_out1;

  Logical_Operator_out3591_out1 <= Logical_Operator_out3079_out1 XOR Logical_Operator_out3143_out1;

  Logical_Operator_out3592_out1 <= Logical_Operator_out3080_out1 XOR Logical_Operator_out3144_out1;

  Logical_Operator_out3593_out1 <= Logical_Operator_out3081_out1 XOR Logical_Operator_out3145_out1;

  Logical_Operator_out3594_out1 <= Logical_Operator_out3082_out1 XOR Logical_Operator_out3146_out1;

  Logical_Operator_out3595_out1 <= Logical_Operator_out3083_out1 XOR Logical_Operator_out3147_out1;

  Logical_Operator_out3596_out1 <= Logical_Operator_out3084_out1 XOR Logical_Operator_out3148_out1;

  Logical_Operator_out3597_out1 <= Logical_Operator_out3085_out1 XOR Logical_Operator_out3149_out1;

  Logical_Operator_out3598_out1 <= Logical_Operator_out3086_out1 XOR Logical_Operator_out3150_out1;

  Logical_Operator_out3599_out1 <= Logical_Operator_out3087_out1 XOR Logical_Operator_out3151_out1;

  Logical_Operator_out3600_out1 <= Logical_Operator_out3088_out1 XOR Logical_Operator_out3152_out1;

  Logical_Operator_out3601_out1 <= Logical_Operator_out3089_out1 XOR Logical_Operator_out3153_out1;

  Logical_Operator_out3602_out1 <= Logical_Operator_out3090_out1 XOR Logical_Operator_out3154_out1;

  Logical_Operator_out3603_out1 <= Logical_Operator_out3091_out1 XOR Logical_Operator_out3155_out1;

  Logical_Operator_out3604_out1 <= Logical_Operator_out3092_out1 XOR Logical_Operator_out3156_out1;

  Logical_Operator_out3605_out1 <= Logical_Operator_out3093_out1 XOR Logical_Operator_out3157_out1;

  Logical_Operator_out3606_out1 <= Logical_Operator_out3094_out1 XOR Logical_Operator_out3158_out1;

  Logical_Operator_out3607_out1 <= Logical_Operator_out3095_out1 XOR Logical_Operator_out3159_out1;

  Logical_Operator_out3608_out1 <= Logical_Operator_out3096_out1 XOR Logical_Operator_out3160_out1;

  Logical_Operator_out3609_out1 <= Logical_Operator_out3097_out1 XOR Logical_Operator_out3161_out1;

  Logical_Operator_out3610_out1 <= Logical_Operator_out3098_out1 XOR Logical_Operator_out3162_out1;

  Logical_Operator_out3611_out1 <= Logical_Operator_out3099_out1 XOR Logical_Operator_out3163_out1;

  Logical_Operator_out3612_out1 <= Logical_Operator_out3100_out1 XOR Logical_Operator_out3164_out1;

  Logical_Operator_out3613_out1 <= Logical_Operator_out3101_out1 XOR Logical_Operator_out3165_out1;

  Logical_Operator_out3614_out1 <= Logical_Operator_out3102_out1 XOR Logical_Operator_out3166_out1;

  Logical_Operator_out3615_out1 <= Logical_Operator_out3103_out1 XOR Logical_Operator_out3167_out1;

  Logical_Operator_out3616_out1 <= Logical_Operator_out3104_out1 XOR Logical_Operator_out3168_out1;

  Logical_Operator_out3617_out1 <= Logical_Operator_out3105_out1 XOR Logical_Operator_out3169_out1;

  Logical_Operator_out3618_out1 <= Logical_Operator_out3106_out1 XOR Logical_Operator_out3170_out1;

  Logical_Operator_out3619_out1 <= Logical_Operator_out3107_out1 XOR Logical_Operator_out3171_out1;

  Logical_Operator_out3620_out1 <= Logical_Operator_out3108_out1 XOR Logical_Operator_out3172_out1;

  Logical_Operator_out3621_out1 <= Logical_Operator_out3109_out1 XOR Logical_Operator_out3173_out1;

  Logical_Operator_out3622_out1 <= Logical_Operator_out3110_out1 XOR Logical_Operator_out3174_out1;

  Logical_Operator_out3623_out1 <= Logical_Operator_out3111_out1 XOR Logical_Operator_out3175_out1;

  Logical_Operator_out3624_out1 <= Logical_Operator_out3112_out1 XOR Logical_Operator_out3176_out1;

  Logical_Operator_out3625_out1 <= Logical_Operator_out3113_out1 XOR Logical_Operator_out3177_out1;

  Logical_Operator_out3626_out1 <= Logical_Operator_out3114_out1 XOR Logical_Operator_out3178_out1;

  Logical_Operator_out3627_out1 <= Logical_Operator_out3115_out1 XOR Logical_Operator_out3179_out1;

  Logical_Operator_out3628_out1 <= Logical_Operator_out3116_out1 XOR Logical_Operator_out3180_out1;

  Logical_Operator_out3629_out1 <= Logical_Operator_out3117_out1 XOR Logical_Operator_out3181_out1;

  Logical_Operator_out3630_out1 <= Logical_Operator_out3118_out1 XOR Logical_Operator_out3182_out1;

  Logical_Operator_out3631_out1 <= Logical_Operator_out3119_out1 XOR Logical_Operator_out3183_out1;

  Logical_Operator_out3632_out1 <= Logical_Operator_out3120_out1 XOR Logical_Operator_out3184_out1;

  Logical_Operator_out3633_out1 <= Logical_Operator_out3121_out1 XOR Logical_Operator_out3185_out1;

  Logical_Operator_out3634_out1 <= Logical_Operator_out3122_out1 XOR Logical_Operator_out3186_out1;

  Logical_Operator_out3635_out1 <= Logical_Operator_out3123_out1 XOR Logical_Operator_out3187_out1;

  Logical_Operator_out3636_out1 <= Logical_Operator_out3124_out1 XOR Logical_Operator_out3188_out1;

  Logical_Operator_out3637_out1 <= Logical_Operator_out3125_out1 XOR Logical_Operator_out3189_out1;

  Logical_Operator_out3638_out1 <= Logical_Operator_out3126_out1 XOR Logical_Operator_out3190_out1;

  Logical_Operator_out3639_out1 <= Logical_Operator_out3127_out1 XOR Logical_Operator_out3191_out1;

  Logical_Operator_out3640_out1 <= Logical_Operator_out3128_out1 XOR Logical_Operator_out3192_out1;

  Logical_Operator_out3641_out1 <= Logical_Operator_out3129_out1 XOR Logical_Operator_out3193_out1;

  Logical_Operator_out3642_out1 <= Logical_Operator_out3130_out1 XOR Logical_Operator_out3194_out1;

  Logical_Operator_out3643_out1 <= Logical_Operator_out3131_out1 XOR Logical_Operator_out3195_out1;

  Logical_Operator_out3644_out1 <= Logical_Operator_out3132_out1 XOR Logical_Operator_out3196_out1;

  Logical_Operator_out3645_out1 <= Logical_Operator_out3133_out1 XOR Logical_Operator_out3197_out1;

  Logical_Operator_out3646_out1 <= Logical_Operator_out3134_out1 XOR Logical_Operator_out3198_out1;

  Logical_Operator_out3647_out1 <= Logical_Operator_out3135_out1 XOR Logical_Operator_out3199_out1;

  Logical_Operator_out3648_out1 <= Logical_Operator_out3136_out1 XOR Logical_Operator_out3200_out1;

  Logical_Operator_out3649_out1 <= Logical_Operator_out2593_out1 XOR Logical_Operator_out2657_out1;

  Logical_Operator_out3650_out1 <= Logical_Operator_out2594_out1 XOR Logical_Operator_out2658_out1;

  Logical_Operator_out3651_out1 <= Logical_Operator_out2595_out1 XOR Logical_Operator_out2659_out1;

  Logical_Operator_out3652_out1 <= Logical_Operator_out2596_out1 XOR Logical_Operator_out2660_out1;

  Logical_Operator_out3653_out1 <= Logical_Operator_out2597_out1 XOR Logical_Operator_out2661_out1;

  Logical_Operator_out3654_out1 <= Logical_Operator_out2598_out1 XOR Logical_Operator_out2662_out1;

  Logical_Operator_out3655_out1 <= Logical_Operator_out2599_out1 XOR Logical_Operator_out2663_out1;

  Logical_Operator_out3656_out1 <= Logical_Operator_out2600_out1 XOR Logical_Operator_out2664_out1;

  Logical_Operator_out3657_out1 <= Logical_Operator_out2601_out1 XOR Logical_Operator_out2665_out1;

  Logical_Operator_out3658_out1 <= Logical_Operator_out2602_out1 XOR Logical_Operator_out2666_out1;

  Logical_Operator_out3659_out1 <= Logical_Operator_out2603_out1 XOR Logical_Operator_out2667_out1;

  Logical_Operator_out3660_out1 <= Logical_Operator_out2604_out1 XOR Logical_Operator_out2668_out1;

  Logical_Operator_out3661_out1 <= Logical_Operator_out2605_out1 XOR Logical_Operator_out2669_out1;

  Logical_Operator_out3662_out1 <= Logical_Operator_out2606_out1 XOR Logical_Operator_out2670_out1;

  Logical_Operator_out3663_out1 <= Logical_Operator_out2607_out1 XOR Logical_Operator_out2671_out1;

  Logical_Operator_out3664_out1 <= Logical_Operator_out2608_out1 XOR Logical_Operator_out2672_out1;

  Logical_Operator_out3665_out1 <= Logical_Operator_out2609_out1 XOR Logical_Operator_out2673_out1;

  Logical_Operator_out3666_out1 <= Logical_Operator_out2610_out1 XOR Logical_Operator_out2674_out1;

  Logical_Operator_out3667_out1 <= Logical_Operator_out2611_out1 XOR Logical_Operator_out2675_out1;

  Logical_Operator_out3668_out1 <= Logical_Operator_out2612_out1 XOR Logical_Operator_out2676_out1;

  Logical_Operator_out3669_out1 <= Logical_Operator_out2613_out1 XOR Logical_Operator_out2677_out1;

  Logical_Operator_out3670_out1 <= Logical_Operator_out2614_out1 XOR Logical_Operator_out2678_out1;

  Logical_Operator_out3671_out1 <= Logical_Operator_out2615_out1 XOR Logical_Operator_out2679_out1;

  Logical_Operator_out3672_out1 <= Logical_Operator_out2616_out1 XOR Logical_Operator_out2680_out1;

  Logical_Operator_out3673_out1 <= Logical_Operator_out2617_out1 XOR Logical_Operator_out2681_out1;

  Logical_Operator_out3674_out1 <= Logical_Operator_out2618_out1 XOR Logical_Operator_out2682_out1;

  Logical_Operator_out3675_out1 <= Logical_Operator_out2619_out1 XOR Logical_Operator_out2683_out1;

  Logical_Operator_out3676_out1 <= Logical_Operator_out2620_out1 XOR Logical_Operator_out2684_out1;

  Logical_Operator_out3677_out1 <= Logical_Operator_out2621_out1 XOR Logical_Operator_out2685_out1;

  Logical_Operator_out3678_out1 <= Logical_Operator_out2622_out1 XOR Logical_Operator_out2686_out1;

  Logical_Operator_out3679_out1 <= Logical_Operator_out2623_out1 XOR Logical_Operator_out2687_out1;

  Logical_Operator_out3680_out1 <= Logical_Operator_out2624_out1 XOR Logical_Operator_out2688_out1;

  Logical_Operator_out3681_out1 <= Logical_Operator_out2097_out1 XOR Logical_Operator_out2161_out1;

  Logical_Operator_out3682_out1 <= Logical_Operator_out2098_out1 XOR Logical_Operator_out2162_out1;

  Logical_Operator_out3683_out1 <= Logical_Operator_out2099_out1 XOR Logical_Operator_out2163_out1;

  Logical_Operator_out3684_out1 <= Logical_Operator_out2100_out1 XOR Logical_Operator_out2164_out1;

  Logical_Operator_out3685_out1 <= Logical_Operator_out2101_out1 XOR Logical_Operator_out2165_out1;

  Logical_Operator_out3686_out1 <= Logical_Operator_out2102_out1 XOR Logical_Operator_out2166_out1;

  Logical_Operator_out3687_out1 <= Logical_Operator_out2103_out1 XOR Logical_Operator_out2167_out1;

  Logical_Operator_out3688_out1 <= Logical_Operator_out2104_out1 XOR Logical_Operator_out2168_out1;

  Logical_Operator_out3689_out1 <= Logical_Operator_out2105_out1 XOR Logical_Operator_out2169_out1;

  Logical_Operator_out3690_out1 <= Logical_Operator_out2106_out1 XOR Logical_Operator_out2170_out1;

  Logical_Operator_out3691_out1 <= Logical_Operator_out2107_out1 XOR Logical_Operator_out2171_out1;

  Logical_Operator_out3692_out1 <= Logical_Operator_out2108_out1 XOR Logical_Operator_out2172_out1;

  Logical_Operator_out3693_out1 <= Logical_Operator_out2109_out1 XOR Logical_Operator_out2173_out1;

  Logical_Operator_out3694_out1 <= Logical_Operator_out2110_out1 XOR Logical_Operator_out2174_out1;

  Logical_Operator_out3695_out1 <= Logical_Operator_out2111_out1 XOR Logical_Operator_out2175_out1;

  Logical_Operator_out3696_out1 <= Logical_Operator_out2112_out1 XOR Logical_Operator_out2176_out1;

  Logical_Operator_out3697_out1 <= Logical_Operator_out1593_out1 XOR Logical_Operator_out1657_out1;

  Logical_Operator_out3698_out1 <= Logical_Operator_out1594_out1 XOR Logical_Operator_out1658_out1;

  Logical_Operator_out3699_out1 <= Logical_Operator_out1595_out1 XOR Logical_Operator_out1659_out1;

  Logical_Operator_out3700_out1 <= Logical_Operator_out1596_out1 XOR Logical_Operator_out1660_out1;

  Logical_Operator_out3701_out1 <= Logical_Operator_out1597_out1 XOR Logical_Operator_out1661_out1;

  Logical_Operator_out3702_out1 <= Logical_Operator_out1598_out1 XOR Logical_Operator_out1662_out1;

  Logical_Operator_out3703_out1 <= Logical_Operator_out1599_out1 XOR Logical_Operator_out1663_out1;

  Logical_Operator_out3704_out1 <= Logical_Operator_out1600_out1 XOR Logical_Operator_out1664_out1;

  Logical_Operator_out3705_out1 <= Logical_Operator_out1085_out1 XOR Logical_Operator_out1149_out1;

  Logical_Operator_out3706_out1 <= Logical_Operator_out1086_out1 XOR Logical_Operator_out1150_out1;

  Logical_Operator_out3707_out1 <= Logical_Operator_out1087_out1 XOR Logical_Operator_out1151_out1;

  Logical_Operator_out3708_out1 <= Logical_Operator_out1088_out1 XOR Logical_Operator_out1152_out1;

  Logical_Operator_out3709_out1 <= Logical_Operator_out575_out1 XOR Logical_Operator_out639_out1;

  Logical_Operator_out3710_out1 <= Logical_Operator_out576_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out3711_out1 <= Logical_Operator_out64_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out3712_out1 <= in128 XOR in256;

  Logical_Operator_out3713_out1 <= Logical_Operator_out3201_out1 XOR Logical_Operator_out3265_out1;

  Logical_Operator_out3714_out1 <= Logical_Operator_out3202_out1 XOR Logical_Operator_out3266_out1;

  Logical_Operator_out3715_out1 <= Logical_Operator_out3203_out1 XOR Logical_Operator_out3267_out1;

  Logical_Operator_out3716_out1 <= Logical_Operator_out3204_out1 XOR Logical_Operator_out3268_out1;

  Logical_Operator_out3717_out1 <= Logical_Operator_out3205_out1 XOR Logical_Operator_out3269_out1;

  Logical_Operator_out3718_out1 <= Logical_Operator_out3206_out1 XOR Logical_Operator_out3270_out1;

  Logical_Operator_out3719_out1 <= Logical_Operator_out3207_out1 XOR Logical_Operator_out3271_out1;

  Logical_Operator_out3720_out1 <= Logical_Operator_out3208_out1 XOR Logical_Operator_out3272_out1;

  Logical_Operator_out3721_out1 <= Logical_Operator_out3209_out1 XOR Logical_Operator_out3273_out1;

  Logical_Operator_out3722_out1 <= Logical_Operator_out3210_out1 XOR Logical_Operator_out3274_out1;

  Logical_Operator_out3723_out1 <= Logical_Operator_out3211_out1 XOR Logical_Operator_out3275_out1;

  Logical_Operator_out3724_out1 <= Logical_Operator_out3212_out1 XOR Logical_Operator_out3276_out1;

  Logical_Operator_out3725_out1 <= Logical_Operator_out3213_out1 XOR Logical_Operator_out3277_out1;

  Logical_Operator_out3726_out1 <= Logical_Operator_out3214_out1 XOR Logical_Operator_out3278_out1;

  Logical_Operator_out3727_out1 <= Logical_Operator_out3215_out1 XOR Logical_Operator_out3279_out1;

  Logical_Operator_out3728_out1 <= Logical_Operator_out3216_out1 XOR Logical_Operator_out3280_out1;

  Logical_Operator_out3729_out1 <= Logical_Operator_out3217_out1 XOR Logical_Operator_out3281_out1;

  Logical_Operator_out3730_out1 <= Logical_Operator_out3218_out1 XOR Logical_Operator_out3282_out1;

  Logical_Operator_out3731_out1 <= Logical_Operator_out3219_out1 XOR Logical_Operator_out3283_out1;

  Logical_Operator_out3732_out1 <= Logical_Operator_out3220_out1 XOR Logical_Operator_out3284_out1;

  Logical_Operator_out3733_out1 <= Logical_Operator_out3221_out1 XOR Logical_Operator_out3285_out1;

  Logical_Operator_out3734_out1 <= Logical_Operator_out3222_out1 XOR Logical_Operator_out3286_out1;

  Logical_Operator_out3735_out1 <= Logical_Operator_out3223_out1 XOR Logical_Operator_out3287_out1;

  Logical_Operator_out3736_out1 <= Logical_Operator_out3224_out1 XOR Logical_Operator_out3288_out1;

  Logical_Operator_out3737_out1 <= Logical_Operator_out3225_out1 XOR Logical_Operator_out3289_out1;

  Logical_Operator_out3738_out1 <= Logical_Operator_out3226_out1 XOR Logical_Operator_out3290_out1;

  Logical_Operator_out3739_out1 <= Logical_Operator_out3227_out1 XOR Logical_Operator_out3291_out1;

  Logical_Operator_out3740_out1 <= Logical_Operator_out3228_out1 XOR Logical_Operator_out3292_out1;

  Logical_Operator_out3741_out1 <= Logical_Operator_out3229_out1 XOR Logical_Operator_out3293_out1;

  Logical_Operator_out3742_out1 <= Logical_Operator_out3230_out1 XOR Logical_Operator_out3294_out1;

  Logical_Operator_out3743_out1 <= Logical_Operator_out3231_out1 XOR Logical_Operator_out3295_out1;

  Logical_Operator_out3744_out1 <= Logical_Operator_out3232_out1 XOR Logical_Operator_out3296_out1;

  Logical_Operator_out3745_out1 <= Logical_Operator_out3233_out1 XOR Logical_Operator_out3297_out1;

  Logical_Operator_out3746_out1 <= Logical_Operator_out3234_out1 XOR Logical_Operator_out3298_out1;

  Logical_Operator_out3747_out1 <= Logical_Operator_out3235_out1 XOR Logical_Operator_out3299_out1;

  Logical_Operator_out3748_out1 <= Logical_Operator_out3236_out1 XOR Logical_Operator_out3300_out1;

  Logical_Operator_out3749_out1 <= Logical_Operator_out3237_out1 XOR Logical_Operator_out3301_out1;

  Logical_Operator_out3750_out1 <= Logical_Operator_out3238_out1 XOR Logical_Operator_out3302_out1;

  Logical_Operator_out3751_out1 <= Logical_Operator_out3239_out1 XOR Logical_Operator_out3303_out1;

  Logical_Operator_out3752_out1 <= Logical_Operator_out3240_out1 XOR Logical_Operator_out3304_out1;

  Logical_Operator_out3753_out1 <= Logical_Operator_out3241_out1 XOR Logical_Operator_out3305_out1;

  Logical_Operator_out3754_out1 <= Logical_Operator_out3242_out1 XOR Logical_Operator_out3306_out1;

  Logical_Operator_out3755_out1 <= Logical_Operator_out3243_out1 XOR Logical_Operator_out3307_out1;

  Logical_Operator_out3756_out1 <= Logical_Operator_out3244_out1 XOR Logical_Operator_out3308_out1;

  Logical_Operator_out3757_out1 <= Logical_Operator_out3245_out1 XOR Logical_Operator_out3309_out1;

  Logical_Operator_out3758_out1 <= Logical_Operator_out3246_out1 XOR Logical_Operator_out3310_out1;

  Logical_Operator_out3759_out1 <= Logical_Operator_out3247_out1 XOR Logical_Operator_out3311_out1;

  Logical_Operator_out3760_out1 <= Logical_Operator_out3248_out1 XOR Logical_Operator_out3312_out1;

  Logical_Operator_out3761_out1 <= Logical_Operator_out3249_out1 XOR Logical_Operator_out3313_out1;

  Logical_Operator_out3762_out1 <= Logical_Operator_out3250_out1 XOR Logical_Operator_out3314_out1;

  Logical_Operator_out3763_out1 <= Logical_Operator_out3251_out1 XOR Logical_Operator_out3315_out1;

  Logical_Operator_out3764_out1 <= Logical_Operator_out3252_out1 XOR Logical_Operator_out3316_out1;

  Logical_Operator_out3765_out1 <= Logical_Operator_out3253_out1 XOR Logical_Operator_out3317_out1;

  Logical_Operator_out3766_out1 <= Logical_Operator_out3254_out1 XOR Logical_Operator_out3318_out1;

  Logical_Operator_out3767_out1 <= Logical_Operator_out3255_out1 XOR Logical_Operator_out3319_out1;

  Logical_Operator_out3768_out1 <= Logical_Operator_out3256_out1 XOR Logical_Operator_out3320_out1;

  Logical_Operator_out3769_out1 <= Logical_Operator_out3257_out1 XOR Logical_Operator_out3321_out1;

  Logical_Operator_out3770_out1 <= Logical_Operator_out3258_out1 XOR Logical_Operator_out3322_out1;

  Logical_Operator_out3771_out1 <= Logical_Operator_out3259_out1 XOR Logical_Operator_out3323_out1;

  Logical_Operator_out3772_out1 <= Logical_Operator_out3260_out1 XOR Logical_Operator_out3324_out1;

  Logical_Operator_out3773_out1 <= Logical_Operator_out3261_out1 XOR Logical_Operator_out3325_out1;

  Logical_Operator_out3774_out1 <= Logical_Operator_out3262_out1 XOR Logical_Operator_out3326_out1;

  Logical_Operator_out3775_out1 <= Logical_Operator_out3263_out1 XOR Logical_Operator_out3327_out1;

  Logical_Operator_out3776_out1 <= Logical_Operator_out3264_out1 XOR Logical_Operator_out3328_out1;

  Logical_Operator_out3777_out1 <= Logical_Operator_out2721_out1 XOR Logical_Operator_out2785_out1;

  Logical_Operator_out3778_out1 <= Logical_Operator_out2722_out1 XOR Logical_Operator_out2786_out1;

  Logical_Operator_out3779_out1 <= Logical_Operator_out2723_out1 XOR Logical_Operator_out2787_out1;

  Logical_Operator_out3780_out1 <= Logical_Operator_out2724_out1 XOR Logical_Operator_out2788_out1;

  Logical_Operator_out3781_out1 <= Logical_Operator_out2725_out1 XOR Logical_Operator_out2789_out1;

  Logical_Operator_out3782_out1 <= Logical_Operator_out2726_out1 XOR Logical_Operator_out2790_out1;

  Logical_Operator_out3783_out1 <= Logical_Operator_out2727_out1 XOR Logical_Operator_out2791_out1;

  Logical_Operator_out3784_out1 <= Logical_Operator_out2728_out1 XOR Logical_Operator_out2792_out1;

  Logical_Operator_out3785_out1 <= Logical_Operator_out2729_out1 XOR Logical_Operator_out2793_out1;

  Logical_Operator_out3786_out1 <= Logical_Operator_out2730_out1 XOR Logical_Operator_out2794_out1;

  Logical_Operator_out3787_out1 <= Logical_Operator_out2731_out1 XOR Logical_Operator_out2795_out1;

  Logical_Operator_out3788_out1 <= Logical_Operator_out2732_out1 XOR Logical_Operator_out2796_out1;

  Logical_Operator_out3789_out1 <= Logical_Operator_out2733_out1 XOR Logical_Operator_out2797_out1;

  Logical_Operator_out3790_out1 <= Logical_Operator_out2734_out1 XOR Logical_Operator_out2798_out1;

  Logical_Operator_out3791_out1 <= Logical_Operator_out2735_out1 XOR Logical_Operator_out2799_out1;

  Logical_Operator_out3792_out1 <= Logical_Operator_out2736_out1 XOR Logical_Operator_out2800_out1;

  Logical_Operator_out3793_out1 <= Logical_Operator_out2737_out1 XOR Logical_Operator_out2801_out1;

  Logical_Operator_out3794_out1 <= Logical_Operator_out2738_out1 XOR Logical_Operator_out2802_out1;

  Logical_Operator_out3795_out1 <= Logical_Operator_out2739_out1 XOR Logical_Operator_out2803_out1;

  Logical_Operator_out3796_out1 <= Logical_Operator_out2740_out1 XOR Logical_Operator_out2804_out1;

  Logical_Operator_out3797_out1 <= Logical_Operator_out2741_out1 XOR Logical_Operator_out2805_out1;

  Logical_Operator_out3798_out1 <= Logical_Operator_out2742_out1 XOR Logical_Operator_out2806_out1;

  Logical_Operator_out3799_out1 <= Logical_Operator_out2743_out1 XOR Logical_Operator_out2807_out1;

  Logical_Operator_out3800_out1 <= Logical_Operator_out2744_out1 XOR Logical_Operator_out2808_out1;

  Logical_Operator_out3801_out1 <= Logical_Operator_out2745_out1 XOR Logical_Operator_out2809_out1;

  Logical_Operator_out3802_out1 <= Logical_Operator_out2746_out1 XOR Logical_Operator_out2810_out1;

  Logical_Operator_out3803_out1 <= Logical_Operator_out2747_out1 XOR Logical_Operator_out2811_out1;

  Logical_Operator_out3804_out1 <= Logical_Operator_out2748_out1 XOR Logical_Operator_out2812_out1;

  Logical_Operator_out3805_out1 <= Logical_Operator_out2749_out1 XOR Logical_Operator_out2813_out1;

  Logical_Operator_out3806_out1 <= Logical_Operator_out2750_out1 XOR Logical_Operator_out2814_out1;

  Logical_Operator_out3807_out1 <= Logical_Operator_out2751_out1 XOR Logical_Operator_out2815_out1;

  Logical_Operator_out3808_out1 <= Logical_Operator_out2752_out1 XOR Logical_Operator_out2816_out1;

  Logical_Operator_out3809_out1 <= Logical_Operator_out2225_out1 XOR Logical_Operator_out2289_out1;

  Logical_Operator_out3810_out1 <= Logical_Operator_out2226_out1 XOR Logical_Operator_out2290_out1;

  Logical_Operator_out3811_out1 <= Logical_Operator_out2227_out1 XOR Logical_Operator_out2291_out1;

  Logical_Operator_out3812_out1 <= Logical_Operator_out2228_out1 XOR Logical_Operator_out2292_out1;

  Logical_Operator_out3813_out1 <= Logical_Operator_out2229_out1 XOR Logical_Operator_out2293_out1;

  Logical_Operator_out3814_out1 <= Logical_Operator_out2230_out1 XOR Logical_Operator_out2294_out1;

  Logical_Operator_out3815_out1 <= Logical_Operator_out2231_out1 XOR Logical_Operator_out2295_out1;

  Logical_Operator_out3816_out1 <= Logical_Operator_out2232_out1 XOR Logical_Operator_out2296_out1;

  Logical_Operator_out3817_out1 <= Logical_Operator_out2233_out1 XOR Logical_Operator_out2297_out1;

  Logical_Operator_out3818_out1 <= Logical_Operator_out2234_out1 XOR Logical_Operator_out2298_out1;

  Logical_Operator_out3819_out1 <= Logical_Operator_out2235_out1 XOR Logical_Operator_out2299_out1;

  Logical_Operator_out3820_out1 <= Logical_Operator_out2236_out1 XOR Logical_Operator_out2300_out1;

  Logical_Operator_out3821_out1 <= Logical_Operator_out2237_out1 XOR Logical_Operator_out2301_out1;

  Logical_Operator_out3822_out1 <= Logical_Operator_out2238_out1 XOR Logical_Operator_out2302_out1;

  Logical_Operator_out3823_out1 <= Logical_Operator_out2239_out1 XOR Logical_Operator_out2303_out1;

  Logical_Operator_out3824_out1 <= Logical_Operator_out2240_out1 XOR Logical_Operator_out2304_out1;

  Logical_Operator_out3825_out1 <= Logical_Operator_out1721_out1 XOR Logical_Operator_out1785_out1;

  Logical_Operator_out3826_out1 <= Logical_Operator_out1722_out1 XOR Logical_Operator_out1786_out1;

  Logical_Operator_out3827_out1 <= Logical_Operator_out1723_out1 XOR Logical_Operator_out1787_out1;

  Logical_Operator_out3828_out1 <= Logical_Operator_out1724_out1 XOR Logical_Operator_out1788_out1;

  Logical_Operator_out3829_out1 <= Logical_Operator_out1725_out1 XOR Logical_Operator_out1789_out1;

  Logical_Operator_out3830_out1 <= Logical_Operator_out1726_out1 XOR Logical_Operator_out1790_out1;

  Logical_Operator_out3831_out1 <= Logical_Operator_out1727_out1 XOR Logical_Operator_out1791_out1;

  Logical_Operator_out3832_out1 <= Logical_Operator_out1728_out1 XOR Logical_Operator_out1792_out1;

  Logical_Operator_out3833_out1 <= Logical_Operator_out1213_out1 XOR Logical_Operator_out1277_out1;

  Logical_Operator_out3834_out1 <= Logical_Operator_out1214_out1 XOR Logical_Operator_out1278_out1;

  Logical_Operator_out3835_out1 <= Logical_Operator_out1215_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out3836_out1 <= Logical_Operator_out1216_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out3837_out1 <= Logical_Operator_out703_out1 XOR Logical_Operator_out767_out1;

  Logical_Operator_out3838_out1 <= Logical_Operator_out704_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out3839_out1 <= Logical_Operator_out192_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out3840_out1 <= in384 XOR in512;

  Logical_Operator_out3841_out1 <= Logical_Operator_out3329_out1 XOR Logical_Operator_out3393_out1;

  Logical_Operator_out3842_out1 <= Logical_Operator_out3330_out1 XOR Logical_Operator_out3394_out1;

  Logical_Operator_out3843_out1 <= Logical_Operator_out3331_out1 XOR Logical_Operator_out3395_out1;

  Logical_Operator_out3844_out1 <= Logical_Operator_out3332_out1 XOR Logical_Operator_out3396_out1;

  Logical_Operator_out3845_out1 <= Logical_Operator_out3333_out1 XOR Logical_Operator_out3397_out1;

  Logical_Operator_out3846_out1 <= Logical_Operator_out3334_out1 XOR Logical_Operator_out3398_out1;

  Logical_Operator_out3847_out1 <= Logical_Operator_out3335_out1 XOR Logical_Operator_out3399_out1;

  Logical_Operator_out3848_out1 <= Logical_Operator_out3336_out1 XOR Logical_Operator_out3400_out1;

  Logical_Operator_out3849_out1 <= Logical_Operator_out3337_out1 XOR Logical_Operator_out3401_out1;

  Logical_Operator_out3850_out1 <= Logical_Operator_out3338_out1 XOR Logical_Operator_out3402_out1;

  Logical_Operator_out3851_out1 <= Logical_Operator_out3339_out1 XOR Logical_Operator_out3403_out1;

  Logical_Operator_out3852_out1 <= Logical_Operator_out3340_out1 XOR Logical_Operator_out3404_out1;

  Logical_Operator_out3853_out1 <= Logical_Operator_out3341_out1 XOR Logical_Operator_out3405_out1;

  Logical_Operator_out3854_out1 <= Logical_Operator_out3342_out1 XOR Logical_Operator_out3406_out1;

  Logical_Operator_out3855_out1 <= Logical_Operator_out3343_out1 XOR Logical_Operator_out3407_out1;

  Logical_Operator_out3856_out1 <= Logical_Operator_out3344_out1 XOR Logical_Operator_out3408_out1;

  Logical_Operator_out3857_out1 <= Logical_Operator_out3345_out1 XOR Logical_Operator_out3409_out1;

  Logical_Operator_out3858_out1 <= Logical_Operator_out3346_out1 XOR Logical_Operator_out3410_out1;

  Logical_Operator_out3859_out1 <= Logical_Operator_out3347_out1 XOR Logical_Operator_out3411_out1;

  Logical_Operator_out3860_out1 <= Logical_Operator_out3348_out1 XOR Logical_Operator_out3412_out1;

  Logical_Operator_out3861_out1 <= Logical_Operator_out3349_out1 XOR Logical_Operator_out3413_out1;

  Logical_Operator_out3862_out1 <= Logical_Operator_out3350_out1 XOR Logical_Operator_out3414_out1;

  Logical_Operator_out3863_out1 <= Logical_Operator_out3351_out1 XOR Logical_Operator_out3415_out1;

  Logical_Operator_out3864_out1 <= Logical_Operator_out3352_out1 XOR Logical_Operator_out3416_out1;

  Logical_Operator_out3865_out1 <= Logical_Operator_out3353_out1 XOR Logical_Operator_out3417_out1;

  Logical_Operator_out3866_out1 <= Logical_Operator_out3354_out1 XOR Logical_Operator_out3418_out1;

  Logical_Operator_out3867_out1 <= Logical_Operator_out3355_out1 XOR Logical_Operator_out3419_out1;

  Logical_Operator_out3868_out1 <= Logical_Operator_out3356_out1 XOR Logical_Operator_out3420_out1;

  Logical_Operator_out3869_out1 <= Logical_Operator_out3357_out1 XOR Logical_Operator_out3421_out1;

  Logical_Operator_out3870_out1 <= Logical_Operator_out3358_out1 XOR Logical_Operator_out3422_out1;

  Logical_Operator_out3871_out1 <= Logical_Operator_out3359_out1 XOR Logical_Operator_out3423_out1;

  Logical_Operator_out3872_out1 <= Logical_Operator_out3360_out1 XOR Logical_Operator_out3424_out1;

  Logical_Operator_out3873_out1 <= Logical_Operator_out3361_out1 XOR Logical_Operator_out3425_out1;

  Logical_Operator_out3874_out1 <= Logical_Operator_out3362_out1 XOR Logical_Operator_out3426_out1;

  Logical_Operator_out3875_out1 <= Logical_Operator_out3363_out1 XOR Logical_Operator_out3427_out1;

  Logical_Operator_out3876_out1 <= Logical_Operator_out3364_out1 XOR Logical_Operator_out3428_out1;

  Logical_Operator_out3877_out1 <= Logical_Operator_out3365_out1 XOR Logical_Operator_out3429_out1;

  Logical_Operator_out3878_out1 <= Logical_Operator_out3366_out1 XOR Logical_Operator_out3430_out1;

  Logical_Operator_out3879_out1 <= Logical_Operator_out3367_out1 XOR Logical_Operator_out3431_out1;

  Logical_Operator_out3880_out1 <= Logical_Operator_out3368_out1 XOR Logical_Operator_out3432_out1;

  Logical_Operator_out3881_out1 <= Logical_Operator_out3369_out1 XOR Logical_Operator_out3433_out1;

  Logical_Operator_out3882_out1 <= Logical_Operator_out3370_out1 XOR Logical_Operator_out3434_out1;

  Logical_Operator_out3883_out1 <= Logical_Operator_out3371_out1 XOR Logical_Operator_out3435_out1;

  Logical_Operator_out3884_out1 <= Logical_Operator_out3372_out1 XOR Logical_Operator_out3436_out1;

  Logical_Operator_out3885_out1 <= Logical_Operator_out3373_out1 XOR Logical_Operator_out3437_out1;

  Logical_Operator_out3886_out1 <= Logical_Operator_out3374_out1 XOR Logical_Operator_out3438_out1;

  Logical_Operator_out3887_out1 <= Logical_Operator_out3375_out1 XOR Logical_Operator_out3439_out1;

  Logical_Operator_out3888_out1 <= Logical_Operator_out3376_out1 XOR Logical_Operator_out3440_out1;

  Logical_Operator_out3889_out1 <= Logical_Operator_out3377_out1 XOR Logical_Operator_out3441_out1;

  Logical_Operator_out3890_out1 <= Logical_Operator_out3378_out1 XOR Logical_Operator_out3442_out1;

  Logical_Operator_out3891_out1 <= Logical_Operator_out3379_out1 XOR Logical_Operator_out3443_out1;

  Logical_Operator_out3892_out1 <= Logical_Operator_out3380_out1 XOR Logical_Operator_out3444_out1;

  Logical_Operator_out3893_out1 <= Logical_Operator_out3381_out1 XOR Logical_Operator_out3445_out1;

  Logical_Operator_out3894_out1 <= Logical_Operator_out3382_out1 XOR Logical_Operator_out3446_out1;

  Logical_Operator_out3895_out1 <= Logical_Operator_out3383_out1 XOR Logical_Operator_out3447_out1;

  Logical_Operator_out3896_out1 <= Logical_Operator_out3384_out1 XOR Logical_Operator_out3448_out1;

  Logical_Operator_out3897_out1 <= Logical_Operator_out3385_out1 XOR Logical_Operator_out3449_out1;

  Logical_Operator_out3898_out1 <= Logical_Operator_out3386_out1 XOR Logical_Operator_out3450_out1;

  Logical_Operator_out3899_out1 <= Logical_Operator_out3387_out1 XOR Logical_Operator_out3451_out1;

  Logical_Operator_out3900_out1 <= Logical_Operator_out3388_out1 XOR Logical_Operator_out3452_out1;

  Logical_Operator_out3901_out1 <= Logical_Operator_out3389_out1 XOR Logical_Operator_out3453_out1;

  Logical_Operator_out3902_out1 <= Logical_Operator_out3390_out1 XOR Logical_Operator_out3454_out1;

  Logical_Operator_out3903_out1 <= Logical_Operator_out3391_out1 XOR Logical_Operator_out3455_out1;

  Logical_Operator_out3904_out1 <= Logical_Operator_out3392_out1 XOR Logical_Operator_out3456_out1;

  Logical_Operator_out3905_out1 <= Logical_Operator_out2849_out1 XOR Logical_Operator_out2913_out1;

  Logical_Operator_out3906_out1 <= Logical_Operator_out2850_out1 XOR Logical_Operator_out2914_out1;

  Logical_Operator_out3907_out1 <= Logical_Operator_out2851_out1 XOR Logical_Operator_out2915_out1;

  Logical_Operator_out3908_out1 <= Logical_Operator_out2852_out1 XOR Logical_Operator_out2916_out1;

  Logical_Operator_out3909_out1 <= Logical_Operator_out2853_out1 XOR Logical_Operator_out2917_out1;

  Logical_Operator_out3910_out1 <= Logical_Operator_out2854_out1 XOR Logical_Operator_out2918_out1;

  Logical_Operator_out3911_out1 <= Logical_Operator_out2855_out1 XOR Logical_Operator_out2919_out1;

  Logical_Operator_out3912_out1 <= Logical_Operator_out2856_out1 XOR Logical_Operator_out2920_out1;

  Logical_Operator_out3913_out1 <= Logical_Operator_out2857_out1 XOR Logical_Operator_out2921_out1;

  Logical_Operator_out3914_out1 <= Logical_Operator_out2858_out1 XOR Logical_Operator_out2922_out1;

  Logical_Operator_out3915_out1 <= Logical_Operator_out2859_out1 XOR Logical_Operator_out2923_out1;

  Logical_Operator_out3916_out1 <= Logical_Operator_out2860_out1 XOR Logical_Operator_out2924_out1;

  Logical_Operator_out3917_out1 <= Logical_Operator_out2861_out1 XOR Logical_Operator_out2925_out1;

  Logical_Operator_out3918_out1 <= Logical_Operator_out2862_out1 XOR Logical_Operator_out2926_out1;

  Logical_Operator_out3919_out1 <= Logical_Operator_out2863_out1 XOR Logical_Operator_out2927_out1;

  Logical_Operator_out3920_out1 <= Logical_Operator_out2864_out1 XOR Logical_Operator_out2928_out1;

  Logical_Operator_out3921_out1 <= Logical_Operator_out2865_out1 XOR Logical_Operator_out2929_out1;

  Logical_Operator_out3922_out1 <= Logical_Operator_out2866_out1 XOR Logical_Operator_out2930_out1;

  Logical_Operator_out3923_out1 <= Logical_Operator_out2867_out1 XOR Logical_Operator_out2931_out1;

  Logical_Operator_out3924_out1 <= Logical_Operator_out2868_out1 XOR Logical_Operator_out2932_out1;

  Logical_Operator_out3925_out1 <= Logical_Operator_out2869_out1 XOR Logical_Operator_out2933_out1;

  Logical_Operator_out3926_out1 <= Logical_Operator_out2870_out1 XOR Logical_Operator_out2934_out1;

  Logical_Operator_out3927_out1 <= Logical_Operator_out2871_out1 XOR Logical_Operator_out2935_out1;

  Logical_Operator_out3928_out1 <= Logical_Operator_out2872_out1 XOR Logical_Operator_out2936_out1;

  Logical_Operator_out3929_out1 <= Logical_Operator_out2873_out1 XOR Logical_Operator_out2937_out1;

  Logical_Operator_out3930_out1 <= Logical_Operator_out2874_out1 XOR Logical_Operator_out2938_out1;

  Logical_Operator_out3931_out1 <= Logical_Operator_out2875_out1 XOR Logical_Operator_out2939_out1;

  Logical_Operator_out3932_out1 <= Logical_Operator_out2876_out1 XOR Logical_Operator_out2940_out1;

  Logical_Operator_out3933_out1 <= Logical_Operator_out2877_out1 XOR Logical_Operator_out2941_out1;

  Logical_Operator_out3934_out1 <= Logical_Operator_out2878_out1 XOR Logical_Operator_out2942_out1;

  Logical_Operator_out3935_out1 <= Logical_Operator_out2879_out1 XOR Logical_Operator_out2943_out1;

  Logical_Operator_out3936_out1 <= Logical_Operator_out2880_out1 XOR Logical_Operator_out2944_out1;

  Logical_Operator_out3937_out1 <= Logical_Operator_out2353_out1 XOR Logical_Operator_out2417_out1;

  Logical_Operator_out3938_out1 <= Logical_Operator_out2354_out1 XOR Logical_Operator_out2418_out1;

  Logical_Operator_out3939_out1 <= Logical_Operator_out2355_out1 XOR Logical_Operator_out2419_out1;

  Logical_Operator_out3940_out1 <= Logical_Operator_out2356_out1 XOR Logical_Operator_out2420_out1;

  Logical_Operator_out3941_out1 <= Logical_Operator_out2357_out1 XOR Logical_Operator_out2421_out1;

  Logical_Operator_out3942_out1 <= Logical_Operator_out2358_out1 XOR Logical_Operator_out2422_out1;

  Logical_Operator_out3943_out1 <= Logical_Operator_out2359_out1 XOR Logical_Operator_out2423_out1;

  Logical_Operator_out3944_out1 <= Logical_Operator_out2360_out1 XOR Logical_Operator_out2424_out1;

  Logical_Operator_out3945_out1 <= Logical_Operator_out2361_out1 XOR Logical_Operator_out2425_out1;

  Logical_Operator_out3946_out1 <= Logical_Operator_out2362_out1 XOR Logical_Operator_out2426_out1;

  Logical_Operator_out3947_out1 <= Logical_Operator_out2363_out1 XOR Logical_Operator_out2427_out1;

  Logical_Operator_out3948_out1 <= Logical_Operator_out2364_out1 XOR Logical_Operator_out2428_out1;

  Logical_Operator_out3949_out1 <= Logical_Operator_out2365_out1 XOR Logical_Operator_out2429_out1;

  Logical_Operator_out3950_out1 <= Logical_Operator_out2366_out1 XOR Logical_Operator_out2430_out1;

  Logical_Operator_out3951_out1 <= Logical_Operator_out2367_out1 XOR Logical_Operator_out2431_out1;

  Logical_Operator_out3952_out1 <= Logical_Operator_out2368_out1 XOR Logical_Operator_out2432_out1;

  Logical_Operator_out3953_out1 <= Logical_Operator_out1849_out1 XOR Logical_Operator_out1913_out1;

  Logical_Operator_out3954_out1 <= Logical_Operator_out1850_out1 XOR Logical_Operator_out1914_out1;

  Logical_Operator_out3955_out1 <= Logical_Operator_out1851_out1 XOR Logical_Operator_out1915_out1;

  Logical_Operator_out3956_out1 <= Logical_Operator_out1852_out1 XOR Logical_Operator_out1916_out1;

  Logical_Operator_out3957_out1 <= Logical_Operator_out1853_out1 XOR Logical_Operator_out1917_out1;

  Logical_Operator_out3958_out1 <= Logical_Operator_out1854_out1 XOR Logical_Operator_out1918_out1;

  Logical_Operator_out3959_out1 <= Logical_Operator_out1855_out1 XOR Logical_Operator_out1919_out1;

  Logical_Operator_out3960_out1 <= Logical_Operator_out1856_out1 XOR Logical_Operator_out1920_out1;

  Logical_Operator_out3961_out1 <= Logical_Operator_out1341_out1 XOR Logical_Operator_out1405_out1;

  Logical_Operator_out3962_out1 <= Logical_Operator_out1342_out1 XOR Logical_Operator_out1406_out1;

  Logical_Operator_out3963_out1 <= Logical_Operator_out1343_out1 XOR Logical_Operator_out1407_out1;

  Logical_Operator_out3964_out1 <= Logical_Operator_out1344_out1 XOR Logical_Operator_out1408_out1;

  Logical_Operator_out3965_out1 <= Logical_Operator_out831_out1 XOR Logical_Operator_out895_out1;

  Logical_Operator_out3966_out1 <= Logical_Operator_out832_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out3967_out1 <= Logical_Operator_out320_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out3968_out1 <= in640 XOR in768;

  Logical_Operator_out3969_out1 <= Logical_Operator_out3457_out1 XOR Logical_Operator_out3521_out1;

  Logical_Operator_out3970_out1 <= Logical_Operator_out3458_out1 XOR Logical_Operator_out3522_out1;

  Logical_Operator_out3971_out1 <= Logical_Operator_out3459_out1 XOR Logical_Operator_out3523_out1;

  Logical_Operator_out3972_out1 <= Logical_Operator_out3460_out1 XOR Logical_Operator_out3524_out1;

  Logical_Operator_out3973_out1 <= Logical_Operator_out3461_out1 XOR Logical_Operator_out3525_out1;

  Logical_Operator_out3974_out1 <= Logical_Operator_out3462_out1 XOR Logical_Operator_out3526_out1;

  Logical_Operator_out3975_out1 <= Logical_Operator_out3463_out1 XOR Logical_Operator_out3527_out1;

  Logical_Operator_out3976_out1 <= Logical_Operator_out3464_out1 XOR Logical_Operator_out3528_out1;

  Logical_Operator_out3977_out1 <= Logical_Operator_out3465_out1 XOR Logical_Operator_out3529_out1;

  Logical_Operator_out3978_out1 <= Logical_Operator_out3466_out1 XOR Logical_Operator_out3530_out1;

  Logical_Operator_out3979_out1 <= Logical_Operator_out3467_out1 XOR Logical_Operator_out3531_out1;

  Logical_Operator_out3980_out1 <= Logical_Operator_out3468_out1 XOR Logical_Operator_out3532_out1;

  Logical_Operator_out3981_out1 <= Logical_Operator_out3469_out1 XOR Logical_Operator_out3533_out1;

  Logical_Operator_out3982_out1 <= Logical_Operator_out3470_out1 XOR Logical_Operator_out3534_out1;

  Logical_Operator_out3983_out1 <= Logical_Operator_out3471_out1 XOR Logical_Operator_out3535_out1;

  Logical_Operator_out3984_out1 <= Logical_Operator_out3472_out1 XOR Logical_Operator_out3536_out1;

  Logical_Operator_out3985_out1 <= Logical_Operator_out3473_out1 XOR Logical_Operator_out3537_out1;

  Logical_Operator_out3986_out1 <= Logical_Operator_out3474_out1 XOR Logical_Operator_out3538_out1;

  Logical_Operator_out3987_out1 <= Logical_Operator_out3475_out1 XOR Logical_Operator_out3539_out1;

  Logical_Operator_out3988_out1 <= Logical_Operator_out3476_out1 XOR Logical_Operator_out3540_out1;

  Logical_Operator_out3989_out1 <= Logical_Operator_out3477_out1 XOR Logical_Operator_out3541_out1;

  Logical_Operator_out3990_out1 <= Logical_Operator_out3478_out1 XOR Logical_Operator_out3542_out1;

  Logical_Operator_out3991_out1 <= Logical_Operator_out3479_out1 XOR Logical_Operator_out3543_out1;

  Logical_Operator_out3992_out1 <= Logical_Operator_out3480_out1 XOR Logical_Operator_out3544_out1;

  Logical_Operator_out3993_out1 <= Logical_Operator_out3481_out1 XOR Logical_Operator_out3545_out1;

  Logical_Operator_out3994_out1 <= Logical_Operator_out3482_out1 XOR Logical_Operator_out3546_out1;

  Logical_Operator_out3995_out1 <= Logical_Operator_out3483_out1 XOR Logical_Operator_out3547_out1;

  Logical_Operator_out3996_out1 <= Logical_Operator_out3484_out1 XOR Logical_Operator_out3548_out1;

  Logical_Operator_out3997_out1 <= Logical_Operator_out3485_out1 XOR Logical_Operator_out3549_out1;

  Logical_Operator_out3998_out1 <= Logical_Operator_out3486_out1 XOR Logical_Operator_out3550_out1;

  Logical_Operator_out3999_out1 <= Logical_Operator_out3487_out1 XOR Logical_Operator_out3551_out1;

  Logical_Operator_out4000_out1 <= Logical_Operator_out3488_out1 XOR Logical_Operator_out3552_out1;

  Logical_Operator_out4001_out1 <= Logical_Operator_out3489_out1 XOR Logical_Operator_out3553_out1;

  Logical_Operator_out4002_out1 <= Logical_Operator_out3490_out1 XOR Logical_Operator_out3554_out1;

  Logical_Operator_out4003_out1 <= Logical_Operator_out3491_out1 XOR Logical_Operator_out3555_out1;

  Logical_Operator_out4004_out1 <= Logical_Operator_out3492_out1 XOR Logical_Operator_out3556_out1;

  Logical_Operator_out4005_out1 <= Logical_Operator_out3493_out1 XOR Logical_Operator_out3557_out1;

  Logical_Operator_out4006_out1 <= Logical_Operator_out3494_out1 XOR Logical_Operator_out3558_out1;

  Logical_Operator_out4007_out1 <= Logical_Operator_out3495_out1 XOR Logical_Operator_out3559_out1;

  Logical_Operator_out4008_out1 <= Logical_Operator_out3496_out1 XOR Logical_Operator_out3560_out1;

  Logical_Operator_out4009_out1 <= Logical_Operator_out3497_out1 XOR Logical_Operator_out3561_out1;

  Logical_Operator_out4010_out1 <= Logical_Operator_out3498_out1 XOR Logical_Operator_out3562_out1;

  Logical_Operator_out4011_out1 <= Logical_Operator_out3499_out1 XOR Logical_Operator_out3563_out1;

  Logical_Operator_out4012_out1 <= Logical_Operator_out3500_out1 XOR Logical_Operator_out3564_out1;

  Logical_Operator_out4013_out1 <= Logical_Operator_out3501_out1 XOR Logical_Operator_out3565_out1;

  Logical_Operator_out4014_out1 <= Logical_Operator_out3502_out1 XOR Logical_Operator_out3566_out1;

  Logical_Operator_out4015_out1 <= Logical_Operator_out3503_out1 XOR Logical_Operator_out3567_out1;

  Logical_Operator_out4016_out1 <= Logical_Operator_out3504_out1 XOR Logical_Operator_out3568_out1;

  Logical_Operator_out4017_out1 <= Logical_Operator_out3505_out1 XOR Logical_Operator_out3569_out1;

  Logical_Operator_out4018_out1 <= Logical_Operator_out3506_out1 XOR Logical_Operator_out3570_out1;

  Logical_Operator_out4019_out1 <= Logical_Operator_out3507_out1 XOR Logical_Operator_out3571_out1;

  Logical_Operator_out4020_out1 <= Logical_Operator_out3508_out1 XOR Logical_Operator_out3572_out1;

  Logical_Operator_out4021_out1 <= Logical_Operator_out3509_out1 XOR Logical_Operator_out3573_out1;

  Logical_Operator_out4022_out1 <= Logical_Operator_out3510_out1 XOR Logical_Operator_out3574_out1;

  Logical_Operator_out4023_out1 <= Logical_Operator_out3511_out1 XOR Logical_Operator_out3575_out1;

  Logical_Operator_out4024_out1 <= Logical_Operator_out3512_out1 XOR Logical_Operator_out3576_out1;

  Logical_Operator_out4025_out1 <= Logical_Operator_out3513_out1 XOR Logical_Operator_out3577_out1;

  Logical_Operator_out4026_out1 <= Logical_Operator_out3514_out1 XOR Logical_Operator_out3578_out1;

  Logical_Operator_out4027_out1 <= Logical_Operator_out3515_out1 XOR Logical_Operator_out3579_out1;

  Logical_Operator_out4028_out1 <= Logical_Operator_out3516_out1 XOR Logical_Operator_out3580_out1;

  Logical_Operator_out4029_out1 <= Logical_Operator_out3517_out1 XOR Logical_Operator_out3581_out1;

  Logical_Operator_out4030_out1 <= Logical_Operator_out3518_out1 XOR Logical_Operator_out3582_out1;

  Logical_Operator_out4031_out1 <= Logical_Operator_out3519_out1 XOR Logical_Operator_out3583_out1;

  Logical_Operator_out4032_out1 <= Logical_Operator_out3520_out1 XOR Logical_Operator_out3584_out1;

  Logical_Operator_out4033_out1 <= Logical_Operator_out2977_out1 XOR Logical_Operator_out3041_out1;

  Logical_Operator_out4034_out1 <= Logical_Operator_out2978_out1 XOR Logical_Operator_out3042_out1;

  Logical_Operator_out4035_out1 <= Logical_Operator_out2979_out1 XOR Logical_Operator_out3043_out1;

  Logical_Operator_out4036_out1 <= Logical_Operator_out2980_out1 XOR Logical_Operator_out3044_out1;

  Logical_Operator_out4037_out1 <= Logical_Operator_out2981_out1 XOR Logical_Operator_out3045_out1;

  Logical_Operator_out4038_out1 <= Logical_Operator_out2982_out1 XOR Logical_Operator_out3046_out1;

  Logical_Operator_out4039_out1 <= Logical_Operator_out2983_out1 XOR Logical_Operator_out3047_out1;

  Logical_Operator_out4040_out1 <= Logical_Operator_out2984_out1 XOR Logical_Operator_out3048_out1;

  Logical_Operator_out4041_out1 <= Logical_Operator_out2985_out1 XOR Logical_Operator_out3049_out1;

  Logical_Operator_out4042_out1 <= Logical_Operator_out2986_out1 XOR Logical_Operator_out3050_out1;

  Logical_Operator_out4043_out1 <= Logical_Operator_out2987_out1 XOR Logical_Operator_out3051_out1;

  Logical_Operator_out4044_out1 <= Logical_Operator_out2988_out1 XOR Logical_Operator_out3052_out1;

  Logical_Operator_out4045_out1 <= Logical_Operator_out2989_out1 XOR Logical_Operator_out3053_out1;

  Logical_Operator_out4046_out1 <= Logical_Operator_out2990_out1 XOR Logical_Operator_out3054_out1;

  Logical_Operator_out4047_out1 <= Logical_Operator_out2991_out1 XOR Logical_Operator_out3055_out1;

  Logical_Operator_out4048_out1 <= Logical_Operator_out2992_out1 XOR Logical_Operator_out3056_out1;

  Logical_Operator_out4049_out1 <= Logical_Operator_out2993_out1 XOR Logical_Operator_out3057_out1;

  Logical_Operator_out4050_out1 <= Logical_Operator_out2994_out1 XOR Logical_Operator_out3058_out1;

  Logical_Operator_out4051_out1 <= Logical_Operator_out2995_out1 XOR Logical_Operator_out3059_out1;

  Logical_Operator_out4052_out1 <= Logical_Operator_out2996_out1 XOR Logical_Operator_out3060_out1;

  Logical_Operator_out4053_out1 <= Logical_Operator_out2997_out1 XOR Logical_Operator_out3061_out1;

  Logical_Operator_out4054_out1 <= Logical_Operator_out2998_out1 XOR Logical_Operator_out3062_out1;

  Logical_Operator_out4055_out1 <= Logical_Operator_out2999_out1 XOR Logical_Operator_out3063_out1;

  Logical_Operator_out4056_out1 <= Logical_Operator_out3000_out1 XOR Logical_Operator_out3064_out1;

  Logical_Operator_out4057_out1 <= Logical_Operator_out3001_out1 XOR Logical_Operator_out3065_out1;

  Logical_Operator_out4058_out1 <= Logical_Operator_out3002_out1 XOR Logical_Operator_out3066_out1;

  Logical_Operator_out4059_out1 <= Logical_Operator_out3003_out1 XOR Logical_Operator_out3067_out1;

  Logical_Operator_out4060_out1 <= Logical_Operator_out3004_out1 XOR Logical_Operator_out3068_out1;

  Logical_Operator_out4061_out1 <= Logical_Operator_out3005_out1 XOR Logical_Operator_out3069_out1;

  Logical_Operator_out4062_out1 <= Logical_Operator_out3006_out1 XOR Logical_Operator_out3070_out1;

  Logical_Operator_out4063_out1 <= Logical_Operator_out3007_out1 XOR Logical_Operator_out3071_out1;

  Logical_Operator_out4064_out1 <= Logical_Operator_out3008_out1 XOR Logical_Operator_out3072_out1;

  Logical_Operator_out4065_out1 <= Logical_Operator_out2481_out1 XOR Logical_Operator_out2545_out1;

  Logical_Operator_out4066_out1 <= Logical_Operator_out2482_out1 XOR Logical_Operator_out2546_out1;

  Logical_Operator_out4067_out1 <= Logical_Operator_out2483_out1 XOR Logical_Operator_out2547_out1;

  Logical_Operator_out4068_out1 <= Logical_Operator_out2484_out1 XOR Logical_Operator_out2548_out1;

  Logical_Operator_out4069_out1 <= Logical_Operator_out2485_out1 XOR Logical_Operator_out2549_out1;

  Logical_Operator_out4070_out1 <= Logical_Operator_out2486_out1 XOR Logical_Operator_out2550_out1;

  Logical_Operator_out4071_out1 <= Logical_Operator_out2487_out1 XOR Logical_Operator_out2551_out1;

  Logical_Operator_out4072_out1 <= Logical_Operator_out2488_out1 XOR Logical_Operator_out2552_out1;

  Logical_Operator_out4073_out1 <= Logical_Operator_out2489_out1 XOR Logical_Operator_out2553_out1;

  Logical_Operator_out4074_out1 <= Logical_Operator_out2490_out1 XOR Logical_Operator_out2554_out1;

  Logical_Operator_out4075_out1 <= Logical_Operator_out2491_out1 XOR Logical_Operator_out2555_out1;

  Logical_Operator_out4076_out1 <= Logical_Operator_out2492_out1 XOR Logical_Operator_out2556_out1;

  Logical_Operator_out4077_out1 <= Logical_Operator_out2493_out1 XOR Logical_Operator_out2557_out1;

  Logical_Operator_out4078_out1 <= Logical_Operator_out2494_out1 XOR Logical_Operator_out2558_out1;

  Logical_Operator_out4079_out1 <= Logical_Operator_out2495_out1 XOR Logical_Operator_out2559_out1;

  Logical_Operator_out4080_out1 <= Logical_Operator_out2496_out1 XOR Logical_Operator_out2560_out1;

  Logical_Operator_out4081_out1 <= Logical_Operator_out1977_out1 XOR Logical_Operator_out2041_out1;

  Logical_Operator_out4082_out1 <= Logical_Operator_out1978_out1 XOR Logical_Operator_out2042_out1;

  Logical_Operator_out4083_out1 <= Logical_Operator_out1979_out1 XOR Logical_Operator_out2043_out1;

  Logical_Operator_out4084_out1 <= Logical_Operator_out1980_out1 XOR Logical_Operator_out2044_out1;

  Logical_Operator_out4085_out1 <= Logical_Operator_out1981_out1 XOR Logical_Operator_out2045_out1;

  Logical_Operator_out4086_out1 <= Logical_Operator_out1982_out1 XOR Logical_Operator_out2046_out1;

  Logical_Operator_out4087_out1 <= Logical_Operator_out1983_out1 XOR Logical_Operator_out2047_out1;

  Logical_Operator_out4088_out1 <= Logical_Operator_out1984_out1 XOR Logical_Operator_out2048_out1;

  Logical_Operator_out4089_out1 <= Logical_Operator_out1469_out1 XOR Logical_Operator_out1533_out1;

  Logical_Operator_out4090_out1 <= Logical_Operator_out1470_out1 XOR Logical_Operator_out1534_out1;

  Logical_Operator_out4091_out1 <= Logical_Operator_out1471_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out4092_out1 <= Logical_Operator_out1472_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out4093_out1 <= Logical_Operator_out959_out1 XOR Logical_Operator_out1023_out1;

  Logical_Operator_out4094_out1 <= Logical_Operator_out960_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out4095_out1 <= Logical_Operator_out448_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out4096_out1 <= in896 XOR in1024;

  Logical_Operator_out4097_out1 <= Logical_Operator_out3585_out1 XOR Logical_Operator_out3713_out1;

  Logical_Operator_out4098_out1 <= Logical_Operator_out3586_out1 XOR Logical_Operator_out3714_out1;

  Logical_Operator_out4099_out1 <= Logical_Operator_out3587_out1 XOR Logical_Operator_out3715_out1;

  Logical_Operator_out4100_out1 <= Logical_Operator_out3588_out1 XOR Logical_Operator_out3716_out1;

  Logical_Operator_out4101_out1 <= Logical_Operator_out3589_out1 XOR Logical_Operator_out3717_out1;

  Logical_Operator_out4102_out1 <= Logical_Operator_out3590_out1 XOR Logical_Operator_out3718_out1;

  Logical_Operator_out4103_out1 <= Logical_Operator_out3591_out1 XOR Logical_Operator_out3719_out1;

  Logical_Operator_out4104_out1 <= Logical_Operator_out3592_out1 XOR Logical_Operator_out3720_out1;

  Logical_Operator_out4105_out1 <= Logical_Operator_out3593_out1 XOR Logical_Operator_out3721_out1;

  Logical_Operator_out4106_out1 <= Logical_Operator_out3594_out1 XOR Logical_Operator_out3722_out1;

  Logical_Operator_out4107_out1 <= Logical_Operator_out3595_out1 XOR Logical_Operator_out3723_out1;

  Logical_Operator_out4108_out1 <= Logical_Operator_out3596_out1 XOR Logical_Operator_out3724_out1;

  Logical_Operator_out4109_out1 <= Logical_Operator_out3597_out1 XOR Logical_Operator_out3725_out1;

  Logical_Operator_out4110_out1 <= Logical_Operator_out3598_out1 XOR Logical_Operator_out3726_out1;

  Logical_Operator_out4111_out1 <= Logical_Operator_out3599_out1 XOR Logical_Operator_out3727_out1;

  Logical_Operator_out4112_out1 <= Logical_Operator_out3600_out1 XOR Logical_Operator_out3728_out1;

  Logical_Operator_out4113_out1 <= Logical_Operator_out3601_out1 XOR Logical_Operator_out3729_out1;

  Logical_Operator_out4114_out1 <= Logical_Operator_out3602_out1 XOR Logical_Operator_out3730_out1;

  Logical_Operator_out4115_out1 <= Logical_Operator_out3603_out1 XOR Logical_Operator_out3731_out1;

  Logical_Operator_out4116_out1 <= Logical_Operator_out3604_out1 XOR Logical_Operator_out3732_out1;

  Logical_Operator_out4117_out1 <= Logical_Operator_out3605_out1 XOR Logical_Operator_out3733_out1;

  Logical_Operator_out4118_out1 <= Logical_Operator_out3606_out1 XOR Logical_Operator_out3734_out1;

  Logical_Operator_out4119_out1 <= Logical_Operator_out3607_out1 XOR Logical_Operator_out3735_out1;

  Logical_Operator_out4120_out1 <= Logical_Operator_out3608_out1 XOR Logical_Operator_out3736_out1;

  Logical_Operator_out4121_out1 <= Logical_Operator_out3609_out1 XOR Logical_Operator_out3737_out1;

  Logical_Operator_out4122_out1 <= Logical_Operator_out3610_out1 XOR Logical_Operator_out3738_out1;

  Logical_Operator_out4123_out1 <= Logical_Operator_out3611_out1 XOR Logical_Operator_out3739_out1;

  Logical_Operator_out4124_out1 <= Logical_Operator_out3612_out1 XOR Logical_Operator_out3740_out1;

  Logical_Operator_out4125_out1 <= Logical_Operator_out3613_out1 XOR Logical_Operator_out3741_out1;

  Logical_Operator_out4126_out1 <= Logical_Operator_out3614_out1 XOR Logical_Operator_out3742_out1;

  Logical_Operator_out4127_out1 <= Logical_Operator_out3615_out1 XOR Logical_Operator_out3743_out1;

  Logical_Operator_out4128_out1 <= Logical_Operator_out3616_out1 XOR Logical_Operator_out3744_out1;

  Logical_Operator_out4129_out1 <= Logical_Operator_out3617_out1 XOR Logical_Operator_out3745_out1;

  Logical_Operator_out4130_out1 <= Logical_Operator_out3618_out1 XOR Logical_Operator_out3746_out1;

  Logical_Operator_out4131_out1 <= Logical_Operator_out3619_out1 XOR Logical_Operator_out3747_out1;

  Logical_Operator_out4132_out1 <= Logical_Operator_out3620_out1 XOR Logical_Operator_out3748_out1;

  Logical_Operator_out4133_out1 <= Logical_Operator_out3621_out1 XOR Logical_Operator_out3749_out1;

  Logical_Operator_out4134_out1 <= Logical_Operator_out3622_out1 XOR Logical_Operator_out3750_out1;

  Logical_Operator_out4135_out1 <= Logical_Operator_out3623_out1 XOR Logical_Operator_out3751_out1;

  Logical_Operator_out4136_out1 <= Logical_Operator_out3624_out1 XOR Logical_Operator_out3752_out1;

  Logical_Operator_out4137_out1 <= Logical_Operator_out3625_out1 XOR Logical_Operator_out3753_out1;

  Logical_Operator_out4138_out1 <= Logical_Operator_out3626_out1 XOR Logical_Operator_out3754_out1;

  Logical_Operator_out4139_out1 <= Logical_Operator_out3627_out1 XOR Logical_Operator_out3755_out1;

  Logical_Operator_out4140_out1 <= Logical_Operator_out3628_out1 XOR Logical_Operator_out3756_out1;

  Logical_Operator_out4141_out1 <= Logical_Operator_out3629_out1 XOR Logical_Operator_out3757_out1;

  Logical_Operator_out4142_out1 <= Logical_Operator_out3630_out1 XOR Logical_Operator_out3758_out1;

  Logical_Operator_out4143_out1 <= Logical_Operator_out3631_out1 XOR Logical_Operator_out3759_out1;

  Logical_Operator_out4144_out1 <= Logical_Operator_out3632_out1 XOR Logical_Operator_out3760_out1;

  Logical_Operator_out4145_out1 <= Logical_Operator_out3633_out1 XOR Logical_Operator_out3761_out1;

  Logical_Operator_out4146_out1 <= Logical_Operator_out3634_out1 XOR Logical_Operator_out3762_out1;

  Logical_Operator_out4147_out1 <= Logical_Operator_out3635_out1 XOR Logical_Operator_out3763_out1;

  Logical_Operator_out4148_out1 <= Logical_Operator_out3636_out1 XOR Logical_Operator_out3764_out1;

  Logical_Operator_out4149_out1 <= Logical_Operator_out3637_out1 XOR Logical_Operator_out3765_out1;

  Logical_Operator_out4150_out1 <= Logical_Operator_out3638_out1 XOR Logical_Operator_out3766_out1;

  Logical_Operator_out4151_out1 <= Logical_Operator_out3639_out1 XOR Logical_Operator_out3767_out1;

  Logical_Operator_out4152_out1 <= Logical_Operator_out3640_out1 XOR Logical_Operator_out3768_out1;

  Logical_Operator_out4153_out1 <= Logical_Operator_out3641_out1 XOR Logical_Operator_out3769_out1;

  Logical_Operator_out4154_out1 <= Logical_Operator_out3642_out1 XOR Logical_Operator_out3770_out1;

  Logical_Operator_out4155_out1 <= Logical_Operator_out3643_out1 XOR Logical_Operator_out3771_out1;

  Logical_Operator_out4156_out1 <= Logical_Operator_out3644_out1 XOR Logical_Operator_out3772_out1;

  Logical_Operator_out4157_out1 <= Logical_Operator_out3645_out1 XOR Logical_Operator_out3773_out1;

  Logical_Operator_out4158_out1 <= Logical_Operator_out3646_out1 XOR Logical_Operator_out3774_out1;

  Logical_Operator_out4159_out1 <= Logical_Operator_out3647_out1 XOR Logical_Operator_out3775_out1;

  Logical_Operator_out4160_out1 <= Logical_Operator_out3648_out1 XOR Logical_Operator_out3776_out1;

  Logical_Operator_out4161_out1 <= Logical_Operator_out3649_out1 XOR Logical_Operator_out3777_out1;

  Logical_Operator_out4162_out1 <= Logical_Operator_out3650_out1 XOR Logical_Operator_out3778_out1;

  Logical_Operator_out4163_out1 <= Logical_Operator_out3651_out1 XOR Logical_Operator_out3779_out1;

  Logical_Operator_out4164_out1 <= Logical_Operator_out3652_out1 XOR Logical_Operator_out3780_out1;

  Logical_Operator_out4165_out1 <= Logical_Operator_out3653_out1 XOR Logical_Operator_out3781_out1;

  Logical_Operator_out4166_out1 <= Logical_Operator_out3654_out1 XOR Logical_Operator_out3782_out1;

  Logical_Operator_out4167_out1 <= Logical_Operator_out3655_out1 XOR Logical_Operator_out3783_out1;

  Logical_Operator_out4168_out1 <= Logical_Operator_out3656_out1 XOR Logical_Operator_out3784_out1;

  Logical_Operator_out4169_out1 <= Logical_Operator_out3657_out1 XOR Logical_Operator_out3785_out1;

  Logical_Operator_out4170_out1 <= Logical_Operator_out3658_out1 XOR Logical_Operator_out3786_out1;

  Logical_Operator_out4171_out1 <= Logical_Operator_out3659_out1 XOR Logical_Operator_out3787_out1;

  Logical_Operator_out4172_out1 <= Logical_Operator_out3660_out1 XOR Logical_Operator_out3788_out1;

  Logical_Operator_out4173_out1 <= Logical_Operator_out3661_out1 XOR Logical_Operator_out3789_out1;

  Logical_Operator_out4174_out1 <= Logical_Operator_out3662_out1 XOR Logical_Operator_out3790_out1;

  Logical_Operator_out4175_out1 <= Logical_Operator_out3663_out1 XOR Logical_Operator_out3791_out1;

  Logical_Operator_out4176_out1 <= Logical_Operator_out3664_out1 XOR Logical_Operator_out3792_out1;

  Logical_Operator_out4177_out1 <= Logical_Operator_out3665_out1 XOR Logical_Operator_out3793_out1;

  Logical_Operator_out4178_out1 <= Logical_Operator_out3666_out1 XOR Logical_Operator_out3794_out1;

  Logical_Operator_out4179_out1 <= Logical_Operator_out3667_out1 XOR Logical_Operator_out3795_out1;

  Logical_Operator_out4180_out1 <= Logical_Operator_out3668_out1 XOR Logical_Operator_out3796_out1;

  Logical_Operator_out4181_out1 <= Logical_Operator_out3669_out1 XOR Logical_Operator_out3797_out1;

  Logical_Operator_out4182_out1 <= Logical_Operator_out3670_out1 XOR Logical_Operator_out3798_out1;

  Logical_Operator_out4183_out1 <= Logical_Operator_out3671_out1 XOR Logical_Operator_out3799_out1;

  Logical_Operator_out4184_out1 <= Logical_Operator_out3672_out1 XOR Logical_Operator_out3800_out1;

  Logical_Operator_out4185_out1 <= Logical_Operator_out3673_out1 XOR Logical_Operator_out3801_out1;

  Logical_Operator_out4186_out1 <= Logical_Operator_out3674_out1 XOR Logical_Operator_out3802_out1;

  Logical_Operator_out4187_out1 <= Logical_Operator_out3675_out1 XOR Logical_Operator_out3803_out1;

  Logical_Operator_out4188_out1 <= Logical_Operator_out3676_out1 XOR Logical_Operator_out3804_out1;

  Logical_Operator_out4189_out1 <= Logical_Operator_out3677_out1 XOR Logical_Operator_out3805_out1;

  Logical_Operator_out4190_out1 <= Logical_Operator_out3678_out1 XOR Logical_Operator_out3806_out1;

  Logical_Operator_out4191_out1 <= Logical_Operator_out3679_out1 XOR Logical_Operator_out3807_out1;

  Logical_Operator_out4192_out1 <= Logical_Operator_out3680_out1 XOR Logical_Operator_out3808_out1;

  Logical_Operator_out4193_out1 <= Logical_Operator_out3681_out1 XOR Logical_Operator_out3809_out1;

  Logical_Operator_out4194_out1 <= Logical_Operator_out3682_out1 XOR Logical_Operator_out3810_out1;

  Logical_Operator_out4195_out1 <= Logical_Operator_out3683_out1 XOR Logical_Operator_out3811_out1;

  Logical_Operator_out4196_out1 <= Logical_Operator_out3684_out1 XOR Logical_Operator_out3812_out1;

  Logical_Operator_out4197_out1 <= Logical_Operator_out3685_out1 XOR Logical_Operator_out3813_out1;

  Logical_Operator_out4198_out1 <= Logical_Operator_out3686_out1 XOR Logical_Operator_out3814_out1;

  Logical_Operator_out4199_out1 <= Logical_Operator_out3687_out1 XOR Logical_Operator_out3815_out1;

  Logical_Operator_out4200_out1 <= Logical_Operator_out3688_out1 XOR Logical_Operator_out3816_out1;

  Logical_Operator_out4201_out1 <= Logical_Operator_out3689_out1 XOR Logical_Operator_out3817_out1;

  Logical_Operator_out4202_out1 <= Logical_Operator_out3690_out1 XOR Logical_Operator_out3818_out1;

  Logical_Operator_out4203_out1 <= Logical_Operator_out3691_out1 XOR Logical_Operator_out3819_out1;

  Logical_Operator_out4204_out1 <= Logical_Operator_out3692_out1 XOR Logical_Operator_out3820_out1;

  Logical_Operator_out4205_out1 <= Logical_Operator_out3693_out1 XOR Logical_Operator_out3821_out1;

  Logical_Operator_out4206_out1 <= Logical_Operator_out3694_out1 XOR Logical_Operator_out3822_out1;

  Logical_Operator_out4207_out1 <= Logical_Operator_out3695_out1 XOR Logical_Operator_out3823_out1;

  Logical_Operator_out4208_out1 <= Logical_Operator_out3696_out1 XOR Logical_Operator_out3824_out1;

  Logical_Operator_out4209_out1 <= Logical_Operator_out3697_out1 XOR Logical_Operator_out3825_out1;

  Logical_Operator_out4210_out1 <= Logical_Operator_out3698_out1 XOR Logical_Operator_out3826_out1;

  Logical_Operator_out4211_out1 <= Logical_Operator_out3699_out1 XOR Logical_Operator_out3827_out1;

  Logical_Operator_out4212_out1 <= Logical_Operator_out3700_out1 XOR Logical_Operator_out3828_out1;

  Logical_Operator_out4213_out1 <= Logical_Operator_out3701_out1 XOR Logical_Operator_out3829_out1;

  Logical_Operator_out4214_out1 <= Logical_Operator_out3702_out1 XOR Logical_Operator_out3830_out1;

  Logical_Operator_out4215_out1 <= Logical_Operator_out3703_out1 XOR Logical_Operator_out3831_out1;

  Logical_Operator_out4216_out1 <= Logical_Operator_out3704_out1 XOR Logical_Operator_out3832_out1;

  Logical_Operator_out4217_out1 <= Logical_Operator_out3705_out1 XOR Logical_Operator_out3833_out1;

  Logical_Operator_out4218_out1 <= Logical_Operator_out3706_out1 XOR Logical_Operator_out3834_out1;

  Logical_Operator_out4219_out1 <= Logical_Operator_out3707_out1 XOR Logical_Operator_out3835_out1;

  Logical_Operator_out4220_out1 <= Logical_Operator_out3708_out1 XOR Logical_Operator_out3836_out1;

  Logical_Operator_out4221_out1 <= Logical_Operator_out3709_out1 XOR Logical_Operator_out3837_out1;

  Logical_Operator_out4222_out1 <= Logical_Operator_out3710_out1 XOR Logical_Operator_out3838_out1;

  Logical_Operator_out4223_out1 <= Logical_Operator_out3711_out1 XOR Logical_Operator_out3839_out1;

  Logical_Operator_out4224_out1 <= Logical_Operator_out3712_out1 XOR Logical_Operator_out3840_out1;

  Logical_Operator_out4225_out1 <= Logical_Operator_out3137_out1 XOR Logical_Operator_out3265_out1;

  Logical_Operator_out4226_out1 <= Logical_Operator_out3138_out1 XOR Logical_Operator_out3266_out1;

  Logical_Operator_out4227_out1 <= Logical_Operator_out3139_out1 XOR Logical_Operator_out3267_out1;

  Logical_Operator_out4228_out1 <= Logical_Operator_out3140_out1 XOR Logical_Operator_out3268_out1;

  Logical_Operator_out4229_out1 <= Logical_Operator_out3141_out1 XOR Logical_Operator_out3269_out1;

  Logical_Operator_out4230_out1 <= Logical_Operator_out3142_out1 XOR Logical_Operator_out3270_out1;

  Logical_Operator_out4231_out1 <= Logical_Operator_out3143_out1 XOR Logical_Operator_out3271_out1;

  Logical_Operator_out4232_out1 <= Logical_Operator_out3144_out1 XOR Logical_Operator_out3272_out1;

  Logical_Operator_out4233_out1 <= Logical_Operator_out3145_out1 XOR Logical_Operator_out3273_out1;

  Logical_Operator_out4234_out1 <= Logical_Operator_out3146_out1 XOR Logical_Operator_out3274_out1;

  Logical_Operator_out4235_out1 <= Logical_Operator_out3147_out1 XOR Logical_Operator_out3275_out1;

  Logical_Operator_out4236_out1 <= Logical_Operator_out3148_out1 XOR Logical_Operator_out3276_out1;

  Logical_Operator_out4237_out1 <= Logical_Operator_out3149_out1 XOR Logical_Operator_out3277_out1;

  Logical_Operator_out4238_out1 <= Logical_Operator_out3150_out1 XOR Logical_Operator_out3278_out1;

  Logical_Operator_out4239_out1 <= Logical_Operator_out3151_out1 XOR Logical_Operator_out3279_out1;

  Logical_Operator_out4240_out1 <= Logical_Operator_out3152_out1 XOR Logical_Operator_out3280_out1;

  Logical_Operator_out4241_out1 <= Logical_Operator_out3153_out1 XOR Logical_Operator_out3281_out1;

  Logical_Operator_out4242_out1 <= Logical_Operator_out3154_out1 XOR Logical_Operator_out3282_out1;

  Logical_Operator_out4243_out1 <= Logical_Operator_out3155_out1 XOR Logical_Operator_out3283_out1;

  Logical_Operator_out4244_out1 <= Logical_Operator_out3156_out1 XOR Logical_Operator_out3284_out1;

  Logical_Operator_out4245_out1 <= Logical_Operator_out3157_out1 XOR Logical_Operator_out3285_out1;

  Logical_Operator_out4246_out1 <= Logical_Operator_out3158_out1 XOR Logical_Operator_out3286_out1;

  Logical_Operator_out4247_out1 <= Logical_Operator_out3159_out1 XOR Logical_Operator_out3287_out1;

  Logical_Operator_out4248_out1 <= Logical_Operator_out3160_out1 XOR Logical_Operator_out3288_out1;

  Logical_Operator_out4249_out1 <= Logical_Operator_out3161_out1 XOR Logical_Operator_out3289_out1;

  Logical_Operator_out4250_out1 <= Logical_Operator_out3162_out1 XOR Logical_Operator_out3290_out1;

  Logical_Operator_out4251_out1 <= Logical_Operator_out3163_out1 XOR Logical_Operator_out3291_out1;

  Logical_Operator_out4252_out1 <= Logical_Operator_out3164_out1 XOR Logical_Operator_out3292_out1;

  Logical_Operator_out4253_out1 <= Logical_Operator_out3165_out1 XOR Logical_Operator_out3293_out1;

  Logical_Operator_out4254_out1 <= Logical_Operator_out3166_out1 XOR Logical_Operator_out3294_out1;

  Logical_Operator_out4255_out1 <= Logical_Operator_out3167_out1 XOR Logical_Operator_out3295_out1;

  Logical_Operator_out4256_out1 <= Logical_Operator_out3168_out1 XOR Logical_Operator_out3296_out1;

  Logical_Operator_out4257_out1 <= Logical_Operator_out3169_out1 XOR Logical_Operator_out3297_out1;

  Logical_Operator_out4258_out1 <= Logical_Operator_out3170_out1 XOR Logical_Operator_out3298_out1;

  Logical_Operator_out4259_out1 <= Logical_Operator_out3171_out1 XOR Logical_Operator_out3299_out1;

  Logical_Operator_out4260_out1 <= Logical_Operator_out3172_out1 XOR Logical_Operator_out3300_out1;

  Logical_Operator_out4261_out1 <= Logical_Operator_out3173_out1 XOR Logical_Operator_out3301_out1;

  Logical_Operator_out4262_out1 <= Logical_Operator_out3174_out1 XOR Logical_Operator_out3302_out1;

  Logical_Operator_out4263_out1 <= Logical_Operator_out3175_out1 XOR Logical_Operator_out3303_out1;

  Logical_Operator_out4264_out1 <= Logical_Operator_out3176_out1 XOR Logical_Operator_out3304_out1;

  Logical_Operator_out4265_out1 <= Logical_Operator_out3177_out1 XOR Logical_Operator_out3305_out1;

  Logical_Operator_out4266_out1 <= Logical_Operator_out3178_out1 XOR Logical_Operator_out3306_out1;

  Logical_Operator_out4267_out1 <= Logical_Operator_out3179_out1 XOR Logical_Operator_out3307_out1;

  Logical_Operator_out4268_out1 <= Logical_Operator_out3180_out1 XOR Logical_Operator_out3308_out1;

  Logical_Operator_out4269_out1 <= Logical_Operator_out3181_out1 XOR Logical_Operator_out3309_out1;

  Logical_Operator_out4270_out1 <= Logical_Operator_out3182_out1 XOR Logical_Operator_out3310_out1;

  Logical_Operator_out4271_out1 <= Logical_Operator_out3183_out1 XOR Logical_Operator_out3311_out1;

  Logical_Operator_out4272_out1 <= Logical_Operator_out3184_out1 XOR Logical_Operator_out3312_out1;

  Logical_Operator_out4273_out1 <= Logical_Operator_out3185_out1 XOR Logical_Operator_out3313_out1;

  Logical_Operator_out4274_out1 <= Logical_Operator_out3186_out1 XOR Logical_Operator_out3314_out1;

  Logical_Operator_out4275_out1 <= Logical_Operator_out3187_out1 XOR Logical_Operator_out3315_out1;

  Logical_Operator_out4276_out1 <= Logical_Operator_out3188_out1 XOR Logical_Operator_out3316_out1;

  Logical_Operator_out4277_out1 <= Logical_Operator_out3189_out1 XOR Logical_Operator_out3317_out1;

  Logical_Operator_out4278_out1 <= Logical_Operator_out3190_out1 XOR Logical_Operator_out3318_out1;

  Logical_Operator_out4279_out1 <= Logical_Operator_out3191_out1 XOR Logical_Operator_out3319_out1;

  Logical_Operator_out4280_out1 <= Logical_Operator_out3192_out1 XOR Logical_Operator_out3320_out1;

  Logical_Operator_out4281_out1 <= Logical_Operator_out3193_out1 XOR Logical_Operator_out3321_out1;

  Logical_Operator_out4282_out1 <= Logical_Operator_out3194_out1 XOR Logical_Operator_out3322_out1;

  Logical_Operator_out4283_out1 <= Logical_Operator_out3195_out1 XOR Logical_Operator_out3323_out1;

  Logical_Operator_out4284_out1 <= Logical_Operator_out3196_out1 XOR Logical_Operator_out3324_out1;

  Logical_Operator_out4285_out1 <= Logical_Operator_out3197_out1 XOR Logical_Operator_out3325_out1;

  Logical_Operator_out4286_out1 <= Logical_Operator_out3198_out1 XOR Logical_Operator_out3326_out1;

  Logical_Operator_out4287_out1 <= Logical_Operator_out3199_out1 XOR Logical_Operator_out3327_out1;

  Logical_Operator_out4288_out1 <= Logical_Operator_out3200_out1 XOR Logical_Operator_out3328_out1;

  Logical_Operator_out4289_out1 <= Logical_Operator_out2657_out1 XOR Logical_Operator_out2785_out1;

  Logical_Operator_out4290_out1 <= Logical_Operator_out2658_out1 XOR Logical_Operator_out2786_out1;

  Logical_Operator_out4291_out1 <= Logical_Operator_out2659_out1 XOR Logical_Operator_out2787_out1;

  Logical_Operator_out4292_out1 <= Logical_Operator_out2660_out1 XOR Logical_Operator_out2788_out1;

  Logical_Operator_out4293_out1 <= Logical_Operator_out2661_out1 XOR Logical_Operator_out2789_out1;

  Logical_Operator_out4294_out1 <= Logical_Operator_out2662_out1 XOR Logical_Operator_out2790_out1;

  Logical_Operator_out4295_out1 <= Logical_Operator_out2663_out1 XOR Logical_Operator_out2791_out1;

  Logical_Operator_out4296_out1 <= Logical_Operator_out2664_out1 XOR Logical_Operator_out2792_out1;

  Logical_Operator_out4297_out1 <= Logical_Operator_out2665_out1 XOR Logical_Operator_out2793_out1;

  Logical_Operator_out4298_out1 <= Logical_Operator_out2666_out1 XOR Logical_Operator_out2794_out1;

  Logical_Operator_out4299_out1 <= Logical_Operator_out2667_out1 XOR Logical_Operator_out2795_out1;

  Logical_Operator_out4300_out1 <= Logical_Operator_out2668_out1 XOR Logical_Operator_out2796_out1;

  Logical_Operator_out4301_out1 <= Logical_Operator_out2669_out1 XOR Logical_Operator_out2797_out1;

  Logical_Operator_out4302_out1 <= Logical_Operator_out2670_out1 XOR Logical_Operator_out2798_out1;

  Logical_Operator_out4303_out1 <= Logical_Operator_out2671_out1 XOR Logical_Operator_out2799_out1;

  Logical_Operator_out4304_out1 <= Logical_Operator_out2672_out1 XOR Logical_Operator_out2800_out1;

  Logical_Operator_out4305_out1 <= Logical_Operator_out2673_out1 XOR Logical_Operator_out2801_out1;

  Logical_Operator_out4306_out1 <= Logical_Operator_out2674_out1 XOR Logical_Operator_out2802_out1;

  Logical_Operator_out4307_out1 <= Logical_Operator_out2675_out1 XOR Logical_Operator_out2803_out1;

  Logical_Operator_out4308_out1 <= Logical_Operator_out2676_out1 XOR Logical_Operator_out2804_out1;

  Logical_Operator_out4309_out1 <= Logical_Operator_out2677_out1 XOR Logical_Operator_out2805_out1;

  Logical_Operator_out4310_out1 <= Logical_Operator_out2678_out1 XOR Logical_Operator_out2806_out1;

  Logical_Operator_out4311_out1 <= Logical_Operator_out2679_out1 XOR Logical_Operator_out2807_out1;

  Logical_Operator_out4312_out1 <= Logical_Operator_out2680_out1 XOR Logical_Operator_out2808_out1;

  Logical_Operator_out4313_out1 <= Logical_Operator_out2681_out1 XOR Logical_Operator_out2809_out1;

  Logical_Operator_out4314_out1 <= Logical_Operator_out2682_out1 XOR Logical_Operator_out2810_out1;

  Logical_Operator_out4315_out1 <= Logical_Operator_out2683_out1 XOR Logical_Operator_out2811_out1;

  Logical_Operator_out4316_out1 <= Logical_Operator_out2684_out1 XOR Logical_Operator_out2812_out1;

  Logical_Operator_out4317_out1 <= Logical_Operator_out2685_out1 XOR Logical_Operator_out2813_out1;

  Logical_Operator_out4318_out1 <= Logical_Operator_out2686_out1 XOR Logical_Operator_out2814_out1;

  Logical_Operator_out4319_out1 <= Logical_Operator_out2687_out1 XOR Logical_Operator_out2815_out1;

  Logical_Operator_out4320_out1 <= Logical_Operator_out2688_out1 XOR Logical_Operator_out2816_out1;

  Logical_Operator_out4321_out1 <= Logical_Operator_out2161_out1 XOR Logical_Operator_out2289_out1;

  Logical_Operator_out4322_out1 <= Logical_Operator_out2162_out1 XOR Logical_Operator_out2290_out1;

  Logical_Operator_out4323_out1 <= Logical_Operator_out2163_out1 XOR Logical_Operator_out2291_out1;

  Logical_Operator_out4324_out1 <= Logical_Operator_out2164_out1 XOR Logical_Operator_out2292_out1;

  Logical_Operator_out4325_out1 <= Logical_Operator_out2165_out1 XOR Logical_Operator_out2293_out1;

  Logical_Operator_out4326_out1 <= Logical_Operator_out2166_out1 XOR Logical_Operator_out2294_out1;

  Logical_Operator_out4327_out1 <= Logical_Operator_out2167_out1 XOR Logical_Operator_out2295_out1;

  Logical_Operator_out4328_out1 <= Logical_Operator_out2168_out1 XOR Logical_Operator_out2296_out1;

  Logical_Operator_out4329_out1 <= Logical_Operator_out2169_out1 XOR Logical_Operator_out2297_out1;

  Logical_Operator_out4330_out1 <= Logical_Operator_out2170_out1 XOR Logical_Operator_out2298_out1;

  Logical_Operator_out4331_out1 <= Logical_Operator_out2171_out1 XOR Logical_Operator_out2299_out1;

  Logical_Operator_out4332_out1 <= Logical_Operator_out2172_out1 XOR Logical_Operator_out2300_out1;

  Logical_Operator_out4333_out1 <= Logical_Operator_out2173_out1 XOR Logical_Operator_out2301_out1;

  Logical_Operator_out4334_out1 <= Logical_Operator_out2174_out1 XOR Logical_Operator_out2302_out1;

  Logical_Operator_out4335_out1 <= Logical_Operator_out2175_out1 XOR Logical_Operator_out2303_out1;

  Logical_Operator_out4336_out1 <= Logical_Operator_out2176_out1 XOR Logical_Operator_out2304_out1;

  Logical_Operator_out4337_out1 <= Logical_Operator_out1657_out1 XOR Logical_Operator_out1785_out1;

  Logical_Operator_out4338_out1 <= Logical_Operator_out1658_out1 XOR Logical_Operator_out1786_out1;

  Logical_Operator_out4339_out1 <= Logical_Operator_out1659_out1 XOR Logical_Operator_out1787_out1;

  Logical_Operator_out4340_out1 <= Logical_Operator_out1660_out1 XOR Logical_Operator_out1788_out1;

  Logical_Operator_out4341_out1 <= Logical_Operator_out1661_out1 XOR Logical_Operator_out1789_out1;

  Logical_Operator_out4342_out1 <= Logical_Operator_out1662_out1 XOR Logical_Operator_out1790_out1;

  Logical_Operator_out4343_out1 <= Logical_Operator_out1663_out1 XOR Logical_Operator_out1791_out1;

  Logical_Operator_out4344_out1 <= Logical_Operator_out1664_out1 XOR Logical_Operator_out1792_out1;

  Logical_Operator_out4345_out1 <= Logical_Operator_out1149_out1 XOR Logical_Operator_out1277_out1;

  Logical_Operator_out4346_out1 <= Logical_Operator_out1150_out1 XOR Logical_Operator_out1278_out1;

  Logical_Operator_out4347_out1 <= Logical_Operator_out1151_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out4348_out1 <= Logical_Operator_out1152_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out4349_out1 <= Logical_Operator_out639_out1 XOR Logical_Operator_out767_out1;

  Logical_Operator_out4350_out1 <= Logical_Operator_out640_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out4351_out1 <= Logical_Operator_out128_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out4352_out1 <= in256 XOR in512;

  Logical_Operator_out4353_out1 <= Logical_Operator_out3841_out1 XOR Logical_Operator_out3969_out1;

  Logical_Operator_out4354_out1 <= Logical_Operator_out3842_out1 XOR Logical_Operator_out3970_out1;

  Logical_Operator_out4355_out1 <= Logical_Operator_out3843_out1 XOR Logical_Operator_out3971_out1;

  Logical_Operator_out4356_out1 <= Logical_Operator_out3844_out1 XOR Logical_Operator_out3972_out1;

  Logical_Operator_out4357_out1 <= Logical_Operator_out3845_out1 XOR Logical_Operator_out3973_out1;

  Logical_Operator_out4358_out1 <= Logical_Operator_out3846_out1 XOR Logical_Operator_out3974_out1;

  Logical_Operator_out4359_out1 <= Logical_Operator_out3847_out1 XOR Logical_Operator_out3975_out1;

  Logical_Operator_out4360_out1 <= Logical_Operator_out3848_out1 XOR Logical_Operator_out3976_out1;

  Logical_Operator_out4361_out1 <= Logical_Operator_out3849_out1 XOR Logical_Operator_out3977_out1;

  Logical_Operator_out4362_out1 <= Logical_Operator_out3850_out1 XOR Logical_Operator_out3978_out1;

  Logical_Operator_out4363_out1 <= Logical_Operator_out3851_out1 XOR Logical_Operator_out3979_out1;

  Logical_Operator_out4364_out1 <= Logical_Operator_out3852_out1 XOR Logical_Operator_out3980_out1;

  Logical_Operator_out4365_out1 <= Logical_Operator_out3853_out1 XOR Logical_Operator_out3981_out1;

  Logical_Operator_out4366_out1 <= Logical_Operator_out3854_out1 XOR Logical_Operator_out3982_out1;

  Logical_Operator_out4367_out1 <= Logical_Operator_out3855_out1 XOR Logical_Operator_out3983_out1;

  Logical_Operator_out4368_out1 <= Logical_Operator_out3856_out1 XOR Logical_Operator_out3984_out1;

  Logical_Operator_out4369_out1 <= Logical_Operator_out3857_out1 XOR Logical_Operator_out3985_out1;

  Logical_Operator_out4370_out1 <= Logical_Operator_out3858_out1 XOR Logical_Operator_out3986_out1;

  Logical_Operator_out4371_out1 <= Logical_Operator_out3859_out1 XOR Logical_Operator_out3987_out1;

  Logical_Operator_out4372_out1 <= Logical_Operator_out3860_out1 XOR Logical_Operator_out3988_out1;

  Logical_Operator_out4373_out1 <= Logical_Operator_out3861_out1 XOR Logical_Operator_out3989_out1;

  Logical_Operator_out4374_out1 <= Logical_Operator_out3862_out1 XOR Logical_Operator_out3990_out1;

  Logical_Operator_out4375_out1 <= Logical_Operator_out3863_out1 XOR Logical_Operator_out3991_out1;

  Logical_Operator_out4376_out1 <= Logical_Operator_out3864_out1 XOR Logical_Operator_out3992_out1;

  Logical_Operator_out4377_out1 <= Logical_Operator_out3865_out1 XOR Logical_Operator_out3993_out1;

  Logical_Operator_out4378_out1 <= Logical_Operator_out3866_out1 XOR Logical_Operator_out3994_out1;

  Logical_Operator_out4379_out1 <= Logical_Operator_out3867_out1 XOR Logical_Operator_out3995_out1;

  Logical_Operator_out4380_out1 <= Logical_Operator_out3868_out1 XOR Logical_Operator_out3996_out1;

  Logical_Operator_out4381_out1 <= Logical_Operator_out3869_out1 XOR Logical_Operator_out3997_out1;

  Logical_Operator_out4382_out1 <= Logical_Operator_out3870_out1 XOR Logical_Operator_out3998_out1;

  Logical_Operator_out4383_out1 <= Logical_Operator_out3871_out1 XOR Logical_Operator_out3999_out1;

  Logical_Operator_out4384_out1 <= Logical_Operator_out3872_out1 XOR Logical_Operator_out4000_out1;

  Logical_Operator_out4385_out1 <= Logical_Operator_out3873_out1 XOR Logical_Operator_out4001_out1;

  Logical_Operator_out4386_out1 <= Logical_Operator_out3874_out1 XOR Logical_Operator_out4002_out1;

  Logical_Operator_out4387_out1 <= Logical_Operator_out3875_out1 XOR Logical_Operator_out4003_out1;

  Logical_Operator_out4388_out1 <= Logical_Operator_out3876_out1 XOR Logical_Operator_out4004_out1;

  Logical_Operator_out4389_out1 <= Logical_Operator_out3877_out1 XOR Logical_Operator_out4005_out1;

  Logical_Operator_out4390_out1 <= Logical_Operator_out3878_out1 XOR Logical_Operator_out4006_out1;

  Logical_Operator_out4391_out1 <= Logical_Operator_out3879_out1 XOR Logical_Operator_out4007_out1;

  Logical_Operator_out4392_out1 <= Logical_Operator_out3880_out1 XOR Logical_Operator_out4008_out1;

  Logical_Operator_out4393_out1 <= Logical_Operator_out3881_out1 XOR Logical_Operator_out4009_out1;

  Logical_Operator_out4394_out1 <= Logical_Operator_out3882_out1 XOR Logical_Operator_out4010_out1;

  Logical_Operator_out4395_out1 <= Logical_Operator_out3883_out1 XOR Logical_Operator_out4011_out1;

  Logical_Operator_out4396_out1 <= Logical_Operator_out3884_out1 XOR Logical_Operator_out4012_out1;

  Logical_Operator_out4397_out1 <= Logical_Operator_out3885_out1 XOR Logical_Operator_out4013_out1;

  Logical_Operator_out4398_out1 <= Logical_Operator_out3886_out1 XOR Logical_Operator_out4014_out1;

  Logical_Operator_out4399_out1 <= Logical_Operator_out3887_out1 XOR Logical_Operator_out4015_out1;

  Logical_Operator_out4400_out1 <= Logical_Operator_out3888_out1 XOR Logical_Operator_out4016_out1;

  Logical_Operator_out4401_out1 <= Logical_Operator_out3889_out1 XOR Logical_Operator_out4017_out1;

  Logical_Operator_out4402_out1 <= Logical_Operator_out3890_out1 XOR Logical_Operator_out4018_out1;

  Logical_Operator_out4403_out1 <= Logical_Operator_out3891_out1 XOR Logical_Operator_out4019_out1;

  Logical_Operator_out4404_out1 <= Logical_Operator_out3892_out1 XOR Logical_Operator_out4020_out1;

  Logical_Operator_out4405_out1 <= Logical_Operator_out3893_out1 XOR Logical_Operator_out4021_out1;

  Logical_Operator_out4406_out1 <= Logical_Operator_out3894_out1 XOR Logical_Operator_out4022_out1;

  Logical_Operator_out4407_out1 <= Logical_Operator_out3895_out1 XOR Logical_Operator_out4023_out1;

  Logical_Operator_out4408_out1 <= Logical_Operator_out3896_out1 XOR Logical_Operator_out4024_out1;

  Logical_Operator_out4409_out1 <= Logical_Operator_out3897_out1 XOR Logical_Operator_out4025_out1;

  Logical_Operator_out4410_out1 <= Logical_Operator_out3898_out1 XOR Logical_Operator_out4026_out1;

  Logical_Operator_out4411_out1 <= Logical_Operator_out3899_out1 XOR Logical_Operator_out4027_out1;

  Logical_Operator_out4412_out1 <= Logical_Operator_out3900_out1 XOR Logical_Operator_out4028_out1;

  Logical_Operator_out4413_out1 <= Logical_Operator_out3901_out1 XOR Logical_Operator_out4029_out1;

  Logical_Operator_out4414_out1 <= Logical_Operator_out3902_out1 XOR Logical_Operator_out4030_out1;

  Logical_Operator_out4415_out1 <= Logical_Operator_out3903_out1 XOR Logical_Operator_out4031_out1;

  Logical_Operator_out4416_out1 <= Logical_Operator_out3904_out1 XOR Logical_Operator_out4032_out1;

  Logical_Operator_out4417_out1 <= Logical_Operator_out3905_out1 XOR Logical_Operator_out4033_out1;

  Logical_Operator_out4418_out1 <= Logical_Operator_out3906_out1 XOR Logical_Operator_out4034_out1;

  Logical_Operator_out4419_out1 <= Logical_Operator_out3907_out1 XOR Logical_Operator_out4035_out1;

  Logical_Operator_out4420_out1 <= Logical_Operator_out3908_out1 XOR Logical_Operator_out4036_out1;

  Logical_Operator_out4421_out1 <= Logical_Operator_out3909_out1 XOR Logical_Operator_out4037_out1;

  Logical_Operator_out4422_out1 <= Logical_Operator_out3910_out1 XOR Logical_Operator_out4038_out1;

  Logical_Operator_out4423_out1 <= Logical_Operator_out3911_out1 XOR Logical_Operator_out4039_out1;

  Logical_Operator_out4424_out1 <= Logical_Operator_out3912_out1 XOR Logical_Operator_out4040_out1;

  Logical_Operator_out4425_out1 <= Logical_Operator_out3913_out1 XOR Logical_Operator_out4041_out1;

  Logical_Operator_out4426_out1 <= Logical_Operator_out3914_out1 XOR Logical_Operator_out4042_out1;

  Logical_Operator_out4427_out1 <= Logical_Operator_out3915_out1 XOR Logical_Operator_out4043_out1;

  Logical_Operator_out4428_out1 <= Logical_Operator_out3916_out1 XOR Logical_Operator_out4044_out1;

  Logical_Operator_out4429_out1 <= Logical_Operator_out3917_out1 XOR Logical_Operator_out4045_out1;

  Logical_Operator_out4430_out1 <= Logical_Operator_out3918_out1 XOR Logical_Operator_out4046_out1;

  Logical_Operator_out4431_out1 <= Logical_Operator_out3919_out1 XOR Logical_Operator_out4047_out1;

  Logical_Operator_out4432_out1 <= Logical_Operator_out3920_out1 XOR Logical_Operator_out4048_out1;

  Logical_Operator_out4433_out1 <= Logical_Operator_out3921_out1 XOR Logical_Operator_out4049_out1;

  Logical_Operator_out4434_out1 <= Logical_Operator_out3922_out1 XOR Logical_Operator_out4050_out1;

  Logical_Operator_out4435_out1 <= Logical_Operator_out3923_out1 XOR Logical_Operator_out4051_out1;

  Logical_Operator_out4436_out1 <= Logical_Operator_out3924_out1 XOR Logical_Operator_out4052_out1;

  Logical_Operator_out4437_out1 <= Logical_Operator_out3925_out1 XOR Logical_Operator_out4053_out1;

  Logical_Operator_out4438_out1 <= Logical_Operator_out3926_out1 XOR Logical_Operator_out4054_out1;

  Logical_Operator_out4439_out1 <= Logical_Operator_out3927_out1 XOR Logical_Operator_out4055_out1;

  Logical_Operator_out4440_out1 <= Logical_Operator_out3928_out1 XOR Logical_Operator_out4056_out1;

  Logical_Operator_out4441_out1 <= Logical_Operator_out3929_out1 XOR Logical_Operator_out4057_out1;

  Logical_Operator_out4442_out1 <= Logical_Operator_out3930_out1 XOR Logical_Operator_out4058_out1;

  Logical_Operator_out4443_out1 <= Logical_Operator_out3931_out1 XOR Logical_Operator_out4059_out1;

  Logical_Operator_out4444_out1 <= Logical_Operator_out3932_out1 XOR Logical_Operator_out4060_out1;

  Logical_Operator_out4445_out1 <= Logical_Operator_out3933_out1 XOR Logical_Operator_out4061_out1;

  Logical_Operator_out4446_out1 <= Logical_Operator_out3934_out1 XOR Logical_Operator_out4062_out1;

  Logical_Operator_out4447_out1 <= Logical_Operator_out3935_out1 XOR Logical_Operator_out4063_out1;

  Logical_Operator_out4448_out1 <= Logical_Operator_out3936_out1 XOR Logical_Operator_out4064_out1;

  Logical_Operator_out4449_out1 <= Logical_Operator_out3937_out1 XOR Logical_Operator_out4065_out1;

  Logical_Operator_out4450_out1 <= Logical_Operator_out3938_out1 XOR Logical_Operator_out4066_out1;

  Logical_Operator_out4451_out1 <= Logical_Operator_out3939_out1 XOR Logical_Operator_out4067_out1;

  Logical_Operator_out4452_out1 <= Logical_Operator_out3940_out1 XOR Logical_Operator_out4068_out1;

  Logical_Operator_out4453_out1 <= Logical_Operator_out3941_out1 XOR Logical_Operator_out4069_out1;

  Logical_Operator_out4454_out1 <= Logical_Operator_out3942_out1 XOR Logical_Operator_out4070_out1;

  Logical_Operator_out4455_out1 <= Logical_Operator_out3943_out1 XOR Logical_Operator_out4071_out1;

  Logical_Operator_out4456_out1 <= Logical_Operator_out3944_out1 XOR Logical_Operator_out4072_out1;

  Logical_Operator_out4457_out1 <= Logical_Operator_out3945_out1 XOR Logical_Operator_out4073_out1;

  Logical_Operator_out4458_out1 <= Logical_Operator_out3946_out1 XOR Logical_Operator_out4074_out1;

  Logical_Operator_out4459_out1 <= Logical_Operator_out3947_out1 XOR Logical_Operator_out4075_out1;

  Logical_Operator_out4460_out1 <= Logical_Operator_out3948_out1 XOR Logical_Operator_out4076_out1;

  Logical_Operator_out4461_out1 <= Logical_Operator_out3949_out1 XOR Logical_Operator_out4077_out1;

  Logical_Operator_out4462_out1 <= Logical_Operator_out3950_out1 XOR Logical_Operator_out4078_out1;

  Logical_Operator_out4463_out1 <= Logical_Operator_out3951_out1 XOR Logical_Operator_out4079_out1;

  Logical_Operator_out4464_out1 <= Logical_Operator_out3952_out1 XOR Logical_Operator_out4080_out1;

  Logical_Operator_out4465_out1 <= Logical_Operator_out3953_out1 XOR Logical_Operator_out4081_out1;

  Logical_Operator_out4466_out1 <= Logical_Operator_out3954_out1 XOR Logical_Operator_out4082_out1;

  Logical_Operator_out4467_out1 <= Logical_Operator_out3955_out1 XOR Logical_Operator_out4083_out1;

  Logical_Operator_out4468_out1 <= Logical_Operator_out3956_out1 XOR Logical_Operator_out4084_out1;

  Logical_Operator_out4469_out1 <= Logical_Operator_out3957_out1 XOR Logical_Operator_out4085_out1;

  Logical_Operator_out4470_out1 <= Logical_Operator_out3958_out1 XOR Logical_Operator_out4086_out1;

  Logical_Operator_out4471_out1 <= Logical_Operator_out3959_out1 XOR Logical_Operator_out4087_out1;

  Logical_Operator_out4472_out1 <= Logical_Operator_out3960_out1 XOR Logical_Operator_out4088_out1;

  Logical_Operator_out4473_out1 <= Logical_Operator_out3961_out1 XOR Logical_Operator_out4089_out1;

  Logical_Operator_out4474_out1 <= Logical_Operator_out3962_out1 XOR Logical_Operator_out4090_out1;

  Logical_Operator_out4475_out1 <= Logical_Operator_out3963_out1 XOR Logical_Operator_out4091_out1;

  Logical_Operator_out4476_out1 <= Logical_Operator_out3964_out1 XOR Logical_Operator_out4092_out1;

  Logical_Operator_out4477_out1 <= Logical_Operator_out3965_out1 XOR Logical_Operator_out4093_out1;

  Logical_Operator_out4478_out1 <= Logical_Operator_out3966_out1 XOR Logical_Operator_out4094_out1;

  Logical_Operator_out4479_out1 <= Logical_Operator_out3967_out1 XOR Logical_Operator_out4095_out1;

  Logical_Operator_out4480_out1 <= Logical_Operator_out3968_out1 XOR Logical_Operator_out4096_out1;

  Logical_Operator_out4481_out1 <= Logical_Operator_out3393_out1 XOR Logical_Operator_out3521_out1;

  Logical_Operator_out4482_out1 <= Logical_Operator_out3394_out1 XOR Logical_Operator_out3522_out1;

  Logical_Operator_out4483_out1 <= Logical_Operator_out3395_out1 XOR Logical_Operator_out3523_out1;

  Logical_Operator_out4484_out1 <= Logical_Operator_out3396_out1 XOR Logical_Operator_out3524_out1;

  Logical_Operator_out4485_out1 <= Logical_Operator_out3397_out1 XOR Logical_Operator_out3525_out1;

  Logical_Operator_out4486_out1 <= Logical_Operator_out3398_out1 XOR Logical_Operator_out3526_out1;

  Logical_Operator_out4487_out1 <= Logical_Operator_out3399_out1 XOR Logical_Operator_out3527_out1;

  Logical_Operator_out4488_out1 <= Logical_Operator_out3400_out1 XOR Logical_Operator_out3528_out1;

  Logical_Operator_out4489_out1 <= Logical_Operator_out3401_out1 XOR Logical_Operator_out3529_out1;

  Logical_Operator_out4490_out1 <= Logical_Operator_out3402_out1 XOR Logical_Operator_out3530_out1;

  Logical_Operator_out4491_out1 <= Logical_Operator_out3403_out1 XOR Logical_Operator_out3531_out1;

  Logical_Operator_out4492_out1 <= Logical_Operator_out3404_out1 XOR Logical_Operator_out3532_out1;

  Logical_Operator_out4493_out1 <= Logical_Operator_out3405_out1 XOR Logical_Operator_out3533_out1;

  Logical_Operator_out4494_out1 <= Logical_Operator_out3406_out1 XOR Logical_Operator_out3534_out1;

  Logical_Operator_out4495_out1 <= Logical_Operator_out3407_out1 XOR Logical_Operator_out3535_out1;

  Logical_Operator_out4496_out1 <= Logical_Operator_out3408_out1 XOR Logical_Operator_out3536_out1;

  Logical_Operator_out4497_out1 <= Logical_Operator_out3409_out1 XOR Logical_Operator_out3537_out1;

  Logical_Operator_out4498_out1 <= Logical_Operator_out3410_out1 XOR Logical_Operator_out3538_out1;

  Logical_Operator_out4499_out1 <= Logical_Operator_out3411_out1 XOR Logical_Operator_out3539_out1;

  Logical_Operator_out4500_out1 <= Logical_Operator_out3412_out1 XOR Logical_Operator_out3540_out1;

  Logical_Operator_out4501_out1 <= Logical_Operator_out3413_out1 XOR Logical_Operator_out3541_out1;

  Logical_Operator_out4502_out1 <= Logical_Operator_out3414_out1 XOR Logical_Operator_out3542_out1;

  Logical_Operator_out4503_out1 <= Logical_Operator_out3415_out1 XOR Logical_Operator_out3543_out1;

  Logical_Operator_out4504_out1 <= Logical_Operator_out3416_out1 XOR Logical_Operator_out3544_out1;

  Logical_Operator_out4505_out1 <= Logical_Operator_out3417_out1 XOR Logical_Operator_out3545_out1;

  Logical_Operator_out4506_out1 <= Logical_Operator_out3418_out1 XOR Logical_Operator_out3546_out1;

  Logical_Operator_out4507_out1 <= Logical_Operator_out3419_out1 XOR Logical_Operator_out3547_out1;

  Logical_Operator_out4508_out1 <= Logical_Operator_out3420_out1 XOR Logical_Operator_out3548_out1;

  Logical_Operator_out4509_out1 <= Logical_Operator_out3421_out1 XOR Logical_Operator_out3549_out1;

  Logical_Operator_out4510_out1 <= Logical_Operator_out3422_out1 XOR Logical_Operator_out3550_out1;

  Logical_Operator_out4511_out1 <= Logical_Operator_out3423_out1 XOR Logical_Operator_out3551_out1;

  Logical_Operator_out4512_out1 <= Logical_Operator_out3424_out1 XOR Logical_Operator_out3552_out1;

  Logical_Operator_out4513_out1 <= Logical_Operator_out3425_out1 XOR Logical_Operator_out3553_out1;

  Logical_Operator_out4514_out1 <= Logical_Operator_out3426_out1 XOR Logical_Operator_out3554_out1;

  Logical_Operator_out4515_out1 <= Logical_Operator_out3427_out1 XOR Logical_Operator_out3555_out1;

  Logical_Operator_out4516_out1 <= Logical_Operator_out3428_out1 XOR Logical_Operator_out3556_out1;

  Logical_Operator_out4517_out1 <= Logical_Operator_out3429_out1 XOR Logical_Operator_out3557_out1;

  Logical_Operator_out4518_out1 <= Logical_Operator_out3430_out1 XOR Logical_Operator_out3558_out1;

  Logical_Operator_out4519_out1 <= Logical_Operator_out3431_out1 XOR Logical_Operator_out3559_out1;

  Logical_Operator_out4520_out1 <= Logical_Operator_out3432_out1 XOR Logical_Operator_out3560_out1;

  Logical_Operator_out4521_out1 <= Logical_Operator_out3433_out1 XOR Logical_Operator_out3561_out1;

  Logical_Operator_out4522_out1 <= Logical_Operator_out3434_out1 XOR Logical_Operator_out3562_out1;

  Logical_Operator_out4523_out1 <= Logical_Operator_out3435_out1 XOR Logical_Operator_out3563_out1;

  Logical_Operator_out4524_out1 <= Logical_Operator_out3436_out1 XOR Logical_Operator_out3564_out1;

  Logical_Operator_out4525_out1 <= Logical_Operator_out3437_out1 XOR Logical_Operator_out3565_out1;

  Logical_Operator_out4526_out1 <= Logical_Operator_out3438_out1 XOR Logical_Operator_out3566_out1;

  Logical_Operator_out4527_out1 <= Logical_Operator_out3439_out1 XOR Logical_Operator_out3567_out1;

  Logical_Operator_out4528_out1 <= Logical_Operator_out3440_out1 XOR Logical_Operator_out3568_out1;

  Logical_Operator_out4529_out1 <= Logical_Operator_out3441_out1 XOR Logical_Operator_out3569_out1;

  Logical_Operator_out4530_out1 <= Logical_Operator_out3442_out1 XOR Logical_Operator_out3570_out1;

  Logical_Operator_out4531_out1 <= Logical_Operator_out3443_out1 XOR Logical_Operator_out3571_out1;

  Logical_Operator_out4532_out1 <= Logical_Operator_out3444_out1 XOR Logical_Operator_out3572_out1;

  Logical_Operator_out4533_out1 <= Logical_Operator_out3445_out1 XOR Logical_Operator_out3573_out1;

  Logical_Operator_out4534_out1 <= Logical_Operator_out3446_out1 XOR Logical_Operator_out3574_out1;

  Logical_Operator_out4535_out1 <= Logical_Operator_out3447_out1 XOR Logical_Operator_out3575_out1;

  Logical_Operator_out4536_out1 <= Logical_Operator_out3448_out1 XOR Logical_Operator_out3576_out1;

  Logical_Operator_out4537_out1 <= Logical_Operator_out3449_out1 XOR Logical_Operator_out3577_out1;

  Logical_Operator_out4538_out1 <= Logical_Operator_out3450_out1 XOR Logical_Operator_out3578_out1;

  Logical_Operator_out4539_out1 <= Logical_Operator_out3451_out1 XOR Logical_Operator_out3579_out1;

  Logical_Operator_out4540_out1 <= Logical_Operator_out3452_out1 XOR Logical_Operator_out3580_out1;

  Logical_Operator_out4541_out1 <= Logical_Operator_out3453_out1 XOR Logical_Operator_out3581_out1;

  Logical_Operator_out4542_out1 <= Logical_Operator_out3454_out1 XOR Logical_Operator_out3582_out1;

  Logical_Operator_out4543_out1 <= Logical_Operator_out3455_out1 XOR Logical_Operator_out3583_out1;

  Logical_Operator_out4544_out1 <= Logical_Operator_out3456_out1 XOR Logical_Operator_out3584_out1;

  Logical_Operator_out4545_out1 <= Logical_Operator_out2913_out1 XOR Logical_Operator_out3041_out1;

  Logical_Operator_out4546_out1 <= Logical_Operator_out2914_out1 XOR Logical_Operator_out3042_out1;

  Logical_Operator_out4547_out1 <= Logical_Operator_out2915_out1 XOR Logical_Operator_out3043_out1;

  Logical_Operator_out4548_out1 <= Logical_Operator_out2916_out1 XOR Logical_Operator_out3044_out1;

  Logical_Operator_out4549_out1 <= Logical_Operator_out2917_out1 XOR Logical_Operator_out3045_out1;

  Logical_Operator_out4550_out1 <= Logical_Operator_out2918_out1 XOR Logical_Operator_out3046_out1;

  Logical_Operator_out4551_out1 <= Logical_Operator_out2919_out1 XOR Logical_Operator_out3047_out1;

  Logical_Operator_out4552_out1 <= Logical_Operator_out2920_out1 XOR Logical_Operator_out3048_out1;

  Logical_Operator_out4553_out1 <= Logical_Operator_out2921_out1 XOR Logical_Operator_out3049_out1;

  Logical_Operator_out4554_out1 <= Logical_Operator_out2922_out1 XOR Logical_Operator_out3050_out1;

  Logical_Operator_out4555_out1 <= Logical_Operator_out2923_out1 XOR Logical_Operator_out3051_out1;

  Logical_Operator_out4556_out1 <= Logical_Operator_out2924_out1 XOR Logical_Operator_out3052_out1;

  Logical_Operator_out4557_out1 <= Logical_Operator_out2925_out1 XOR Logical_Operator_out3053_out1;

  Logical_Operator_out4558_out1 <= Logical_Operator_out2926_out1 XOR Logical_Operator_out3054_out1;

  Logical_Operator_out4559_out1 <= Logical_Operator_out2927_out1 XOR Logical_Operator_out3055_out1;

  Logical_Operator_out4560_out1 <= Logical_Operator_out2928_out1 XOR Logical_Operator_out3056_out1;

  Logical_Operator_out4561_out1 <= Logical_Operator_out2929_out1 XOR Logical_Operator_out3057_out1;

  Logical_Operator_out4562_out1 <= Logical_Operator_out2930_out1 XOR Logical_Operator_out3058_out1;

  Logical_Operator_out4563_out1 <= Logical_Operator_out2931_out1 XOR Logical_Operator_out3059_out1;

  Logical_Operator_out4564_out1 <= Logical_Operator_out2932_out1 XOR Logical_Operator_out3060_out1;

  Logical_Operator_out4565_out1 <= Logical_Operator_out2933_out1 XOR Logical_Operator_out3061_out1;

  Logical_Operator_out4566_out1 <= Logical_Operator_out2934_out1 XOR Logical_Operator_out3062_out1;

  Logical_Operator_out4567_out1 <= Logical_Operator_out2935_out1 XOR Logical_Operator_out3063_out1;

  Logical_Operator_out4568_out1 <= Logical_Operator_out2936_out1 XOR Logical_Operator_out3064_out1;

  Logical_Operator_out4569_out1 <= Logical_Operator_out2937_out1 XOR Logical_Operator_out3065_out1;

  Logical_Operator_out4570_out1 <= Logical_Operator_out2938_out1 XOR Logical_Operator_out3066_out1;

  Logical_Operator_out4571_out1 <= Logical_Operator_out2939_out1 XOR Logical_Operator_out3067_out1;

  Logical_Operator_out4572_out1 <= Logical_Operator_out2940_out1 XOR Logical_Operator_out3068_out1;

  Logical_Operator_out4573_out1 <= Logical_Operator_out2941_out1 XOR Logical_Operator_out3069_out1;

  Logical_Operator_out4574_out1 <= Logical_Operator_out2942_out1 XOR Logical_Operator_out3070_out1;

  Logical_Operator_out4575_out1 <= Logical_Operator_out2943_out1 XOR Logical_Operator_out3071_out1;

  Logical_Operator_out4576_out1 <= Logical_Operator_out2944_out1 XOR Logical_Operator_out3072_out1;

  Logical_Operator_out4577_out1 <= Logical_Operator_out2417_out1 XOR Logical_Operator_out2545_out1;

  Logical_Operator_out4578_out1 <= Logical_Operator_out2418_out1 XOR Logical_Operator_out2546_out1;

  Logical_Operator_out4579_out1 <= Logical_Operator_out2419_out1 XOR Logical_Operator_out2547_out1;

  Logical_Operator_out4580_out1 <= Logical_Operator_out2420_out1 XOR Logical_Operator_out2548_out1;

  Logical_Operator_out4581_out1 <= Logical_Operator_out2421_out1 XOR Logical_Operator_out2549_out1;

  Logical_Operator_out4582_out1 <= Logical_Operator_out2422_out1 XOR Logical_Operator_out2550_out1;

  Logical_Operator_out4583_out1 <= Logical_Operator_out2423_out1 XOR Logical_Operator_out2551_out1;

  Logical_Operator_out4584_out1 <= Logical_Operator_out2424_out1 XOR Logical_Operator_out2552_out1;

  Logical_Operator_out4585_out1 <= Logical_Operator_out2425_out1 XOR Logical_Operator_out2553_out1;

  Logical_Operator_out4586_out1 <= Logical_Operator_out2426_out1 XOR Logical_Operator_out2554_out1;

  Logical_Operator_out4587_out1 <= Logical_Operator_out2427_out1 XOR Logical_Operator_out2555_out1;

  Logical_Operator_out4588_out1 <= Logical_Operator_out2428_out1 XOR Logical_Operator_out2556_out1;

  Logical_Operator_out4589_out1 <= Logical_Operator_out2429_out1 XOR Logical_Operator_out2557_out1;

  Logical_Operator_out4590_out1 <= Logical_Operator_out2430_out1 XOR Logical_Operator_out2558_out1;

  Logical_Operator_out4591_out1 <= Logical_Operator_out2431_out1 XOR Logical_Operator_out2559_out1;

  Logical_Operator_out4592_out1 <= Logical_Operator_out2432_out1 XOR Logical_Operator_out2560_out1;

  Logical_Operator_out4593_out1 <= Logical_Operator_out1913_out1 XOR Logical_Operator_out2041_out1;

  Logical_Operator_out4594_out1 <= Logical_Operator_out1914_out1 XOR Logical_Operator_out2042_out1;

  Logical_Operator_out4595_out1 <= Logical_Operator_out1915_out1 XOR Logical_Operator_out2043_out1;

  Logical_Operator_out4596_out1 <= Logical_Operator_out1916_out1 XOR Logical_Operator_out2044_out1;

  Logical_Operator_out4597_out1 <= Logical_Operator_out1917_out1 XOR Logical_Operator_out2045_out1;

  Logical_Operator_out4598_out1 <= Logical_Operator_out1918_out1 XOR Logical_Operator_out2046_out1;

  Logical_Operator_out4599_out1 <= Logical_Operator_out1919_out1 XOR Logical_Operator_out2047_out1;

  Logical_Operator_out4600_out1 <= Logical_Operator_out1920_out1 XOR Logical_Operator_out2048_out1;

  Logical_Operator_out4601_out1 <= Logical_Operator_out1405_out1 XOR Logical_Operator_out1533_out1;

  Logical_Operator_out4602_out1 <= Logical_Operator_out1406_out1 XOR Logical_Operator_out1534_out1;

  Logical_Operator_out4603_out1 <= Logical_Operator_out1407_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out4604_out1 <= Logical_Operator_out1408_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out4605_out1 <= Logical_Operator_out895_out1 XOR Logical_Operator_out1023_out1;

  Logical_Operator_out4606_out1 <= Logical_Operator_out896_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out4607_out1 <= Logical_Operator_out384_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out4608_out1 <= in768 XOR in1024;

  Logical_Operator_out4609_out1 <= Logical_Operator_out4097_out1 XOR Logical_Operator_out4353_out1;

  Logical_Operator_out4610_out1 <= Logical_Operator_out4098_out1 XOR Logical_Operator_out4354_out1;

  Logical_Operator_out4611_out1 <= Logical_Operator_out4099_out1 XOR Logical_Operator_out4355_out1;

  Logical_Operator_out4612_out1 <= Logical_Operator_out4100_out1 XOR Logical_Operator_out4356_out1;

  Logical_Operator_out4613_out1 <= Logical_Operator_out4101_out1 XOR Logical_Operator_out4357_out1;

  Logical_Operator_out4614_out1 <= Logical_Operator_out4102_out1 XOR Logical_Operator_out4358_out1;

  Logical_Operator_out4615_out1 <= Logical_Operator_out4103_out1 XOR Logical_Operator_out4359_out1;

  Logical_Operator_out4616_out1 <= Logical_Operator_out4104_out1 XOR Logical_Operator_out4360_out1;

  Logical_Operator_out4617_out1 <= Logical_Operator_out4105_out1 XOR Logical_Operator_out4361_out1;

  Logical_Operator_out4618_out1 <= Logical_Operator_out4106_out1 XOR Logical_Operator_out4362_out1;

  Logical_Operator_out4619_out1 <= Logical_Operator_out4107_out1 XOR Logical_Operator_out4363_out1;

  Logical_Operator_out4620_out1 <= Logical_Operator_out4108_out1 XOR Logical_Operator_out4364_out1;

  Logical_Operator_out4621_out1 <= Logical_Operator_out4109_out1 XOR Logical_Operator_out4365_out1;

  Logical_Operator_out4622_out1 <= Logical_Operator_out4110_out1 XOR Logical_Operator_out4366_out1;

  Logical_Operator_out4623_out1 <= Logical_Operator_out4111_out1 XOR Logical_Operator_out4367_out1;

  Logical_Operator_out4624_out1 <= Logical_Operator_out4112_out1 XOR Logical_Operator_out4368_out1;

  Logical_Operator_out4625_out1 <= Logical_Operator_out4113_out1 XOR Logical_Operator_out4369_out1;

  Logical_Operator_out4626_out1 <= Logical_Operator_out4114_out1 XOR Logical_Operator_out4370_out1;

  Logical_Operator_out4627_out1 <= Logical_Operator_out4115_out1 XOR Logical_Operator_out4371_out1;

  Logical_Operator_out4628_out1 <= Logical_Operator_out4116_out1 XOR Logical_Operator_out4372_out1;

  Logical_Operator_out4629_out1 <= Logical_Operator_out4117_out1 XOR Logical_Operator_out4373_out1;

  Logical_Operator_out4630_out1 <= Logical_Operator_out4118_out1 XOR Logical_Operator_out4374_out1;

  Logical_Operator_out4631_out1 <= Logical_Operator_out4119_out1 XOR Logical_Operator_out4375_out1;

  Logical_Operator_out4632_out1 <= Logical_Operator_out4120_out1 XOR Logical_Operator_out4376_out1;

  Logical_Operator_out4633_out1 <= Logical_Operator_out4121_out1 XOR Logical_Operator_out4377_out1;

  Logical_Operator_out4634_out1 <= Logical_Operator_out4122_out1 XOR Logical_Operator_out4378_out1;

  Logical_Operator_out4635_out1 <= Logical_Operator_out4123_out1 XOR Logical_Operator_out4379_out1;

  Logical_Operator_out4636_out1 <= Logical_Operator_out4124_out1 XOR Logical_Operator_out4380_out1;

  Logical_Operator_out4637_out1 <= Logical_Operator_out4125_out1 XOR Logical_Operator_out4381_out1;

  Logical_Operator_out4638_out1 <= Logical_Operator_out4126_out1 XOR Logical_Operator_out4382_out1;

  Logical_Operator_out4639_out1 <= Logical_Operator_out4127_out1 XOR Logical_Operator_out4383_out1;

  Logical_Operator_out4640_out1 <= Logical_Operator_out4128_out1 XOR Logical_Operator_out4384_out1;

  Logical_Operator_out4641_out1 <= Logical_Operator_out4129_out1 XOR Logical_Operator_out4385_out1;

  Logical_Operator_out4642_out1 <= Logical_Operator_out4130_out1 XOR Logical_Operator_out4386_out1;

  Logical_Operator_out4643_out1 <= Logical_Operator_out4131_out1 XOR Logical_Operator_out4387_out1;

  Logical_Operator_out4644_out1 <= Logical_Operator_out4132_out1 XOR Logical_Operator_out4388_out1;

  Logical_Operator_out4645_out1 <= Logical_Operator_out4133_out1 XOR Logical_Operator_out4389_out1;

  Logical_Operator_out4646_out1 <= Logical_Operator_out4134_out1 XOR Logical_Operator_out4390_out1;

  Logical_Operator_out4647_out1 <= Logical_Operator_out4135_out1 XOR Logical_Operator_out4391_out1;

  Logical_Operator_out4648_out1 <= Logical_Operator_out4136_out1 XOR Logical_Operator_out4392_out1;

  Logical_Operator_out4649_out1 <= Logical_Operator_out4137_out1 XOR Logical_Operator_out4393_out1;

  Logical_Operator_out4650_out1 <= Logical_Operator_out4138_out1 XOR Logical_Operator_out4394_out1;

  Logical_Operator_out4651_out1 <= Logical_Operator_out4139_out1 XOR Logical_Operator_out4395_out1;

  Logical_Operator_out4652_out1 <= Logical_Operator_out4140_out1 XOR Logical_Operator_out4396_out1;

  Logical_Operator_out4653_out1 <= Logical_Operator_out4141_out1 XOR Logical_Operator_out4397_out1;

  Logical_Operator_out4654_out1 <= Logical_Operator_out4142_out1 XOR Logical_Operator_out4398_out1;

  Logical_Operator_out4655_out1 <= Logical_Operator_out4143_out1 XOR Logical_Operator_out4399_out1;

  Logical_Operator_out4656_out1 <= Logical_Operator_out4144_out1 XOR Logical_Operator_out4400_out1;

  Logical_Operator_out4657_out1 <= Logical_Operator_out4145_out1 XOR Logical_Operator_out4401_out1;

  Logical_Operator_out4658_out1 <= Logical_Operator_out4146_out1 XOR Logical_Operator_out4402_out1;

  Logical_Operator_out4659_out1 <= Logical_Operator_out4147_out1 XOR Logical_Operator_out4403_out1;

  Logical_Operator_out4660_out1 <= Logical_Operator_out4148_out1 XOR Logical_Operator_out4404_out1;

  Logical_Operator_out4661_out1 <= Logical_Operator_out4149_out1 XOR Logical_Operator_out4405_out1;

  Logical_Operator_out4662_out1 <= Logical_Operator_out4150_out1 XOR Logical_Operator_out4406_out1;

  Logical_Operator_out4663_out1 <= Logical_Operator_out4151_out1 XOR Logical_Operator_out4407_out1;

  Logical_Operator_out4664_out1 <= Logical_Operator_out4152_out1 XOR Logical_Operator_out4408_out1;

  Logical_Operator_out4665_out1 <= Logical_Operator_out4153_out1 XOR Logical_Operator_out4409_out1;

  Logical_Operator_out4666_out1 <= Logical_Operator_out4154_out1 XOR Logical_Operator_out4410_out1;

  Logical_Operator_out4667_out1 <= Logical_Operator_out4155_out1 XOR Logical_Operator_out4411_out1;

  Logical_Operator_out4668_out1 <= Logical_Operator_out4156_out1 XOR Logical_Operator_out4412_out1;

  Logical_Operator_out4669_out1 <= Logical_Operator_out4157_out1 XOR Logical_Operator_out4413_out1;

  Logical_Operator_out4670_out1 <= Logical_Operator_out4158_out1 XOR Logical_Operator_out4414_out1;

  Logical_Operator_out4671_out1 <= Logical_Operator_out4159_out1 XOR Logical_Operator_out4415_out1;

  Logical_Operator_out4672_out1 <= Logical_Operator_out4160_out1 XOR Logical_Operator_out4416_out1;

  Logical_Operator_out4673_out1 <= Logical_Operator_out4161_out1 XOR Logical_Operator_out4417_out1;

  Logical_Operator_out4674_out1 <= Logical_Operator_out4162_out1 XOR Logical_Operator_out4418_out1;

  Logical_Operator_out4675_out1 <= Logical_Operator_out4163_out1 XOR Logical_Operator_out4419_out1;

  Logical_Operator_out4676_out1 <= Logical_Operator_out4164_out1 XOR Logical_Operator_out4420_out1;

  Logical_Operator_out4677_out1 <= Logical_Operator_out4165_out1 XOR Logical_Operator_out4421_out1;

  Logical_Operator_out4678_out1 <= Logical_Operator_out4166_out1 XOR Logical_Operator_out4422_out1;

  Logical_Operator_out4679_out1 <= Logical_Operator_out4167_out1 XOR Logical_Operator_out4423_out1;

  Logical_Operator_out4680_out1 <= Logical_Operator_out4168_out1 XOR Logical_Operator_out4424_out1;

  Logical_Operator_out4681_out1 <= Logical_Operator_out4169_out1 XOR Logical_Operator_out4425_out1;

  Logical_Operator_out4682_out1 <= Logical_Operator_out4170_out1 XOR Logical_Operator_out4426_out1;

  Logical_Operator_out4683_out1 <= Logical_Operator_out4171_out1 XOR Logical_Operator_out4427_out1;

  Logical_Operator_out4684_out1 <= Logical_Operator_out4172_out1 XOR Logical_Operator_out4428_out1;

  Logical_Operator_out4685_out1 <= Logical_Operator_out4173_out1 XOR Logical_Operator_out4429_out1;

  Logical_Operator_out4686_out1 <= Logical_Operator_out4174_out1 XOR Logical_Operator_out4430_out1;

  Logical_Operator_out4687_out1 <= Logical_Operator_out4175_out1 XOR Logical_Operator_out4431_out1;

  Logical_Operator_out4688_out1 <= Logical_Operator_out4176_out1 XOR Logical_Operator_out4432_out1;

  Logical_Operator_out4689_out1 <= Logical_Operator_out4177_out1 XOR Logical_Operator_out4433_out1;

  Logical_Operator_out4690_out1 <= Logical_Operator_out4178_out1 XOR Logical_Operator_out4434_out1;

  Logical_Operator_out4691_out1 <= Logical_Operator_out4179_out1 XOR Logical_Operator_out4435_out1;

  Logical_Operator_out4692_out1 <= Logical_Operator_out4180_out1 XOR Logical_Operator_out4436_out1;

  Logical_Operator_out4693_out1 <= Logical_Operator_out4181_out1 XOR Logical_Operator_out4437_out1;

  Logical_Operator_out4694_out1 <= Logical_Operator_out4182_out1 XOR Logical_Operator_out4438_out1;

  Logical_Operator_out4695_out1 <= Logical_Operator_out4183_out1 XOR Logical_Operator_out4439_out1;

  Logical_Operator_out4696_out1 <= Logical_Operator_out4184_out1 XOR Logical_Operator_out4440_out1;

  Logical_Operator_out4697_out1 <= Logical_Operator_out4185_out1 XOR Logical_Operator_out4441_out1;

  Logical_Operator_out4698_out1 <= Logical_Operator_out4186_out1 XOR Logical_Operator_out4442_out1;

  Logical_Operator_out4699_out1 <= Logical_Operator_out4187_out1 XOR Logical_Operator_out4443_out1;

  Logical_Operator_out4700_out1 <= Logical_Operator_out4188_out1 XOR Logical_Operator_out4444_out1;

  Logical_Operator_out4701_out1 <= Logical_Operator_out4189_out1 XOR Logical_Operator_out4445_out1;

  Logical_Operator_out4702_out1 <= Logical_Operator_out4190_out1 XOR Logical_Operator_out4446_out1;

  Logical_Operator_out4703_out1 <= Logical_Operator_out4191_out1 XOR Logical_Operator_out4447_out1;

  Logical_Operator_out4704_out1 <= Logical_Operator_out4192_out1 XOR Logical_Operator_out4448_out1;

  Logical_Operator_out4705_out1 <= Logical_Operator_out4193_out1 XOR Logical_Operator_out4449_out1;

  Logical_Operator_out4706_out1 <= Logical_Operator_out4194_out1 XOR Logical_Operator_out4450_out1;

  Logical_Operator_out4707_out1 <= Logical_Operator_out4195_out1 XOR Logical_Operator_out4451_out1;

  Logical_Operator_out4708_out1 <= Logical_Operator_out4196_out1 XOR Logical_Operator_out4452_out1;

  Logical_Operator_out4709_out1 <= Logical_Operator_out4197_out1 XOR Logical_Operator_out4453_out1;

  Logical_Operator_out4710_out1 <= Logical_Operator_out4198_out1 XOR Logical_Operator_out4454_out1;

  Logical_Operator_out4711_out1 <= Logical_Operator_out4199_out1 XOR Logical_Operator_out4455_out1;

  Logical_Operator_out4712_out1 <= Logical_Operator_out4200_out1 XOR Logical_Operator_out4456_out1;

  Logical_Operator_out4713_out1 <= Logical_Operator_out4201_out1 XOR Logical_Operator_out4457_out1;

  Logical_Operator_out4714_out1 <= Logical_Operator_out4202_out1 XOR Logical_Operator_out4458_out1;

  Logical_Operator_out4715_out1 <= Logical_Operator_out4203_out1 XOR Logical_Operator_out4459_out1;

  Logical_Operator_out4716_out1 <= Logical_Operator_out4204_out1 XOR Logical_Operator_out4460_out1;

  Logical_Operator_out4717_out1 <= Logical_Operator_out4205_out1 XOR Logical_Operator_out4461_out1;

  Logical_Operator_out4718_out1 <= Logical_Operator_out4206_out1 XOR Logical_Operator_out4462_out1;

  Logical_Operator_out4719_out1 <= Logical_Operator_out4207_out1 XOR Logical_Operator_out4463_out1;

  Logical_Operator_out4720_out1 <= Logical_Operator_out4208_out1 XOR Logical_Operator_out4464_out1;

  Logical_Operator_out4721_out1 <= Logical_Operator_out4209_out1 XOR Logical_Operator_out4465_out1;

  Logical_Operator_out4722_out1 <= Logical_Operator_out4210_out1 XOR Logical_Operator_out4466_out1;

  Logical_Operator_out4723_out1 <= Logical_Operator_out4211_out1 XOR Logical_Operator_out4467_out1;

  Logical_Operator_out4724_out1 <= Logical_Operator_out4212_out1 XOR Logical_Operator_out4468_out1;

  Logical_Operator_out4725_out1 <= Logical_Operator_out4213_out1 XOR Logical_Operator_out4469_out1;

  Logical_Operator_out4726_out1 <= Logical_Operator_out4214_out1 XOR Logical_Operator_out4470_out1;

  Logical_Operator_out4727_out1 <= Logical_Operator_out4215_out1 XOR Logical_Operator_out4471_out1;

  Logical_Operator_out4728_out1 <= Logical_Operator_out4216_out1 XOR Logical_Operator_out4472_out1;

  Logical_Operator_out4729_out1 <= Logical_Operator_out4217_out1 XOR Logical_Operator_out4473_out1;

  Logical_Operator_out4730_out1 <= Logical_Operator_out4218_out1 XOR Logical_Operator_out4474_out1;

  Logical_Operator_out4731_out1 <= Logical_Operator_out4219_out1 XOR Logical_Operator_out4475_out1;

  Logical_Operator_out4732_out1 <= Logical_Operator_out4220_out1 XOR Logical_Operator_out4476_out1;

  Logical_Operator_out4733_out1 <= Logical_Operator_out4221_out1 XOR Logical_Operator_out4477_out1;

  Logical_Operator_out4734_out1 <= Logical_Operator_out4222_out1 XOR Logical_Operator_out4478_out1;

  Logical_Operator_out4735_out1 <= Logical_Operator_out4223_out1 XOR Logical_Operator_out4479_out1;

  Logical_Operator_out4736_out1 <= Logical_Operator_out4224_out1 XOR Logical_Operator_out4480_out1;

  Logical_Operator_out4737_out1 <= Logical_Operator_out4225_out1 XOR Logical_Operator_out4481_out1;

  Logical_Operator_out4738_out1 <= Logical_Operator_out4226_out1 XOR Logical_Operator_out4482_out1;

  Logical_Operator_out4739_out1 <= Logical_Operator_out4227_out1 XOR Logical_Operator_out4483_out1;

  Logical_Operator_out4740_out1 <= Logical_Operator_out4228_out1 XOR Logical_Operator_out4484_out1;

  Logical_Operator_out4741_out1 <= Logical_Operator_out4229_out1 XOR Logical_Operator_out4485_out1;

  Logical_Operator_out4742_out1 <= Logical_Operator_out4230_out1 XOR Logical_Operator_out4486_out1;

  Logical_Operator_out4743_out1 <= Logical_Operator_out4231_out1 XOR Logical_Operator_out4487_out1;

  Logical_Operator_out4744_out1 <= Logical_Operator_out4232_out1 XOR Logical_Operator_out4488_out1;

  Logical_Operator_out4745_out1 <= Logical_Operator_out4233_out1 XOR Logical_Operator_out4489_out1;

  Logical_Operator_out4746_out1 <= Logical_Operator_out4234_out1 XOR Logical_Operator_out4490_out1;

  Logical_Operator_out4747_out1 <= Logical_Operator_out4235_out1 XOR Logical_Operator_out4491_out1;

  Logical_Operator_out4748_out1 <= Logical_Operator_out4236_out1 XOR Logical_Operator_out4492_out1;

  Logical_Operator_out4749_out1 <= Logical_Operator_out4237_out1 XOR Logical_Operator_out4493_out1;

  Logical_Operator_out4750_out1 <= Logical_Operator_out4238_out1 XOR Logical_Operator_out4494_out1;

  Logical_Operator_out4751_out1 <= Logical_Operator_out4239_out1 XOR Logical_Operator_out4495_out1;

  Logical_Operator_out4752_out1 <= Logical_Operator_out4240_out1 XOR Logical_Operator_out4496_out1;

  Logical_Operator_out4753_out1 <= Logical_Operator_out4241_out1 XOR Logical_Operator_out4497_out1;

  Logical_Operator_out4754_out1 <= Logical_Operator_out4242_out1 XOR Logical_Operator_out4498_out1;

  Logical_Operator_out4755_out1 <= Logical_Operator_out4243_out1 XOR Logical_Operator_out4499_out1;

  Logical_Operator_out4756_out1 <= Logical_Operator_out4244_out1 XOR Logical_Operator_out4500_out1;

  Logical_Operator_out4757_out1 <= Logical_Operator_out4245_out1 XOR Logical_Operator_out4501_out1;

  Logical_Operator_out4758_out1 <= Logical_Operator_out4246_out1 XOR Logical_Operator_out4502_out1;

  Logical_Operator_out4759_out1 <= Logical_Operator_out4247_out1 XOR Logical_Operator_out4503_out1;

  Logical_Operator_out4760_out1 <= Logical_Operator_out4248_out1 XOR Logical_Operator_out4504_out1;

  Logical_Operator_out4761_out1 <= Logical_Operator_out4249_out1 XOR Logical_Operator_out4505_out1;

  Logical_Operator_out4762_out1 <= Logical_Operator_out4250_out1 XOR Logical_Operator_out4506_out1;

  Logical_Operator_out4763_out1 <= Logical_Operator_out4251_out1 XOR Logical_Operator_out4507_out1;

  Logical_Operator_out4764_out1 <= Logical_Operator_out4252_out1 XOR Logical_Operator_out4508_out1;

  Logical_Operator_out4765_out1 <= Logical_Operator_out4253_out1 XOR Logical_Operator_out4509_out1;

  Logical_Operator_out4766_out1 <= Logical_Operator_out4254_out1 XOR Logical_Operator_out4510_out1;

  Logical_Operator_out4767_out1 <= Logical_Operator_out4255_out1 XOR Logical_Operator_out4511_out1;

  Logical_Operator_out4768_out1 <= Logical_Operator_out4256_out1 XOR Logical_Operator_out4512_out1;

  Logical_Operator_out4769_out1 <= Logical_Operator_out4257_out1 XOR Logical_Operator_out4513_out1;

  Logical_Operator_out4770_out1 <= Logical_Operator_out4258_out1 XOR Logical_Operator_out4514_out1;

  Logical_Operator_out4771_out1 <= Logical_Operator_out4259_out1 XOR Logical_Operator_out4515_out1;

  Logical_Operator_out4772_out1 <= Logical_Operator_out4260_out1 XOR Logical_Operator_out4516_out1;

  Logical_Operator_out4773_out1 <= Logical_Operator_out4261_out1 XOR Logical_Operator_out4517_out1;

  Logical_Operator_out4774_out1 <= Logical_Operator_out4262_out1 XOR Logical_Operator_out4518_out1;

  Logical_Operator_out4775_out1 <= Logical_Operator_out4263_out1 XOR Logical_Operator_out4519_out1;

  Logical_Operator_out4776_out1 <= Logical_Operator_out4264_out1 XOR Logical_Operator_out4520_out1;

  Logical_Operator_out4777_out1 <= Logical_Operator_out4265_out1 XOR Logical_Operator_out4521_out1;

  Logical_Operator_out4778_out1 <= Logical_Operator_out4266_out1 XOR Logical_Operator_out4522_out1;

  Logical_Operator_out4779_out1 <= Logical_Operator_out4267_out1 XOR Logical_Operator_out4523_out1;

  Logical_Operator_out4780_out1 <= Logical_Operator_out4268_out1 XOR Logical_Operator_out4524_out1;

  Logical_Operator_out4781_out1 <= Logical_Operator_out4269_out1 XOR Logical_Operator_out4525_out1;

  Logical_Operator_out4782_out1 <= Logical_Operator_out4270_out1 XOR Logical_Operator_out4526_out1;

  Logical_Operator_out4783_out1 <= Logical_Operator_out4271_out1 XOR Logical_Operator_out4527_out1;

  Logical_Operator_out4784_out1 <= Logical_Operator_out4272_out1 XOR Logical_Operator_out4528_out1;

  Logical_Operator_out4785_out1 <= Logical_Operator_out4273_out1 XOR Logical_Operator_out4529_out1;

  Logical_Operator_out4786_out1 <= Logical_Operator_out4274_out1 XOR Logical_Operator_out4530_out1;

  Logical_Operator_out4787_out1 <= Logical_Operator_out4275_out1 XOR Logical_Operator_out4531_out1;

  Logical_Operator_out4788_out1 <= Logical_Operator_out4276_out1 XOR Logical_Operator_out4532_out1;

  Logical_Operator_out4789_out1 <= Logical_Operator_out4277_out1 XOR Logical_Operator_out4533_out1;

  Logical_Operator_out4790_out1 <= Logical_Operator_out4278_out1 XOR Logical_Operator_out4534_out1;

  Logical_Operator_out4791_out1 <= Logical_Operator_out4279_out1 XOR Logical_Operator_out4535_out1;

  Logical_Operator_out4792_out1 <= Logical_Operator_out4280_out1 XOR Logical_Operator_out4536_out1;

  Logical_Operator_out4793_out1 <= Logical_Operator_out4281_out1 XOR Logical_Operator_out4537_out1;

  Logical_Operator_out4794_out1 <= Logical_Operator_out4282_out1 XOR Logical_Operator_out4538_out1;

  Logical_Operator_out4795_out1 <= Logical_Operator_out4283_out1 XOR Logical_Operator_out4539_out1;

  Logical_Operator_out4796_out1 <= Logical_Operator_out4284_out1 XOR Logical_Operator_out4540_out1;

  Logical_Operator_out4797_out1 <= Logical_Operator_out4285_out1 XOR Logical_Operator_out4541_out1;

  Logical_Operator_out4798_out1 <= Logical_Operator_out4286_out1 XOR Logical_Operator_out4542_out1;

  Logical_Operator_out4799_out1 <= Logical_Operator_out4287_out1 XOR Logical_Operator_out4543_out1;

  Logical_Operator_out4800_out1 <= Logical_Operator_out4288_out1 XOR Logical_Operator_out4544_out1;

  Logical_Operator_out4801_out1 <= Logical_Operator_out4289_out1 XOR Logical_Operator_out4545_out1;

  Logical_Operator_out4802_out1 <= Logical_Operator_out4290_out1 XOR Logical_Operator_out4546_out1;

  Logical_Operator_out4803_out1 <= Logical_Operator_out4291_out1 XOR Logical_Operator_out4547_out1;

  Logical_Operator_out4804_out1 <= Logical_Operator_out4292_out1 XOR Logical_Operator_out4548_out1;

  Logical_Operator_out4805_out1 <= Logical_Operator_out4293_out1 XOR Logical_Operator_out4549_out1;

  Logical_Operator_out4806_out1 <= Logical_Operator_out4294_out1 XOR Logical_Operator_out4550_out1;

  Logical_Operator_out4807_out1 <= Logical_Operator_out4295_out1 XOR Logical_Operator_out4551_out1;

  Logical_Operator_out4808_out1 <= Logical_Operator_out4296_out1 XOR Logical_Operator_out4552_out1;

  Logical_Operator_out4809_out1 <= Logical_Operator_out4297_out1 XOR Logical_Operator_out4553_out1;

  Logical_Operator_out4810_out1 <= Logical_Operator_out4298_out1 XOR Logical_Operator_out4554_out1;

  Logical_Operator_out4811_out1 <= Logical_Operator_out4299_out1 XOR Logical_Operator_out4555_out1;

  Logical_Operator_out4812_out1 <= Logical_Operator_out4300_out1 XOR Logical_Operator_out4556_out1;

  Logical_Operator_out4813_out1 <= Logical_Operator_out4301_out1 XOR Logical_Operator_out4557_out1;

  Logical_Operator_out4814_out1 <= Logical_Operator_out4302_out1 XOR Logical_Operator_out4558_out1;

  Logical_Operator_out4815_out1 <= Logical_Operator_out4303_out1 XOR Logical_Operator_out4559_out1;

  Logical_Operator_out4816_out1 <= Logical_Operator_out4304_out1 XOR Logical_Operator_out4560_out1;

  Logical_Operator_out4817_out1 <= Logical_Operator_out4305_out1 XOR Logical_Operator_out4561_out1;

  Logical_Operator_out4818_out1 <= Logical_Operator_out4306_out1 XOR Logical_Operator_out4562_out1;

  Logical_Operator_out4819_out1 <= Logical_Operator_out4307_out1 XOR Logical_Operator_out4563_out1;

  Logical_Operator_out4820_out1 <= Logical_Operator_out4308_out1 XOR Logical_Operator_out4564_out1;

  Logical_Operator_out4821_out1 <= Logical_Operator_out4309_out1 XOR Logical_Operator_out4565_out1;

  Logical_Operator_out4822_out1 <= Logical_Operator_out4310_out1 XOR Logical_Operator_out4566_out1;

  Logical_Operator_out4823_out1 <= Logical_Operator_out4311_out1 XOR Logical_Operator_out4567_out1;

  Logical_Operator_out4824_out1 <= Logical_Operator_out4312_out1 XOR Logical_Operator_out4568_out1;

  Logical_Operator_out4825_out1 <= Logical_Operator_out4313_out1 XOR Logical_Operator_out4569_out1;

  Logical_Operator_out4826_out1 <= Logical_Operator_out4314_out1 XOR Logical_Operator_out4570_out1;

  Logical_Operator_out4827_out1 <= Logical_Operator_out4315_out1 XOR Logical_Operator_out4571_out1;

  Logical_Operator_out4828_out1 <= Logical_Operator_out4316_out1 XOR Logical_Operator_out4572_out1;

  Logical_Operator_out4829_out1 <= Logical_Operator_out4317_out1 XOR Logical_Operator_out4573_out1;

  Logical_Operator_out4830_out1 <= Logical_Operator_out4318_out1 XOR Logical_Operator_out4574_out1;

  Logical_Operator_out4831_out1 <= Logical_Operator_out4319_out1 XOR Logical_Operator_out4575_out1;

  Logical_Operator_out4832_out1 <= Logical_Operator_out4320_out1 XOR Logical_Operator_out4576_out1;

  Logical_Operator_out4833_out1 <= Logical_Operator_out4321_out1 XOR Logical_Operator_out4577_out1;

  Logical_Operator_out4834_out1 <= Logical_Operator_out4322_out1 XOR Logical_Operator_out4578_out1;

  Logical_Operator_out4835_out1 <= Logical_Operator_out4323_out1 XOR Logical_Operator_out4579_out1;

  Logical_Operator_out4836_out1 <= Logical_Operator_out4324_out1 XOR Logical_Operator_out4580_out1;

  Logical_Operator_out4837_out1 <= Logical_Operator_out4325_out1 XOR Logical_Operator_out4581_out1;

  Logical_Operator_out4838_out1 <= Logical_Operator_out4326_out1 XOR Logical_Operator_out4582_out1;

  Logical_Operator_out4839_out1 <= Logical_Operator_out4327_out1 XOR Logical_Operator_out4583_out1;

  Logical_Operator_out4840_out1 <= Logical_Operator_out4328_out1 XOR Logical_Operator_out4584_out1;

  Logical_Operator_out4841_out1 <= Logical_Operator_out4329_out1 XOR Logical_Operator_out4585_out1;

  Logical_Operator_out4842_out1 <= Logical_Operator_out4330_out1 XOR Logical_Operator_out4586_out1;

  Logical_Operator_out4843_out1 <= Logical_Operator_out4331_out1 XOR Logical_Operator_out4587_out1;

  Logical_Operator_out4844_out1 <= Logical_Operator_out4332_out1 XOR Logical_Operator_out4588_out1;

  Logical_Operator_out4845_out1 <= Logical_Operator_out4333_out1 XOR Logical_Operator_out4589_out1;

  Logical_Operator_out4846_out1 <= Logical_Operator_out4334_out1 XOR Logical_Operator_out4590_out1;

  Logical_Operator_out4847_out1 <= Logical_Operator_out4335_out1 XOR Logical_Operator_out4591_out1;

  Logical_Operator_out4848_out1 <= Logical_Operator_out4336_out1 XOR Logical_Operator_out4592_out1;

  Logical_Operator_out4849_out1 <= Logical_Operator_out4337_out1 XOR Logical_Operator_out4593_out1;

  Logical_Operator_out4850_out1 <= Logical_Operator_out4338_out1 XOR Logical_Operator_out4594_out1;

  Logical_Operator_out4851_out1 <= Logical_Operator_out4339_out1 XOR Logical_Operator_out4595_out1;

  Logical_Operator_out4852_out1 <= Logical_Operator_out4340_out1 XOR Logical_Operator_out4596_out1;

  Logical_Operator_out4853_out1 <= Logical_Operator_out4341_out1 XOR Logical_Operator_out4597_out1;

  Logical_Operator_out4854_out1 <= Logical_Operator_out4342_out1 XOR Logical_Operator_out4598_out1;

  Logical_Operator_out4855_out1 <= Logical_Operator_out4343_out1 XOR Logical_Operator_out4599_out1;

  Logical_Operator_out4856_out1 <= Logical_Operator_out4344_out1 XOR Logical_Operator_out4600_out1;

  Logical_Operator_out4857_out1 <= Logical_Operator_out4345_out1 XOR Logical_Operator_out4601_out1;

  Logical_Operator_out4858_out1 <= Logical_Operator_out4346_out1 XOR Logical_Operator_out4602_out1;

  Logical_Operator_out4859_out1 <= Logical_Operator_out4347_out1 XOR Logical_Operator_out4603_out1;

  Logical_Operator_out4860_out1 <= Logical_Operator_out4348_out1 XOR Logical_Operator_out4604_out1;

  Logical_Operator_out4861_out1 <= Logical_Operator_out4349_out1 XOR Logical_Operator_out4605_out1;

  Logical_Operator_out4862_out1 <= Logical_Operator_out4350_out1 XOR Logical_Operator_out4606_out1;

  Logical_Operator_out4863_out1 <= Logical_Operator_out4351_out1 XOR Logical_Operator_out4607_out1;

  Logical_Operator_out4864_out1 <= Logical_Operator_out4352_out1 XOR Logical_Operator_out4608_out1;

  Logical_Operator_out4865_out1 <= Logical_Operator_out3713_out1 XOR Logical_Operator_out3969_out1;

  Logical_Operator_out4866_out1 <= Logical_Operator_out3714_out1 XOR Logical_Operator_out3970_out1;

  Logical_Operator_out4867_out1 <= Logical_Operator_out3715_out1 XOR Logical_Operator_out3971_out1;

  Logical_Operator_out4868_out1 <= Logical_Operator_out3716_out1 XOR Logical_Operator_out3972_out1;

  Logical_Operator_out4869_out1 <= Logical_Operator_out3717_out1 XOR Logical_Operator_out3973_out1;

  Logical_Operator_out4870_out1 <= Logical_Operator_out3718_out1 XOR Logical_Operator_out3974_out1;

  Logical_Operator_out4871_out1 <= Logical_Operator_out3719_out1 XOR Logical_Operator_out3975_out1;

  Logical_Operator_out4872_out1 <= Logical_Operator_out3720_out1 XOR Logical_Operator_out3976_out1;

  Logical_Operator_out4873_out1 <= Logical_Operator_out3721_out1 XOR Logical_Operator_out3977_out1;

  Logical_Operator_out4874_out1 <= Logical_Operator_out3722_out1 XOR Logical_Operator_out3978_out1;

  Logical_Operator_out4875_out1 <= Logical_Operator_out3723_out1 XOR Logical_Operator_out3979_out1;

  Logical_Operator_out4876_out1 <= Logical_Operator_out3724_out1 XOR Logical_Operator_out3980_out1;

  Logical_Operator_out4877_out1 <= Logical_Operator_out3725_out1 XOR Logical_Operator_out3981_out1;

  Logical_Operator_out4878_out1 <= Logical_Operator_out3726_out1 XOR Logical_Operator_out3982_out1;

  Logical_Operator_out4879_out1 <= Logical_Operator_out3727_out1 XOR Logical_Operator_out3983_out1;

  Logical_Operator_out4880_out1 <= Logical_Operator_out3728_out1 XOR Logical_Operator_out3984_out1;

  Logical_Operator_out4881_out1 <= Logical_Operator_out3729_out1 XOR Logical_Operator_out3985_out1;

  Logical_Operator_out4882_out1 <= Logical_Operator_out3730_out1 XOR Logical_Operator_out3986_out1;

  Logical_Operator_out4883_out1 <= Logical_Operator_out3731_out1 XOR Logical_Operator_out3987_out1;

  Logical_Operator_out4884_out1 <= Logical_Operator_out3732_out1 XOR Logical_Operator_out3988_out1;

  Logical_Operator_out4885_out1 <= Logical_Operator_out3733_out1 XOR Logical_Operator_out3989_out1;

  Logical_Operator_out4886_out1 <= Logical_Operator_out3734_out1 XOR Logical_Operator_out3990_out1;

  Logical_Operator_out4887_out1 <= Logical_Operator_out3735_out1 XOR Logical_Operator_out3991_out1;

  Logical_Operator_out4888_out1 <= Logical_Operator_out3736_out1 XOR Logical_Operator_out3992_out1;

  Logical_Operator_out4889_out1 <= Logical_Operator_out3737_out1 XOR Logical_Operator_out3993_out1;

  Logical_Operator_out4890_out1 <= Logical_Operator_out3738_out1 XOR Logical_Operator_out3994_out1;

  Logical_Operator_out4891_out1 <= Logical_Operator_out3739_out1 XOR Logical_Operator_out3995_out1;

  Logical_Operator_out4892_out1 <= Logical_Operator_out3740_out1 XOR Logical_Operator_out3996_out1;

  Logical_Operator_out4893_out1 <= Logical_Operator_out3741_out1 XOR Logical_Operator_out3997_out1;

  Logical_Operator_out4894_out1 <= Logical_Operator_out3742_out1 XOR Logical_Operator_out3998_out1;

  Logical_Operator_out4895_out1 <= Logical_Operator_out3743_out1 XOR Logical_Operator_out3999_out1;

  Logical_Operator_out4896_out1 <= Logical_Operator_out3744_out1 XOR Logical_Operator_out4000_out1;

  Logical_Operator_out4897_out1 <= Logical_Operator_out3745_out1 XOR Logical_Operator_out4001_out1;

  Logical_Operator_out4898_out1 <= Logical_Operator_out3746_out1 XOR Logical_Operator_out4002_out1;

  Logical_Operator_out4899_out1 <= Logical_Operator_out3747_out1 XOR Logical_Operator_out4003_out1;

  Logical_Operator_out4900_out1 <= Logical_Operator_out3748_out1 XOR Logical_Operator_out4004_out1;

  Logical_Operator_out4901_out1 <= Logical_Operator_out3749_out1 XOR Logical_Operator_out4005_out1;

  Logical_Operator_out4902_out1 <= Logical_Operator_out3750_out1 XOR Logical_Operator_out4006_out1;

  Logical_Operator_out4903_out1 <= Logical_Operator_out3751_out1 XOR Logical_Operator_out4007_out1;

  Logical_Operator_out4904_out1 <= Logical_Operator_out3752_out1 XOR Logical_Operator_out4008_out1;

  Logical_Operator_out4905_out1 <= Logical_Operator_out3753_out1 XOR Logical_Operator_out4009_out1;

  Logical_Operator_out4906_out1 <= Logical_Operator_out3754_out1 XOR Logical_Operator_out4010_out1;

  Logical_Operator_out4907_out1 <= Logical_Operator_out3755_out1 XOR Logical_Operator_out4011_out1;

  Logical_Operator_out4908_out1 <= Logical_Operator_out3756_out1 XOR Logical_Operator_out4012_out1;

  Logical_Operator_out4909_out1 <= Logical_Operator_out3757_out1 XOR Logical_Operator_out4013_out1;

  Logical_Operator_out4910_out1 <= Logical_Operator_out3758_out1 XOR Logical_Operator_out4014_out1;

  Logical_Operator_out4911_out1 <= Logical_Operator_out3759_out1 XOR Logical_Operator_out4015_out1;

  Logical_Operator_out4912_out1 <= Logical_Operator_out3760_out1 XOR Logical_Operator_out4016_out1;

  Logical_Operator_out4913_out1 <= Logical_Operator_out3761_out1 XOR Logical_Operator_out4017_out1;

  Logical_Operator_out4914_out1 <= Logical_Operator_out3762_out1 XOR Logical_Operator_out4018_out1;

  Logical_Operator_out4915_out1 <= Logical_Operator_out3763_out1 XOR Logical_Operator_out4019_out1;

  Logical_Operator_out4916_out1 <= Logical_Operator_out3764_out1 XOR Logical_Operator_out4020_out1;

  Logical_Operator_out4917_out1 <= Logical_Operator_out3765_out1 XOR Logical_Operator_out4021_out1;

  Logical_Operator_out4918_out1 <= Logical_Operator_out3766_out1 XOR Logical_Operator_out4022_out1;

  Logical_Operator_out4919_out1 <= Logical_Operator_out3767_out1 XOR Logical_Operator_out4023_out1;

  Logical_Operator_out4920_out1 <= Logical_Operator_out3768_out1 XOR Logical_Operator_out4024_out1;

  Logical_Operator_out4921_out1 <= Logical_Operator_out3769_out1 XOR Logical_Operator_out4025_out1;

  Logical_Operator_out4922_out1 <= Logical_Operator_out3770_out1 XOR Logical_Operator_out4026_out1;

  Logical_Operator_out4923_out1 <= Logical_Operator_out3771_out1 XOR Logical_Operator_out4027_out1;

  Logical_Operator_out4924_out1 <= Logical_Operator_out3772_out1 XOR Logical_Operator_out4028_out1;

  Logical_Operator_out4925_out1 <= Logical_Operator_out3773_out1 XOR Logical_Operator_out4029_out1;

  Logical_Operator_out4926_out1 <= Logical_Operator_out3774_out1 XOR Logical_Operator_out4030_out1;

  Logical_Operator_out4927_out1 <= Logical_Operator_out3775_out1 XOR Logical_Operator_out4031_out1;

  Logical_Operator_out4928_out1 <= Logical_Operator_out3776_out1 XOR Logical_Operator_out4032_out1;

  Logical_Operator_out4929_out1 <= Logical_Operator_out3777_out1 XOR Logical_Operator_out4033_out1;

  Logical_Operator_out4930_out1 <= Logical_Operator_out3778_out1 XOR Logical_Operator_out4034_out1;

  Logical_Operator_out4931_out1 <= Logical_Operator_out3779_out1 XOR Logical_Operator_out4035_out1;

  Logical_Operator_out4932_out1 <= Logical_Operator_out3780_out1 XOR Logical_Operator_out4036_out1;

  Logical_Operator_out4933_out1 <= Logical_Operator_out3781_out1 XOR Logical_Operator_out4037_out1;

  Logical_Operator_out4934_out1 <= Logical_Operator_out3782_out1 XOR Logical_Operator_out4038_out1;

  Logical_Operator_out4935_out1 <= Logical_Operator_out3783_out1 XOR Logical_Operator_out4039_out1;

  Logical_Operator_out4936_out1 <= Logical_Operator_out3784_out1 XOR Logical_Operator_out4040_out1;

  Logical_Operator_out4937_out1 <= Logical_Operator_out3785_out1 XOR Logical_Operator_out4041_out1;

  Logical_Operator_out4938_out1 <= Logical_Operator_out3786_out1 XOR Logical_Operator_out4042_out1;

  Logical_Operator_out4939_out1 <= Logical_Operator_out3787_out1 XOR Logical_Operator_out4043_out1;

  Logical_Operator_out4940_out1 <= Logical_Operator_out3788_out1 XOR Logical_Operator_out4044_out1;

  Logical_Operator_out4941_out1 <= Logical_Operator_out3789_out1 XOR Logical_Operator_out4045_out1;

  Logical_Operator_out4942_out1 <= Logical_Operator_out3790_out1 XOR Logical_Operator_out4046_out1;

  Logical_Operator_out4943_out1 <= Logical_Operator_out3791_out1 XOR Logical_Operator_out4047_out1;

  Logical_Operator_out4944_out1 <= Logical_Operator_out3792_out1 XOR Logical_Operator_out4048_out1;

  Logical_Operator_out4945_out1 <= Logical_Operator_out3793_out1 XOR Logical_Operator_out4049_out1;

  Logical_Operator_out4946_out1 <= Logical_Operator_out3794_out1 XOR Logical_Operator_out4050_out1;

  Logical_Operator_out4947_out1 <= Logical_Operator_out3795_out1 XOR Logical_Operator_out4051_out1;

  Logical_Operator_out4948_out1 <= Logical_Operator_out3796_out1 XOR Logical_Operator_out4052_out1;

  Logical_Operator_out4949_out1 <= Logical_Operator_out3797_out1 XOR Logical_Operator_out4053_out1;

  Logical_Operator_out4950_out1 <= Logical_Operator_out3798_out1 XOR Logical_Operator_out4054_out1;

  Logical_Operator_out4951_out1 <= Logical_Operator_out3799_out1 XOR Logical_Operator_out4055_out1;

  Logical_Operator_out4952_out1 <= Logical_Operator_out3800_out1 XOR Logical_Operator_out4056_out1;

  Logical_Operator_out4953_out1 <= Logical_Operator_out3801_out1 XOR Logical_Operator_out4057_out1;

  Logical_Operator_out4954_out1 <= Logical_Operator_out3802_out1 XOR Logical_Operator_out4058_out1;

  Logical_Operator_out4955_out1 <= Logical_Operator_out3803_out1 XOR Logical_Operator_out4059_out1;

  Logical_Operator_out4956_out1 <= Logical_Operator_out3804_out1 XOR Logical_Operator_out4060_out1;

  Logical_Operator_out4957_out1 <= Logical_Operator_out3805_out1 XOR Logical_Operator_out4061_out1;

  Logical_Operator_out4958_out1 <= Logical_Operator_out3806_out1 XOR Logical_Operator_out4062_out1;

  Logical_Operator_out4959_out1 <= Logical_Operator_out3807_out1 XOR Logical_Operator_out4063_out1;

  Logical_Operator_out4960_out1 <= Logical_Operator_out3808_out1 XOR Logical_Operator_out4064_out1;

  Logical_Operator_out4961_out1 <= Logical_Operator_out3809_out1 XOR Logical_Operator_out4065_out1;

  Logical_Operator_out4962_out1 <= Logical_Operator_out3810_out1 XOR Logical_Operator_out4066_out1;

  Logical_Operator_out4963_out1 <= Logical_Operator_out3811_out1 XOR Logical_Operator_out4067_out1;

  Logical_Operator_out4964_out1 <= Logical_Operator_out3812_out1 XOR Logical_Operator_out4068_out1;

  Logical_Operator_out4965_out1 <= Logical_Operator_out3813_out1 XOR Logical_Operator_out4069_out1;

  Logical_Operator_out4966_out1 <= Logical_Operator_out3814_out1 XOR Logical_Operator_out4070_out1;

  Logical_Operator_out4967_out1 <= Logical_Operator_out3815_out1 XOR Logical_Operator_out4071_out1;

  Logical_Operator_out4968_out1 <= Logical_Operator_out3816_out1 XOR Logical_Operator_out4072_out1;

  Logical_Operator_out4969_out1 <= Logical_Operator_out3817_out1 XOR Logical_Operator_out4073_out1;

  Logical_Operator_out4970_out1 <= Logical_Operator_out3818_out1 XOR Logical_Operator_out4074_out1;

  Logical_Operator_out4971_out1 <= Logical_Operator_out3819_out1 XOR Logical_Operator_out4075_out1;

  Logical_Operator_out4972_out1 <= Logical_Operator_out3820_out1 XOR Logical_Operator_out4076_out1;

  Logical_Operator_out4973_out1 <= Logical_Operator_out3821_out1 XOR Logical_Operator_out4077_out1;

  Logical_Operator_out4974_out1 <= Logical_Operator_out3822_out1 XOR Logical_Operator_out4078_out1;

  Logical_Operator_out4975_out1 <= Logical_Operator_out3823_out1 XOR Logical_Operator_out4079_out1;

  Logical_Operator_out4976_out1 <= Logical_Operator_out3824_out1 XOR Logical_Operator_out4080_out1;

  Logical_Operator_out4977_out1 <= Logical_Operator_out3825_out1 XOR Logical_Operator_out4081_out1;

  Logical_Operator_out4978_out1 <= Logical_Operator_out3826_out1 XOR Logical_Operator_out4082_out1;

  Logical_Operator_out4979_out1 <= Logical_Operator_out3827_out1 XOR Logical_Operator_out4083_out1;

  Logical_Operator_out4980_out1 <= Logical_Operator_out3828_out1 XOR Logical_Operator_out4084_out1;

  Logical_Operator_out4981_out1 <= Logical_Operator_out3829_out1 XOR Logical_Operator_out4085_out1;

  Logical_Operator_out4982_out1 <= Logical_Operator_out3830_out1 XOR Logical_Operator_out4086_out1;

  Logical_Operator_out4983_out1 <= Logical_Operator_out3831_out1 XOR Logical_Operator_out4087_out1;

  Logical_Operator_out4984_out1 <= Logical_Operator_out3832_out1 XOR Logical_Operator_out4088_out1;

  Logical_Operator_out4985_out1 <= Logical_Operator_out3833_out1 XOR Logical_Operator_out4089_out1;

  Logical_Operator_out4986_out1 <= Logical_Operator_out3834_out1 XOR Logical_Operator_out4090_out1;

  Logical_Operator_out4987_out1 <= Logical_Operator_out3835_out1 XOR Logical_Operator_out4091_out1;

  Logical_Operator_out4988_out1 <= Logical_Operator_out3836_out1 XOR Logical_Operator_out4092_out1;

  Logical_Operator_out4989_out1 <= Logical_Operator_out3837_out1 XOR Logical_Operator_out4093_out1;

  Logical_Operator_out4990_out1 <= Logical_Operator_out3838_out1 XOR Logical_Operator_out4094_out1;

  Logical_Operator_out4991_out1 <= Logical_Operator_out3839_out1 XOR Logical_Operator_out4095_out1;

  Logical_Operator_out4992_out1 <= Logical_Operator_out3840_out1 XOR Logical_Operator_out4096_out1;

  Logical_Operator_out4993_out1 <= Logical_Operator_out3265_out1 XOR Logical_Operator_out3521_out1;

  Logical_Operator_out4994_out1 <= Logical_Operator_out3266_out1 XOR Logical_Operator_out3522_out1;

  Logical_Operator_out4995_out1 <= Logical_Operator_out3267_out1 XOR Logical_Operator_out3523_out1;

  Logical_Operator_out4996_out1 <= Logical_Operator_out3268_out1 XOR Logical_Operator_out3524_out1;

  Logical_Operator_out4997_out1 <= Logical_Operator_out3269_out1 XOR Logical_Operator_out3525_out1;

  Logical_Operator_out4998_out1 <= Logical_Operator_out3270_out1 XOR Logical_Operator_out3526_out1;

  Logical_Operator_out4999_out1 <= Logical_Operator_out3271_out1 XOR Logical_Operator_out3527_out1;

  Logical_Operator_out5000_out1 <= Logical_Operator_out3272_out1 XOR Logical_Operator_out3528_out1;

  Logical_Operator_out5001_out1 <= Logical_Operator_out3273_out1 XOR Logical_Operator_out3529_out1;

  Logical_Operator_out5002_out1 <= Logical_Operator_out3274_out1 XOR Logical_Operator_out3530_out1;

  Logical_Operator_out5003_out1 <= Logical_Operator_out3275_out1 XOR Logical_Operator_out3531_out1;

  Logical_Operator_out5004_out1 <= Logical_Operator_out3276_out1 XOR Logical_Operator_out3532_out1;

  Logical_Operator_out5005_out1 <= Logical_Operator_out3277_out1 XOR Logical_Operator_out3533_out1;

  Logical_Operator_out5006_out1 <= Logical_Operator_out3278_out1 XOR Logical_Operator_out3534_out1;

  Logical_Operator_out5007_out1 <= Logical_Operator_out3279_out1 XOR Logical_Operator_out3535_out1;

  Logical_Operator_out5008_out1 <= Logical_Operator_out3280_out1 XOR Logical_Operator_out3536_out1;

  Logical_Operator_out5009_out1 <= Logical_Operator_out3281_out1 XOR Logical_Operator_out3537_out1;

  Logical_Operator_out5010_out1 <= Logical_Operator_out3282_out1 XOR Logical_Operator_out3538_out1;

  Logical_Operator_out5011_out1 <= Logical_Operator_out3283_out1 XOR Logical_Operator_out3539_out1;

  Logical_Operator_out5012_out1 <= Logical_Operator_out3284_out1 XOR Logical_Operator_out3540_out1;

  Logical_Operator_out5013_out1 <= Logical_Operator_out3285_out1 XOR Logical_Operator_out3541_out1;

  Logical_Operator_out5014_out1 <= Logical_Operator_out3286_out1 XOR Logical_Operator_out3542_out1;

  Logical_Operator_out5015_out1 <= Logical_Operator_out3287_out1 XOR Logical_Operator_out3543_out1;

  Logical_Operator_out5016_out1 <= Logical_Operator_out3288_out1 XOR Logical_Operator_out3544_out1;

  Logical_Operator_out5017_out1 <= Logical_Operator_out3289_out1 XOR Logical_Operator_out3545_out1;

  Logical_Operator_out5018_out1 <= Logical_Operator_out3290_out1 XOR Logical_Operator_out3546_out1;

  Logical_Operator_out5019_out1 <= Logical_Operator_out3291_out1 XOR Logical_Operator_out3547_out1;

  Logical_Operator_out5020_out1 <= Logical_Operator_out3292_out1 XOR Logical_Operator_out3548_out1;

  Logical_Operator_out5021_out1 <= Logical_Operator_out3293_out1 XOR Logical_Operator_out3549_out1;

  Logical_Operator_out5022_out1 <= Logical_Operator_out3294_out1 XOR Logical_Operator_out3550_out1;

  Logical_Operator_out5023_out1 <= Logical_Operator_out3295_out1 XOR Logical_Operator_out3551_out1;

  Logical_Operator_out5024_out1 <= Logical_Operator_out3296_out1 XOR Logical_Operator_out3552_out1;

  Logical_Operator_out5025_out1 <= Logical_Operator_out3297_out1 XOR Logical_Operator_out3553_out1;

  Logical_Operator_out5026_out1 <= Logical_Operator_out3298_out1 XOR Logical_Operator_out3554_out1;

  Logical_Operator_out5027_out1 <= Logical_Operator_out3299_out1 XOR Logical_Operator_out3555_out1;

  Logical_Operator_out5028_out1 <= Logical_Operator_out3300_out1 XOR Logical_Operator_out3556_out1;

  Logical_Operator_out5029_out1 <= Logical_Operator_out3301_out1 XOR Logical_Operator_out3557_out1;

  Logical_Operator_out5030_out1 <= Logical_Operator_out3302_out1 XOR Logical_Operator_out3558_out1;

  Logical_Operator_out5031_out1 <= Logical_Operator_out3303_out1 XOR Logical_Operator_out3559_out1;

  Logical_Operator_out5032_out1 <= Logical_Operator_out3304_out1 XOR Logical_Operator_out3560_out1;

  Logical_Operator_out5033_out1 <= Logical_Operator_out3305_out1 XOR Logical_Operator_out3561_out1;

  Logical_Operator_out5034_out1 <= Logical_Operator_out3306_out1 XOR Logical_Operator_out3562_out1;

  Logical_Operator_out5035_out1 <= Logical_Operator_out3307_out1 XOR Logical_Operator_out3563_out1;

  Logical_Operator_out5036_out1 <= Logical_Operator_out3308_out1 XOR Logical_Operator_out3564_out1;

  Logical_Operator_out5037_out1 <= Logical_Operator_out3309_out1 XOR Logical_Operator_out3565_out1;

  Logical_Operator_out5038_out1 <= Logical_Operator_out3310_out1 XOR Logical_Operator_out3566_out1;

  Logical_Operator_out5039_out1 <= Logical_Operator_out3311_out1 XOR Logical_Operator_out3567_out1;

  Logical_Operator_out5040_out1 <= Logical_Operator_out3312_out1 XOR Logical_Operator_out3568_out1;

  Logical_Operator_out5041_out1 <= Logical_Operator_out3313_out1 XOR Logical_Operator_out3569_out1;

  Logical_Operator_out5042_out1 <= Logical_Operator_out3314_out1 XOR Logical_Operator_out3570_out1;

  Logical_Operator_out5043_out1 <= Logical_Operator_out3315_out1 XOR Logical_Operator_out3571_out1;

  Logical_Operator_out5044_out1 <= Logical_Operator_out3316_out1 XOR Logical_Operator_out3572_out1;

  Logical_Operator_out5045_out1 <= Logical_Operator_out3317_out1 XOR Logical_Operator_out3573_out1;

  Logical_Operator_out5046_out1 <= Logical_Operator_out3318_out1 XOR Logical_Operator_out3574_out1;

  Logical_Operator_out5047_out1 <= Logical_Operator_out3319_out1 XOR Logical_Operator_out3575_out1;

  Logical_Operator_out5048_out1 <= Logical_Operator_out3320_out1 XOR Logical_Operator_out3576_out1;

  Logical_Operator_out5049_out1 <= Logical_Operator_out3321_out1 XOR Logical_Operator_out3577_out1;

  Logical_Operator_out5050_out1 <= Logical_Operator_out3322_out1 XOR Logical_Operator_out3578_out1;

  Logical_Operator_out5051_out1 <= Logical_Operator_out3323_out1 XOR Logical_Operator_out3579_out1;

  Logical_Operator_out5052_out1 <= Logical_Operator_out3324_out1 XOR Logical_Operator_out3580_out1;

  Logical_Operator_out5053_out1 <= Logical_Operator_out3325_out1 XOR Logical_Operator_out3581_out1;

  Logical_Operator_out5054_out1 <= Logical_Operator_out3326_out1 XOR Logical_Operator_out3582_out1;

  Logical_Operator_out5055_out1 <= Logical_Operator_out3327_out1 XOR Logical_Operator_out3583_out1;

  Logical_Operator_out5056_out1 <= Logical_Operator_out3328_out1 XOR Logical_Operator_out3584_out1;

  Logical_Operator_out5057_out1 <= Logical_Operator_out2785_out1 XOR Logical_Operator_out3041_out1;

  Logical_Operator_out5058_out1 <= Logical_Operator_out2786_out1 XOR Logical_Operator_out3042_out1;

  Logical_Operator_out5059_out1 <= Logical_Operator_out2787_out1 XOR Logical_Operator_out3043_out1;

  Logical_Operator_out5060_out1 <= Logical_Operator_out2788_out1 XOR Logical_Operator_out3044_out1;

  Logical_Operator_out5061_out1 <= Logical_Operator_out2789_out1 XOR Logical_Operator_out3045_out1;

  Logical_Operator_out5062_out1 <= Logical_Operator_out2790_out1 XOR Logical_Operator_out3046_out1;

  Logical_Operator_out5063_out1 <= Logical_Operator_out2791_out1 XOR Logical_Operator_out3047_out1;

  Logical_Operator_out5064_out1 <= Logical_Operator_out2792_out1 XOR Logical_Operator_out3048_out1;

  Logical_Operator_out5065_out1 <= Logical_Operator_out2793_out1 XOR Logical_Operator_out3049_out1;

  Logical_Operator_out5066_out1 <= Logical_Operator_out2794_out1 XOR Logical_Operator_out3050_out1;

  Logical_Operator_out5067_out1 <= Logical_Operator_out2795_out1 XOR Logical_Operator_out3051_out1;

  Logical_Operator_out5068_out1 <= Logical_Operator_out2796_out1 XOR Logical_Operator_out3052_out1;

  Logical_Operator_out5069_out1 <= Logical_Operator_out2797_out1 XOR Logical_Operator_out3053_out1;

  Logical_Operator_out5070_out1 <= Logical_Operator_out2798_out1 XOR Logical_Operator_out3054_out1;

  Logical_Operator_out5071_out1 <= Logical_Operator_out2799_out1 XOR Logical_Operator_out3055_out1;

  Logical_Operator_out5072_out1 <= Logical_Operator_out2800_out1 XOR Logical_Operator_out3056_out1;

  Logical_Operator_out5073_out1 <= Logical_Operator_out2801_out1 XOR Logical_Operator_out3057_out1;

  Logical_Operator_out5074_out1 <= Logical_Operator_out2802_out1 XOR Logical_Operator_out3058_out1;

  Logical_Operator_out5075_out1 <= Logical_Operator_out2803_out1 XOR Logical_Operator_out3059_out1;

  Logical_Operator_out5076_out1 <= Logical_Operator_out2804_out1 XOR Logical_Operator_out3060_out1;

  Logical_Operator_out5077_out1 <= Logical_Operator_out2805_out1 XOR Logical_Operator_out3061_out1;

  Logical_Operator_out5078_out1 <= Logical_Operator_out2806_out1 XOR Logical_Operator_out3062_out1;

  Logical_Operator_out5079_out1 <= Logical_Operator_out2807_out1 XOR Logical_Operator_out3063_out1;

  Logical_Operator_out5080_out1 <= Logical_Operator_out2808_out1 XOR Logical_Operator_out3064_out1;

  Logical_Operator_out5081_out1 <= Logical_Operator_out2809_out1 XOR Logical_Operator_out3065_out1;

  Logical_Operator_out5082_out1 <= Logical_Operator_out2810_out1 XOR Logical_Operator_out3066_out1;

  Logical_Operator_out5083_out1 <= Logical_Operator_out2811_out1 XOR Logical_Operator_out3067_out1;

  Logical_Operator_out5084_out1 <= Logical_Operator_out2812_out1 XOR Logical_Operator_out3068_out1;

  Logical_Operator_out5085_out1 <= Logical_Operator_out2813_out1 XOR Logical_Operator_out3069_out1;

  Logical_Operator_out5086_out1 <= Logical_Operator_out2814_out1 XOR Logical_Operator_out3070_out1;

  Logical_Operator_out5087_out1 <= Logical_Operator_out2815_out1 XOR Logical_Operator_out3071_out1;

  Logical_Operator_out5088_out1 <= Logical_Operator_out2816_out1 XOR Logical_Operator_out3072_out1;

  Logical_Operator_out5089_out1 <= Logical_Operator_out2289_out1 XOR Logical_Operator_out2545_out1;

  Logical_Operator_out5090_out1 <= Logical_Operator_out2290_out1 XOR Logical_Operator_out2546_out1;

  Logical_Operator_out5091_out1 <= Logical_Operator_out2291_out1 XOR Logical_Operator_out2547_out1;

  Logical_Operator_out5092_out1 <= Logical_Operator_out2292_out1 XOR Logical_Operator_out2548_out1;

  Logical_Operator_out5093_out1 <= Logical_Operator_out2293_out1 XOR Logical_Operator_out2549_out1;

  Logical_Operator_out5094_out1 <= Logical_Operator_out2294_out1 XOR Logical_Operator_out2550_out1;

  Logical_Operator_out5095_out1 <= Logical_Operator_out2295_out1 XOR Logical_Operator_out2551_out1;

  Logical_Operator_out5096_out1 <= Logical_Operator_out2296_out1 XOR Logical_Operator_out2552_out1;

  Logical_Operator_out5097_out1 <= Logical_Operator_out2297_out1 XOR Logical_Operator_out2553_out1;

  Logical_Operator_out5098_out1 <= Logical_Operator_out2298_out1 XOR Logical_Operator_out2554_out1;

  Logical_Operator_out5099_out1 <= Logical_Operator_out2299_out1 XOR Logical_Operator_out2555_out1;

  Logical_Operator_out5100_out1 <= Logical_Operator_out2300_out1 XOR Logical_Operator_out2556_out1;

  Logical_Operator_out5101_out1 <= Logical_Operator_out2301_out1 XOR Logical_Operator_out2557_out1;

  Logical_Operator_out5102_out1 <= Logical_Operator_out2302_out1 XOR Logical_Operator_out2558_out1;

  Logical_Operator_out5103_out1 <= Logical_Operator_out2303_out1 XOR Logical_Operator_out2559_out1;

  Logical_Operator_out5104_out1 <= Logical_Operator_out2304_out1 XOR Logical_Operator_out2560_out1;

  Logical_Operator_out5105_out1 <= Logical_Operator_out1785_out1 XOR Logical_Operator_out2041_out1;

  Logical_Operator_out5106_out1 <= Logical_Operator_out1786_out1 XOR Logical_Operator_out2042_out1;

  Logical_Operator_out5107_out1 <= Logical_Operator_out1787_out1 XOR Logical_Operator_out2043_out1;

  Logical_Operator_out5108_out1 <= Logical_Operator_out1788_out1 XOR Logical_Operator_out2044_out1;

  Logical_Operator_out5109_out1 <= Logical_Operator_out1789_out1 XOR Logical_Operator_out2045_out1;

  Logical_Operator_out5110_out1 <= Logical_Operator_out1790_out1 XOR Logical_Operator_out2046_out1;

  Logical_Operator_out5111_out1 <= Logical_Operator_out1791_out1 XOR Logical_Operator_out2047_out1;

  Logical_Operator_out5112_out1 <= Logical_Operator_out1792_out1 XOR Logical_Operator_out2048_out1;

  Logical_Operator_out5113_out1 <= Logical_Operator_out1277_out1 XOR Logical_Operator_out1533_out1;

  Logical_Operator_out5114_out1 <= Logical_Operator_out1278_out1 XOR Logical_Operator_out1534_out1;

  Logical_Operator_out5115_out1 <= Logical_Operator_out1279_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out5116_out1 <= Logical_Operator_out1280_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out5117_out1 <= Logical_Operator_out767_out1 XOR Logical_Operator_out1023_out1;

  Logical_Operator_out5118_out1 <= Logical_Operator_out768_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out5119_out1 <= Logical_Operator_out256_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out5120_out1 <= in512 XOR in1024;

  out1 <= Logical_Operator_out4609_out1;

  out2 <= Logical_Operator_out4610_out1;

  out3 <= Logical_Operator_out4611_out1;

  out4 <= Logical_Operator_out4612_out1;

  out5 <= Logical_Operator_out4613_out1;

  out6 <= Logical_Operator_out4614_out1;

  out7 <= Logical_Operator_out4615_out1;

  out8 <= Logical_Operator_out4616_out1;

  out9 <= Logical_Operator_out4617_out1;

  out10 <= Logical_Operator_out4618_out1;

  out11 <= Logical_Operator_out4619_out1;

  out12 <= Logical_Operator_out4620_out1;

  out13 <= Logical_Operator_out4621_out1;

  out14 <= Logical_Operator_out4622_out1;

  out15 <= Logical_Operator_out4623_out1;

  out16 <= Logical_Operator_out4624_out1;

  out17 <= Logical_Operator_out4625_out1;

  out18 <= Logical_Operator_out4626_out1;

  out19 <= Logical_Operator_out4627_out1;

  out20 <= Logical_Operator_out4628_out1;

  out21 <= Logical_Operator_out4629_out1;

  out22 <= Logical_Operator_out4630_out1;

  out23 <= Logical_Operator_out4631_out1;

  out24 <= Logical_Operator_out4632_out1;

  out25 <= Logical_Operator_out4633_out1;

  out26 <= Logical_Operator_out4634_out1;

  out27 <= Logical_Operator_out4635_out1;

  out28 <= Logical_Operator_out4636_out1;

  out29 <= Logical_Operator_out4637_out1;

  out30 <= Logical_Operator_out4638_out1;

  out31 <= Logical_Operator_out4639_out1;

  out32 <= Logical_Operator_out4640_out1;

  out33 <= Logical_Operator_out4641_out1;

  out34 <= Logical_Operator_out4642_out1;

  out35 <= Logical_Operator_out4643_out1;

  out36 <= Logical_Operator_out4644_out1;

  out37 <= Logical_Operator_out4645_out1;

  out38 <= Logical_Operator_out4646_out1;

  out39 <= Logical_Operator_out4647_out1;

  out40 <= Logical_Operator_out4648_out1;

  out41 <= Logical_Operator_out4649_out1;

  out42 <= Logical_Operator_out4650_out1;

  out43 <= Logical_Operator_out4651_out1;

  out44 <= Logical_Operator_out4652_out1;

  out45 <= Logical_Operator_out4653_out1;

  out46 <= Logical_Operator_out4654_out1;

  out47 <= Logical_Operator_out4655_out1;

  out48 <= Logical_Operator_out4656_out1;

  out49 <= Logical_Operator_out4657_out1;

  out50 <= Logical_Operator_out4658_out1;

  out51 <= Logical_Operator_out4659_out1;

  out52 <= Logical_Operator_out4660_out1;

  out53 <= Logical_Operator_out4661_out1;

  out54 <= Logical_Operator_out4662_out1;

  out55 <= Logical_Operator_out4663_out1;

  out56 <= Logical_Operator_out4664_out1;

  out57 <= Logical_Operator_out4665_out1;

  out58 <= Logical_Operator_out4666_out1;

  out59 <= Logical_Operator_out4667_out1;

  out60 <= Logical_Operator_out4668_out1;

  out61 <= Logical_Operator_out4669_out1;

  out62 <= Logical_Operator_out4670_out1;

  out63 <= Logical_Operator_out4671_out1;

  out64 <= Logical_Operator_out4672_out1;

  out65 <= Logical_Operator_out4673_out1;

  out66 <= Logical_Operator_out4674_out1;

  out67 <= Logical_Operator_out4675_out1;

  out68 <= Logical_Operator_out4676_out1;

  out69 <= Logical_Operator_out4677_out1;

  out70 <= Logical_Operator_out4678_out1;

  out71 <= Logical_Operator_out4679_out1;

  out72 <= Logical_Operator_out4680_out1;

  out73 <= Logical_Operator_out4681_out1;

  out74 <= Logical_Operator_out4682_out1;

  out75 <= Logical_Operator_out4683_out1;

  out76 <= Logical_Operator_out4684_out1;

  out77 <= Logical_Operator_out4685_out1;

  out78 <= Logical_Operator_out4686_out1;

  out79 <= Logical_Operator_out4687_out1;

  out80 <= Logical_Operator_out4688_out1;

  out81 <= Logical_Operator_out4689_out1;

  out82 <= Logical_Operator_out4690_out1;

  out83 <= Logical_Operator_out4691_out1;

  out84 <= Logical_Operator_out4692_out1;

  out85 <= Logical_Operator_out4693_out1;

  out86 <= Logical_Operator_out4694_out1;

  out87 <= Logical_Operator_out4695_out1;

  out88 <= Logical_Operator_out4696_out1;

  out89 <= Logical_Operator_out4697_out1;

  out90 <= Logical_Operator_out4698_out1;

  out91 <= Logical_Operator_out4699_out1;

  out92 <= Logical_Operator_out4700_out1;

  out93 <= Logical_Operator_out4701_out1;

  out94 <= Logical_Operator_out4702_out1;

  out95 <= Logical_Operator_out4703_out1;

  out96 <= Logical_Operator_out4704_out1;

  out97 <= Logical_Operator_out4705_out1;

  out98 <= Logical_Operator_out4706_out1;

  out99 <= Logical_Operator_out4707_out1;

  out100 <= Logical_Operator_out4708_out1;

  out101 <= Logical_Operator_out4709_out1;

  out102 <= Logical_Operator_out4710_out1;

  out103 <= Logical_Operator_out4711_out1;

  out104 <= Logical_Operator_out4712_out1;

  out105 <= Logical_Operator_out4713_out1;

  out106 <= Logical_Operator_out4714_out1;

  out107 <= Logical_Operator_out4715_out1;

  out108 <= Logical_Operator_out4716_out1;

  out109 <= Logical_Operator_out4717_out1;

  out110 <= Logical_Operator_out4718_out1;

  out111 <= Logical_Operator_out4719_out1;

  out112 <= Logical_Operator_out4720_out1;

  out113 <= Logical_Operator_out4721_out1;

  out114 <= Logical_Operator_out4722_out1;

  out115 <= Logical_Operator_out4723_out1;

  out116 <= Logical_Operator_out4724_out1;

  out117 <= Logical_Operator_out4725_out1;

  out118 <= Logical_Operator_out4726_out1;

  out119 <= Logical_Operator_out4727_out1;

  out120 <= Logical_Operator_out4728_out1;

  out121 <= Logical_Operator_out4729_out1;

  out122 <= Logical_Operator_out4730_out1;

  out123 <= Logical_Operator_out4731_out1;

  out124 <= Logical_Operator_out4732_out1;

  out125 <= Logical_Operator_out4733_out1;

  out126 <= Logical_Operator_out4734_out1;

  out127 <= Logical_Operator_out4735_out1;

  out128 <= Logical_Operator_out4736_out1;

  out129 <= Logical_Operator_out4737_out1;

  out130 <= Logical_Operator_out4738_out1;

  out131 <= Logical_Operator_out4739_out1;

  out132 <= Logical_Operator_out4740_out1;

  out133 <= Logical_Operator_out4741_out1;

  out134 <= Logical_Operator_out4742_out1;

  out135 <= Logical_Operator_out4743_out1;

  out136 <= Logical_Operator_out4744_out1;

  out137 <= Logical_Operator_out4745_out1;

  out138 <= Logical_Operator_out4746_out1;

  out139 <= Logical_Operator_out4747_out1;

  out140 <= Logical_Operator_out4748_out1;

  out141 <= Logical_Operator_out4749_out1;

  out142 <= Logical_Operator_out4750_out1;

  out143 <= Logical_Operator_out4751_out1;

  out144 <= Logical_Operator_out4752_out1;

  out145 <= Logical_Operator_out4753_out1;

  out146 <= Logical_Operator_out4754_out1;

  out147 <= Logical_Operator_out4755_out1;

  out148 <= Logical_Operator_out4756_out1;

  out149 <= Logical_Operator_out4757_out1;

  out150 <= Logical_Operator_out4758_out1;

  out151 <= Logical_Operator_out4759_out1;

  out152 <= Logical_Operator_out4760_out1;

  out153 <= Logical_Operator_out4761_out1;

  out154 <= Logical_Operator_out4762_out1;

  out155 <= Logical_Operator_out4763_out1;

  out156 <= Logical_Operator_out4764_out1;

  out157 <= Logical_Operator_out4765_out1;

  out158 <= Logical_Operator_out4766_out1;

  out159 <= Logical_Operator_out4767_out1;

  out160 <= Logical_Operator_out4768_out1;

  out161 <= Logical_Operator_out4769_out1;

  out162 <= Logical_Operator_out4770_out1;

  out163 <= Logical_Operator_out4771_out1;

  out164 <= Logical_Operator_out4772_out1;

  out165 <= Logical_Operator_out4773_out1;

  out166 <= Logical_Operator_out4774_out1;

  out167 <= Logical_Operator_out4775_out1;

  out168 <= Logical_Operator_out4776_out1;

  out169 <= Logical_Operator_out4777_out1;

  out170 <= Logical_Operator_out4778_out1;

  out171 <= Logical_Operator_out4779_out1;

  out172 <= Logical_Operator_out4780_out1;

  out173 <= Logical_Operator_out4781_out1;

  out174 <= Logical_Operator_out4782_out1;

  out175 <= Logical_Operator_out4783_out1;

  out176 <= Logical_Operator_out4784_out1;

  out177 <= Logical_Operator_out4785_out1;

  out178 <= Logical_Operator_out4786_out1;

  out179 <= Logical_Operator_out4787_out1;

  out180 <= Logical_Operator_out4788_out1;

  out181 <= Logical_Operator_out4789_out1;

  out182 <= Logical_Operator_out4790_out1;

  out183 <= Logical_Operator_out4791_out1;

  out184 <= Logical_Operator_out4792_out1;

  out185 <= Logical_Operator_out4793_out1;

  out186 <= Logical_Operator_out4794_out1;

  out187 <= Logical_Operator_out4795_out1;

  out188 <= Logical_Operator_out4796_out1;

  out189 <= Logical_Operator_out4797_out1;

  out190 <= Logical_Operator_out4798_out1;

  out191 <= Logical_Operator_out4799_out1;

  out192 <= Logical_Operator_out4800_out1;

  out193 <= Logical_Operator_out4801_out1;

  out194 <= Logical_Operator_out4802_out1;

  out195 <= Logical_Operator_out4803_out1;

  out196 <= Logical_Operator_out4804_out1;

  out197 <= Logical_Operator_out4805_out1;

  out198 <= Logical_Operator_out4806_out1;

  out199 <= Logical_Operator_out4807_out1;

  out200 <= Logical_Operator_out4808_out1;

  out201 <= Logical_Operator_out4809_out1;

  out202 <= Logical_Operator_out4810_out1;

  out203 <= Logical_Operator_out4811_out1;

  out204 <= Logical_Operator_out4812_out1;

  out205 <= Logical_Operator_out4813_out1;

  out206 <= Logical_Operator_out4814_out1;

  out207 <= Logical_Operator_out4815_out1;

  out208 <= Logical_Operator_out4816_out1;

  out209 <= Logical_Operator_out4817_out1;

  out210 <= Logical_Operator_out4818_out1;

  out211 <= Logical_Operator_out4819_out1;

  out212 <= Logical_Operator_out4820_out1;

  out213 <= Logical_Operator_out4821_out1;

  out214 <= Logical_Operator_out4822_out1;

  out215 <= Logical_Operator_out4823_out1;

  out216 <= Logical_Operator_out4824_out1;

  out217 <= Logical_Operator_out4825_out1;

  out218 <= Logical_Operator_out4826_out1;

  out219 <= Logical_Operator_out4827_out1;

  out220 <= Logical_Operator_out4828_out1;

  out221 <= Logical_Operator_out4829_out1;

  out222 <= Logical_Operator_out4830_out1;

  out223 <= Logical_Operator_out4831_out1;

  out224 <= Logical_Operator_out4832_out1;

  out225 <= Logical_Operator_out4833_out1;

  out226 <= Logical_Operator_out4834_out1;

  out227 <= Logical_Operator_out4835_out1;

  out228 <= Logical_Operator_out4836_out1;

  out229 <= Logical_Operator_out4837_out1;

  out230 <= Logical_Operator_out4838_out1;

  out231 <= Logical_Operator_out4839_out1;

  out232 <= Logical_Operator_out4840_out1;

  out233 <= Logical_Operator_out4841_out1;

  out234 <= Logical_Operator_out4842_out1;

  out235 <= Logical_Operator_out4843_out1;

  out236 <= Logical_Operator_out4844_out1;

  out237 <= Logical_Operator_out4845_out1;

  out238 <= Logical_Operator_out4846_out1;

  out239 <= Logical_Operator_out4847_out1;

  out240 <= Logical_Operator_out4848_out1;

  out241 <= Logical_Operator_out4849_out1;

  out242 <= Logical_Operator_out4850_out1;

  out243 <= Logical_Operator_out4851_out1;

  out244 <= Logical_Operator_out4852_out1;

  out245 <= Logical_Operator_out4853_out1;

  out246 <= Logical_Operator_out4854_out1;

  out247 <= Logical_Operator_out4855_out1;

  out248 <= Logical_Operator_out4856_out1;

  out249 <= Logical_Operator_out4857_out1;

  out250 <= Logical_Operator_out4858_out1;

  out251 <= Logical_Operator_out4859_out1;

  out252 <= Logical_Operator_out4860_out1;

  out253 <= Logical_Operator_out4861_out1;

  out254 <= Logical_Operator_out4862_out1;

  out255 <= Logical_Operator_out4863_out1;

  out256 <= Logical_Operator_out4864_out1;

  out257 <= Logical_Operator_out4865_out1;

  out258 <= Logical_Operator_out4866_out1;

  out259 <= Logical_Operator_out4867_out1;

  out260 <= Logical_Operator_out4868_out1;

  out261 <= Logical_Operator_out4869_out1;

  out262 <= Logical_Operator_out4870_out1;

  out263 <= Logical_Operator_out4871_out1;

  out264 <= Logical_Operator_out4872_out1;

  out265 <= Logical_Operator_out4873_out1;

  out266 <= Logical_Operator_out4874_out1;

  out267 <= Logical_Operator_out4875_out1;

  out268 <= Logical_Operator_out4876_out1;

  out269 <= Logical_Operator_out4877_out1;

  out270 <= Logical_Operator_out4878_out1;

  out271 <= Logical_Operator_out4879_out1;

  out272 <= Logical_Operator_out4880_out1;

  out273 <= Logical_Operator_out4881_out1;

  out274 <= Logical_Operator_out4882_out1;

  out275 <= Logical_Operator_out4883_out1;

  out276 <= Logical_Operator_out4884_out1;

  out277 <= Logical_Operator_out4885_out1;

  out278 <= Logical_Operator_out4886_out1;

  out279 <= Logical_Operator_out4887_out1;

  out280 <= Logical_Operator_out4888_out1;

  out281 <= Logical_Operator_out4889_out1;

  out282 <= Logical_Operator_out4890_out1;

  out283 <= Logical_Operator_out4891_out1;

  out284 <= Logical_Operator_out4892_out1;

  out285 <= Logical_Operator_out4893_out1;

  out286 <= Logical_Operator_out4894_out1;

  out287 <= Logical_Operator_out4895_out1;

  out288 <= Logical_Operator_out4896_out1;

  out289 <= Logical_Operator_out4897_out1;

  out290 <= Logical_Operator_out4898_out1;

  out291 <= Logical_Operator_out4899_out1;

  out292 <= Logical_Operator_out4900_out1;

  out293 <= Logical_Operator_out4901_out1;

  out294 <= Logical_Operator_out4902_out1;

  out295 <= Logical_Operator_out4903_out1;

  out296 <= Logical_Operator_out4904_out1;

  out297 <= Logical_Operator_out4905_out1;

  out298 <= Logical_Operator_out4906_out1;

  out299 <= Logical_Operator_out4907_out1;

  out300 <= Logical_Operator_out4908_out1;

  out301 <= Logical_Operator_out4909_out1;

  out302 <= Logical_Operator_out4910_out1;

  out303 <= Logical_Operator_out4911_out1;

  out304 <= Logical_Operator_out4912_out1;

  out305 <= Logical_Operator_out4913_out1;

  out306 <= Logical_Operator_out4914_out1;

  out307 <= Logical_Operator_out4915_out1;

  out308 <= Logical_Operator_out4916_out1;

  out309 <= Logical_Operator_out4917_out1;

  out310 <= Logical_Operator_out4918_out1;

  out311 <= Logical_Operator_out4919_out1;

  out312 <= Logical_Operator_out4920_out1;

  out313 <= Logical_Operator_out4921_out1;

  out314 <= Logical_Operator_out4922_out1;

  out315 <= Logical_Operator_out4923_out1;

  out316 <= Logical_Operator_out4924_out1;

  out317 <= Logical_Operator_out4925_out1;

  out318 <= Logical_Operator_out4926_out1;

  out319 <= Logical_Operator_out4927_out1;

  out320 <= Logical_Operator_out4928_out1;

  out321 <= Logical_Operator_out4929_out1;

  out322 <= Logical_Operator_out4930_out1;

  out323 <= Logical_Operator_out4931_out1;

  out324 <= Logical_Operator_out4932_out1;

  out325 <= Logical_Operator_out4933_out1;

  out326 <= Logical_Operator_out4934_out1;

  out327 <= Logical_Operator_out4935_out1;

  out328 <= Logical_Operator_out4936_out1;

  out329 <= Logical_Operator_out4937_out1;

  out330 <= Logical_Operator_out4938_out1;

  out331 <= Logical_Operator_out4939_out1;

  out332 <= Logical_Operator_out4940_out1;

  out333 <= Logical_Operator_out4941_out1;

  out334 <= Logical_Operator_out4942_out1;

  out335 <= Logical_Operator_out4943_out1;

  out336 <= Logical_Operator_out4944_out1;

  out337 <= Logical_Operator_out4945_out1;

  out338 <= Logical_Operator_out4946_out1;

  out339 <= Logical_Operator_out4947_out1;

  out340 <= Logical_Operator_out4948_out1;

  out341 <= Logical_Operator_out4949_out1;

  out342 <= Logical_Operator_out4950_out1;

  out343 <= Logical_Operator_out4951_out1;

  out344 <= Logical_Operator_out4952_out1;

  out345 <= Logical_Operator_out4953_out1;

  out346 <= Logical_Operator_out4954_out1;

  out347 <= Logical_Operator_out4955_out1;

  out348 <= Logical_Operator_out4956_out1;

  out349 <= Logical_Operator_out4957_out1;

  out350 <= Logical_Operator_out4958_out1;

  out351 <= Logical_Operator_out4959_out1;

  out352 <= Logical_Operator_out4960_out1;

  out353 <= Logical_Operator_out4961_out1;

  out354 <= Logical_Operator_out4962_out1;

  out355 <= Logical_Operator_out4963_out1;

  out356 <= Logical_Operator_out4964_out1;

  out357 <= Logical_Operator_out4965_out1;

  out358 <= Logical_Operator_out4966_out1;

  out359 <= Logical_Operator_out4967_out1;

  out360 <= Logical_Operator_out4968_out1;

  out361 <= Logical_Operator_out4969_out1;

  out362 <= Logical_Operator_out4970_out1;

  out363 <= Logical_Operator_out4971_out1;

  out364 <= Logical_Operator_out4972_out1;

  out365 <= Logical_Operator_out4973_out1;

  out366 <= Logical_Operator_out4974_out1;

  out367 <= Logical_Operator_out4975_out1;

  out368 <= Logical_Operator_out4976_out1;

  out369 <= Logical_Operator_out4977_out1;

  out370 <= Logical_Operator_out4978_out1;

  out371 <= Logical_Operator_out4979_out1;

  out372 <= Logical_Operator_out4980_out1;

  out373 <= Logical_Operator_out4981_out1;

  out374 <= Logical_Operator_out4982_out1;

  out375 <= Logical_Operator_out4983_out1;

  out376 <= Logical_Operator_out4984_out1;

  out377 <= Logical_Operator_out4985_out1;

  out378 <= Logical_Operator_out4986_out1;

  out379 <= Logical_Operator_out4987_out1;

  out380 <= Logical_Operator_out4988_out1;

  out381 <= Logical_Operator_out4989_out1;

  out382 <= Logical_Operator_out4990_out1;

  out383 <= Logical_Operator_out4991_out1;

  out384 <= Logical_Operator_out4992_out1;

  out385 <= Logical_Operator_out4993_out1;

  out386 <= Logical_Operator_out4994_out1;

  out387 <= Logical_Operator_out4995_out1;

  out388 <= Logical_Operator_out4996_out1;

  out389 <= Logical_Operator_out4997_out1;

  out390 <= Logical_Operator_out4998_out1;

  out391 <= Logical_Operator_out4999_out1;

  out392 <= Logical_Operator_out5000_out1;

  out393 <= Logical_Operator_out5001_out1;

  out394 <= Logical_Operator_out5002_out1;

  out395 <= Logical_Operator_out5003_out1;

  out396 <= Logical_Operator_out5004_out1;

  out397 <= Logical_Operator_out5005_out1;

  out398 <= Logical_Operator_out5006_out1;

  out399 <= Logical_Operator_out5007_out1;

  out400 <= Logical_Operator_out5008_out1;

  out401 <= Logical_Operator_out5009_out1;

  out402 <= Logical_Operator_out5010_out1;

  out403 <= Logical_Operator_out5011_out1;

  out404 <= Logical_Operator_out5012_out1;

  out405 <= Logical_Operator_out5013_out1;

  out406 <= Logical_Operator_out5014_out1;

  out407 <= Logical_Operator_out5015_out1;

  out408 <= Logical_Operator_out5016_out1;

  out409 <= Logical_Operator_out5017_out1;

  out410 <= Logical_Operator_out5018_out1;

  out411 <= Logical_Operator_out5019_out1;

  out412 <= Logical_Operator_out5020_out1;

  out413 <= Logical_Operator_out5021_out1;

  out414 <= Logical_Operator_out5022_out1;

  out415 <= Logical_Operator_out5023_out1;

  out416 <= Logical_Operator_out5024_out1;

  out417 <= Logical_Operator_out5025_out1;

  out418 <= Logical_Operator_out5026_out1;

  out419 <= Logical_Operator_out5027_out1;

  out420 <= Logical_Operator_out5028_out1;

  out421 <= Logical_Operator_out5029_out1;

  out422 <= Logical_Operator_out5030_out1;

  out423 <= Logical_Operator_out5031_out1;

  out424 <= Logical_Operator_out5032_out1;

  out425 <= Logical_Operator_out5033_out1;

  out426 <= Logical_Operator_out5034_out1;

  out427 <= Logical_Operator_out5035_out1;

  out428 <= Logical_Operator_out5036_out1;

  out429 <= Logical_Operator_out5037_out1;

  out430 <= Logical_Operator_out5038_out1;

  out431 <= Logical_Operator_out5039_out1;

  out432 <= Logical_Operator_out5040_out1;

  out433 <= Logical_Operator_out5041_out1;

  out434 <= Logical_Operator_out5042_out1;

  out435 <= Logical_Operator_out5043_out1;

  out436 <= Logical_Operator_out5044_out1;

  out437 <= Logical_Operator_out5045_out1;

  out438 <= Logical_Operator_out5046_out1;

  out439 <= Logical_Operator_out5047_out1;

  out440 <= Logical_Operator_out5048_out1;

  out441 <= Logical_Operator_out5049_out1;

  out442 <= Logical_Operator_out5050_out1;

  out443 <= Logical_Operator_out5051_out1;

  out444 <= Logical_Operator_out5052_out1;

  out445 <= Logical_Operator_out5053_out1;

  out446 <= Logical_Operator_out5054_out1;

  out447 <= Logical_Operator_out5055_out1;

  out448 <= Logical_Operator_out5056_out1;

  out449 <= Logical_Operator_out5057_out1;

  out450 <= Logical_Operator_out5058_out1;

  out451 <= Logical_Operator_out5059_out1;

  out452 <= Logical_Operator_out5060_out1;

  out453 <= Logical_Operator_out5061_out1;

  out454 <= Logical_Operator_out5062_out1;

  out455 <= Logical_Operator_out5063_out1;

  out456 <= Logical_Operator_out5064_out1;

  out457 <= Logical_Operator_out5065_out1;

  out458 <= Logical_Operator_out5066_out1;

  out459 <= Logical_Operator_out5067_out1;

  out460 <= Logical_Operator_out5068_out1;

  out461 <= Logical_Operator_out5069_out1;

  out462 <= Logical_Operator_out5070_out1;

  out463 <= Logical_Operator_out5071_out1;

  out464 <= Logical_Operator_out5072_out1;

  out465 <= Logical_Operator_out5073_out1;

  out466 <= Logical_Operator_out5074_out1;

  out467 <= Logical_Operator_out5075_out1;

  out468 <= Logical_Operator_out5076_out1;

  out469 <= Logical_Operator_out5077_out1;

  out470 <= Logical_Operator_out5078_out1;

  out471 <= Logical_Operator_out5079_out1;

  out472 <= Logical_Operator_out5080_out1;

  out473 <= Logical_Operator_out5081_out1;

  out474 <= Logical_Operator_out5082_out1;

  out475 <= Logical_Operator_out5083_out1;

  out476 <= Logical_Operator_out5084_out1;

  out477 <= Logical_Operator_out5085_out1;

  out478 <= Logical_Operator_out5086_out1;

  out479 <= Logical_Operator_out5087_out1;

  out480 <= Logical_Operator_out5088_out1;

  out481 <= Logical_Operator_out5089_out1;

  out482 <= Logical_Operator_out5090_out1;

  out483 <= Logical_Operator_out5091_out1;

  out484 <= Logical_Operator_out5092_out1;

  out485 <= Logical_Operator_out5093_out1;

  out486 <= Logical_Operator_out5094_out1;

  out487 <= Logical_Operator_out5095_out1;

  out488 <= Logical_Operator_out5096_out1;

  out489 <= Logical_Operator_out5097_out1;

  out490 <= Logical_Operator_out5098_out1;

  out491 <= Logical_Operator_out5099_out1;

  out492 <= Logical_Operator_out5100_out1;

  out493 <= Logical_Operator_out5101_out1;

  out494 <= Logical_Operator_out5102_out1;

  out495 <= Logical_Operator_out5103_out1;

  out496 <= Logical_Operator_out5104_out1;

  out497 <= Logical_Operator_out5105_out1;

  out498 <= Logical_Operator_out5106_out1;

  out499 <= Logical_Operator_out5107_out1;

  out500 <= Logical_Operator_out5108_out1;

  out501 <= Logical_Operator_out5109_out1;

  out502 <= Logical_Operator_out5110_out1;

  out503 <= Logical_Operator_out5111_out1;

  out504 <= Logical_Operator_out5112_out1;

  out505 <= Logical_Operator_out5113_out1;

  out506 <= Logical_Operator_out5114_out1;

  out507 <= Logical_Operator_out5115_out1;

  out508 <= Logical_Operator_out5116_out1;

  out509 <= Logical_Operator_out5117_out1;

  out510 <= Logical_Operator_out5118_out1;

  out511 <= Logical_Operator_out5119_out1;

  out512 <= Logical_Operator_out5120_out1;

  out513 <= Logical_Operator_out4353_out1;

  out514 <= Logical_Operator_out4354_out1;

  out515 <= Logical_Operator_out4355_out1;

  out516 <= Logical_Operator_out4356_out1;

  out517 <= Logical_Operator_out4357_out1;

  out518 <= Logical_Operator_out4358_out1;

  out519 <= Logical_Operator_out4359_out1;

  out520 <= Logical_Operator_out4360_out1;

  out521 <= Logical_Operator_out4361_out1;

  out522 <= Logical_Operator_out4362_out1;

  out523 <= Logical_Operator_out4363_out1;

  out524 <= Logical_Operator_out4364_out1;

  out525 <= Logical_Operator_out4365_out1;

  out526 <= Logical_Operator_out4366_out1;

  out527 <= Logical_Operator_out4367_out1;

  out528 <= Logical_Operator_out4368_out1;

  out529 <= Logical_Operator_out4369_out1;

  out530 <= Logical_Operator_out4370_out1;

  out531 <= Logical_Operator_out4371_out1;

  out532 <= Logical_Operator_out4372_out1;

  out533 <= Logical_Operator_out4373_out1;

  out534 <= Logical_Operator_out4374_out1;

  out535 <= Logical_Operator_out4375_out1;

  out536 <= Logical_Operator_out4376_out1;

  out537 <= Logical_Operator_out4377_out1;

  out538 <= Logical_Operator_out4378_out1;

  out539 <= Logical_Operator_out4379_out1;

  out540 <= Logical_Operator_out4380_out1;

  out541 <= Logical_Operator_out4381_out1;

  out542 <= Logical_Operator_out4382_out1;

  out543 <= Logical_Operator_out4383_out1;

  out544 <= Logical_Operator_out4384_out1;

  out545 <= Logical_Operator_out4385_out1;

  out546 <= Logical_Operator_out4386_out1;

  out547 <= Logical_Operator_out4387_out1;

  out548 <= Logical_Operator_out4388_out1;

  out549 <= Logical_Operator_out4389_out1;

  out550 <= Logical_Operator_out4390_out1;

  out551 <= Logical_Operator_out4391_out1;

  out552 <= Logical_Operator_out4392_out1;

  out553 <= Logical_Operator_out4393_out1;

  out554 <= Logical_Operator_out4394_out1;

  out555 <= Logical_Operator_out4395_out1;

  out556 <= Logical_Operator_out4396_out1;

  out557 <= Logical_Operator_out4397_out1;

  out558 <= Logical_Operator_out4398_out1;

  out559 <= Logical_Operator_out4399_out1;

  out560 <= Logical_Operator_out4400_out1;

  out561 <= Logical_Operator_out4401_out1;

  out562 <= Logical_Operator_out4402_out1;

  out563 <= Logical_Operator_out4403_out1;

  out564 <= Logical_Operator_out4404_out1;

  out565 <= Logical_Operator_out4405_out1;

  out566 <= Logical_Operator_out4406_out1;

  out567 <= Logical_Operator_out4407_out1;

  out568 <= Logical_Operator_out4408_out1;

  out569 <= Logical_Operator_out4409_out1;

  out570 <= Logical_Operator_out4410_out1;

  out571 <= Logical_Operator_out4411_out1;

  out572 <= Logical_Operator_out4412_out1;

  out573 <= Logical_Operator_out4413_out1;

  out574 <= Logical_Operator_out4414_out1;

  out575 <= Logical_Operator_out4415_out1;

  out576 <= Logical_Operator_out4416_out1;

  out577 <= Logical_Operator_out4417_out1;

  out578 <= Logical_Operator_out4418_out1;

  out579 <= Logical_Operator_out4419_out1;

  out580 <= Logical_Operator_out4420_out1;

  out581 <= Logical_Operator_out4421_out1;

  out582 <= Logical_Operator_out4422_out1;

  out583 <= Logical_Operator_out4423_out1;

  out584 <= Logical_Operator_out4424_out1;

  out585 <= Logical_Operator_out4425_out1;

  out586 <= Logical_Operator_out4426_out1;

  out587 <= Logical_Operator_out4427_out1;

  out588 <= Logical_Operator_out4428_out1;

  out589 <= Logical_Operator_out4429_out1;

  out590 <= Logical_Operator_out4430_out1;

  out591 <= Logical_Operator_out4431_out1;

  out592 <= Logical_Operator_out4432_out1;

  out593 <= Logical_Operator_out4433_out1;

  out594 <= Logical_Operator_out4434_out1;

  out595 <= Logical_Operator_out4435_out1;

  out596 <= Logical_Operator_out4436_out1;

  out597 <= Logical_Operator_out4437_out1;

  out598 <= Logical_Operator_out4438_out1;

  out599 <= Logical_Operator_out4439_out1;

  out600 <= Logical_Operator_out4440_out1;

  out601 <= Logical_Operator_out4441_out1;

  out602 <= Logical_Operator_out4442_out1;

  out603 <= Logical_Operator_out4443_out1;

  out604 <= Logical_Operator_out4444_out1;

  out605 <= Logical_Operator_out4445_out1;

  out606 <= Logical_Operator_out4446_out1;

  out607 <= Logical_Operator_out4447_out1;

  out608 <= Logical_Operator_out4448_out1;

  out609 <= Logical_Operator_out4449_out1;

  out610 <= Logical_Operator_out4450_out1;

  out611 <= Logical_Operator_out4451_out1;

  out612 <= Logical_Operator_out4452_out1;

  out613 <= Logical_Operator_out4453_out1;

  out614 <= Logical_Operator_out4454_out1;

  out615 <= Logical_Operator_out4455_out1;

  out616 <= Logical_Operator_out4456_out1;

  out617 <= Logical_Operator_out4457_out1;

  out618 <= Logical_Operator_out4458_out1;

  out619 <= Logical_Operator_out4459_out1;

  out620 <= Logical_Operator_out4460_out1;

  out621 <= Logical_Operator_out4461_out1;

  out622 <= Logical_Operator_out4462_out1;

  out623 <= Logical_Operator_out4463_out1;

  out624 <= Logical_Operator_out4464_out1;

  out625 <= Logical_Operator_out4465_out1;

  out626 <= Logical_Operator_out4466_out1;

  out627 <= Logical_Operator_out4467_out1;

  out628 <= Logical_Operator_out4468_out1;

  out629 <= Logical_Operator_out4469_out1;

  out630 <= Logical_Operator_out4470_out1;

  out631 <= Logical_Operator_out4471_out1;

  out632 <= Logical_Operator_out4472_out1;

  out633 <= Logical_Operator_out4473_out1;

  out634 <= Logical_Operator_out4474_out1;

  out635 <= Logical_Operator_out4475_out1;

  out636 <= Logical_Operator_out4476_out1;

  out637 <= Logical_Operator_out4477_out1;

  out638 <= Logical_Operator_out4478_out1;

  out639 <= Logical_Operator_out4479_out1;

  out640 <= Logical_Operator_out4480_out1;

  out641 <= Logical_Operator_out4481_out1;

  out642 <= Logical_Operator_out4482_out1;

  out643 <= Logical_Operator_out4483_out1;

  out644 <= Logical_Operator_out4484_out1;

  out645 <= Logical_Operator_out4485_out1;

  out646 <= Logical_Operator_out4486_out1;

  out647 <= Logical_Operator_out4487_out1;

  out648 <= Logical_Operator_out4488_out1;

  out649 <= Logical_Operator_out4489_out1;

  out650 <= Logical_Operator_out4490_out1;

  out651 <= Logical_Operator_out4491_out1;

  out652 <= Logical_Operator_out4492_out1;

  out653 <= Logical_Operator_out4493_out1;

  out654 <= Logical_Operator_out4494_out1;

  out655 <= Logical_Operator_out4495_out1;

  out656 <= Logical_Operator_out4496_out1;

  out657 <= Logical_Operator_out4497_out1;

  out658 <= Logical_Operator_out4498_out1;

  out659 <= Logical_Operator_out4499_out1;

  out660 <= Logical_Operator_out4500_out1;

  out661 <= Logical_Operator_out4501_out1;

  out662 <= Logical_Operator_out4502_out1;

  out663 <= Logical_Operator_out4503_out1;

  out664 <= Logical_Operator_out4504_out1;

  out665 <= Logical_Operator_out4505_out1;

  out666 <= Logical_Operator_out4506_out1;

  out667 <= Logical_Operator_out4507_out1;

  out668 <= Logical_Operator_out4508_out1;

  out669 <= Logical_Operator_out4509_out1;

  out670 <= Logical_Operator_out4510_out1;

  out671 <= Logical_Operator_out4511_out1;

  out672 <= Logical_Operator_out4512_out1;

  out673 <= Logical_Operator_out4513_out1;

  out674 <= Logical_Operator_out4514_out1;

  out675 <= Logical_Operator_out4515_out1;

  out676 <= Logical_Operator_out4516_out1;

  out677 <= Logical_Operator_out4517_out1;

  out678 <= Logical_Operator_out4518_out1;

  out679 <= Logical_Operator_out4519_out1;

  out680 <= Logical_Operator_out4520_out1;

  out681 <= Logical_Operator_out4521_out1;

  out682 <= Logical_Operator_out4522_out1;

  out683 <= Logical_Operator_out4523_out1;

  out684 <= Logical_Operator_out4524_out1;

  out685 <= Logical_Operator_out4525_out1;

  out686 <= Logical_Operator_out4526_out1;

  out687 <= Logical_Operator_out4527_out1;

  out688 <= Logical_Operator_out4528_out1;

  out689 <= Logical_Operator_out4529_out1;

  out690 <= Logical_Operator_out4530_out1;

  out691 <= Logical_Operator_out4531_out1;

  out692 <= Logical_Operator_out4532_out1;

  out693 <= Logical_Operator_out4533_out1;

  out694 <= Logical_Operator_out4534_out1;

  out695 <= Logical_Operator_out4535_out1;

  out696 <= Logical_Operator_out4536_out1;

  out697 <= Logical_Operator_out4537_out1;

  out698 <= Logical_Operator_out4538_out1;

  out699 <= Logical_Operator_out4539_out1;

  out700 <= Logical_Operator_out4540_out1;

  out701 <= Logical_Operator_out4541_out1;

  out702 <= Logical_Operator_out4542_out1;

  out703 <= Logical_Operator_out4543_out1;

  out704 <= Logical_Operator_out4544_out1;

  out705 <= Logical_Operator_out4545_out1;

  out706 <= Logical_Operator_out4546_out1;

  out707 <= Logical_Operator_out4547_out1;

  out708 <= Logical_Operator_out4548_out1;

  out709 <= Logical_Operator_out4549_out1;

  out710 <= Logical_Operator_out4550_out1;

  out711 <= Logical_Operator_out4551_out1;

  out712 <= Logical_Operator_out4552_out1;

  out713 <= Logical_Operator_out4553_out1;

  out714 <= Logical_Operator_out4554_out1;

  out715 <= Logical_Operator_out4555_out1;

  out716 <= Logical_Operator_out4556_out1;

  out717 <= Logical_Operator_out4557_out1;

  out718 <= Logical_Operator_out4558_out1;

  out719 <= Logical_Operator_out4559_out1;

  out720 <= Logical_Operator_out4560_out1;

  out721 <= Logical_Operator_out4561_out1;

  out722 <= Logical_Operator_out4562_out1;

  out723 <= Logical_Operator_out4563_out1;

  out724 <= Logical_Operator_out4564_out1;

  out725 <= Logical_Operator_out4565_out1;

  out726 <= Logical_Operator_out4566_out1;

  out727 <= Logical_Operator_out4567_out1;

  out728 <= Logical_Operator_out4568_out1;

  out729 <= Logical_Operator_out4569_out1;

  out730 <= Logical_Operator_out4570_out1;

  out731 <= Logical_Operator_out4571_out1;

  out732 <= Logical_Operator_out4572_out1;

  out733 <= Logical_Operator_out4573_out1;

  out734 <= Logical_Operator_out4574_out1;

  out735 <= Logical_Operator_out4575_out1;

  out736 <= Logical_Operator_out4576_out1;

  out737 <= Logical_Operator_out4577_out1;

  out738 <= Logical_Operator_out4578_out1;

  out739 <= Logical_Operator_out4579_out1;

  out740 <= Logical_Operator_out4580_out1;

  out741 <= Logical_Operator_out4581_out1;

  out742 <= Logical_Operator_out4582_out1;

  out743 <= Logical_Operator_out4583_out1;

  out744 <= Logical_Operator_out4584_out1;

  out745 <= Logical_Operator_out4585_out1;

  out746 <= Logical_Operator_out4586_out1;

  out747 <= Logical_Operator_out4587_out1;

  out748 <= Logical_Operator_out4588_out1;

  out749 <= Logical_Operator_out4589_out1;

  out750 <= Logical_Operator_out4590_out1;

  out751 <= Logical_Operator_out4591_out1;

  out752 <= Logical_Operator_out4592_out1;

  out753 <= Logical_Operator_out4593_out1;

  out754 <= Logical_Operator_out4594_out1;

  out755 <= Logical_Operator_out4595_out1;

  out756 <= Logical_Operator_out4596_out1;

  out757 <= Logical_Operator_out4597_out1;

  out758 <= Logical_Operator_out4598_out1;

  out759 <= Logical_Operator_out4599_out1;

  out760 <= Logical_Operator_out4600_out1;

  out761 <= Logical_Operator_out4601_out1;

  out762 <= Logical_Operator_out4602_out1;

  out763 <= Logical_Operator_out4603_out1;

  out764 <= Logical_Operator_out4604_out1;

  out765 <= Logical_Operator_out4605_out1;

  out766 <= Logical_Operator_out4606_out1;

  out767 <= Logical_Operator_out4607_out1;

  out768 <= Logical_Operator_out4608_out1;

  out769 <= Logical_Operator_out3969_out1;

  out770 <= Logical_Operator_out3970_out1;

  out771 <= Logical_Operator_out3971_out1;

  out772 <= Logical_Operator_out3972_out1;

  out773 <= Logical_Operator_out3973_out1;

  out774 <= Logical_Operator_out3974_out1;

  out775 <= Logical_Operator_out3975_out1;

  out776 <= Logical_Operator_out3976_out1;

  out777 <= Logical_Operator_out3977_out1;

  out778 <= Logical_Operator_out3978_out1;

  out779 <= Logical_Operator_out3979_out1;

  out780 <= Logical_Operator_out3980_out1;

  out781 <= Logical_Operator_out3981_out1;

  out782 <= Logical_Operator_out3982_out1;

  out783 <= Logical_Operator_out3983_out1;

  out784 <= Logical_Operator_out3984_out1;

  out785 <= Logical_Operator_out3985_out1;

  out786 <= Logical_Operator_out3986_out1;

  out787 <= Logical_Operator_out3987_out1;

  out788 <= Logical_Operator_out3988_out1;

  out789 <= Logical_Operator_out3989_out1;

  out790 <= Logical_Operator_out3990_out1;

  out791 <= Logical_Operator_out3991_out1;

  out792 <= Logical_Operator_out3992_out1;

  out793 <= Logical_Operator_out3993_out1;

  out794 <= Logical_Operator_out3994_out1;

  out795 <= Logical_Operator_out3995_out1;

  out796 <= Logical_Operator_out3996_out1;

  out797 <= Logical_Operator_out3997_out1;

  out798 <= Logical_Operator_out3998_out1;

  out799 <= Logical_Operator_out3999_out1;

  out800 <= Logical_Operator_out4000_out1;

  out801 <= Logical_Operator_out4001_out1;

  out802 <= Logical_Operator_out4002_out1;

  out803 <= Logical_Operator_out4003_out1;

  out804 <= Logical_Operator_out4004_out1;

  out805 <= Logical_Operator_out4005_out1;

  out806 <= Logical_Operator_out4006_out1;

  out807 <= Logical_Operator_out4007_out1;

  out808 <= Logical_Operator_out4008_out1;

  out809 <= Logical_Operator_out4009_out1;

  out810 <= Logical_Operator_out4010_out1;

  out811 <= Logical_Operator_out4011_out1;

  out812 <= Logical_Operator_out4012_out1;

  out813 <= Logical_Operator_out4013_out1;

  out814 <= Logical_Operator_out4014_out1;

  out815 <= Logical_Operator_out4015_out1;

  out816 <= Logical_Operator_out4016_out1;

  out817 <= Logical_Operator_out4017_out1;

  out818 <= Logical_Operator_out4018_out1;

  out819 <= Logical_Operator_out4019_out1;

  out820 <= Logical_Operator_out4020_out1;

  out821 <= Logical_Operator_out4021_out1;

  out822 <= Logical_Operator_out4022_out1;

  out823 <= Logical_Operator_out4023_out1;

  out824 <= Logical_Operator_out4024_out1;

  out825 <= Logical_Operator_out4025_out1;

  out826 <= Logical_Operator_out4026_out1;

  out827 <= Logical_Operator_out4027_out1;

  out828 <= Logical_Operator_out4028_out1;

  out829 <= Logical_Operator_out4029_out1;

  out830 <= Logical_Operator_out4030_out1;

  out831 <= Logical_Operator_out4031_out1;

  out832 <= Logical_Operator_out4032_out1;

  out833 <= Logical_Operator_out4033_out1;

  out834 <= Logical_Operator_out4034_out1;

  out835 <= Logical_Operator_out4035_out1;

  out836 <= Logical_Operator_out4036_out1;

  out837 <= Logical_Operator_out4037_out1;

  out838 <= Logical_Operator_out4038_out1;

  out839 <= Logical_Operator_out4039_out1;

  out840 <= Logical_Operator_out4040_out1;

  out841 <= Logical_Operator_out4041_out1;

  out842 <= Logical_Operator_out4042_out1;

  out843 <= Logical_Operator_out4043_out1;

  out844 <= Logical_Operator_out4044_out1;

  out845 <= Logical_Operator_out4045_out1;

  out846 <= Logical_Operator_out4046_out1;

  out847 <= Logical_Operator_out4047_out1;

  out848 <= Logical_Operator_out4048_out1;

  out849 <= Logical_Operator_out4049_out1;

  out850 <= Logical_Operator_out4050_out1;

  out851 <= Logical_Operator_out4051_out1;

  out852 <= Logical_Operator_out4052_out1;

  out853 <= Logical_Operator_out4053_out1;

  out854 <= Logical_Operator_out4054_out1;

  out855 <= Logical_Operator_out4055_out1;

  out856 <= Logical_Operator_out4056_out1;

  out857 <= Logical_Operator_out4057_out1;

  out858 <= Logical_Operator_out4058_out1;

  out859 <= Logical_Operator_out4059_out1;

  out860 <= Logical_Operator_out4060_out1;

  out861 <= Logical_Operator_out4061_out1;

  out862 <= Logical_Operator_out4062_out1;

  out863 <= Logical_Operator_out4063_out1;

  out864 <= Logical_Operator_out4064_out1;

  out865 <= Logical_Operator_out4065_out1;

  out866 <= Logical_Operator_out4066_out1;

  out867 <= Logical_Operator_out4067_out1;

  out868 <= Logical_Operator_out4068_out1;

  out869 <= Logical_Operator_out4069_out1;

  out870 <= Logical_Operator_out4070_out1;

  out871 <= Logical_Operator_out4071_out1;

  out872 <= Logical_Operator_out4072_out1;

  out873 <= Logical_Operator_out4073_out1;

  out874 <= Logical_Operator_out4074_out1;

  out875 <= Logical_Operator_out4075_out1;

  out876 <= Logical_Operator_out4076_out1;

  out877 <= Logical_Operator_out4077_out1;

  out878 <= Logical_Operator_out4078_out1;

  out879 <= Logical_Operator_out4079_out1;

  out880 <= Logical_Operator_out4080_out1;

  out881 <= Logical_Operator_out4081_out1;

  out882 <= Logical_Operator_out4082_out1;

  out883 <= Logical_Operator_out4083_out1;

  out884 <= Logical_Operator_out4084_out1;

  out885 <= Logical_Operator_out4085_out1;

  out886 <= Logical_Operator_out4086_out1;

  out887 <= Logical_Operator_out4087_out1;

  out888 <= Logical_Operator_out4088_out1;

  out889 <= Logical_Operator_out4089_out1;

  out890 <= Logical_Operator_out4090_out1;

  out891 <= Logical_Operator_out4091_out1;

  out892 <= Logical_Operator_out4092_out1;

  out893 <= Logical_Operator_out4093_out1;

  out894 <= Logical_Operator_out4094_out1;

  out895 <= Logical_Operator_out4095_out1;

  out896 <= Logical_Operator_out4096_out1;

  out897 <= Logical_Operator_out3521_out1;

  out898 <= Logical_Operator_out3522_out1;

  out899 <= Logical_Operator_out3523_out1;

  out900 <= Logical_Operator_out3524_out1;

  out901 <= Logical_Operator_out3525_out1;

  out902 <= Logical_Operator_out3526_out1;

  out903 <= Logical_Operator_out3527_out1;

  out904 <= Logical_Operator_out3528_out1;

  out905 <= Logical_Operator_out3529_out1;

  out906 <= Logical_Operator_out3530_out1;

  out907 <= Logical_Operator_out3531_out1;

  out908 <= Logical_Operator_out3532_out1;

  out909 <= Logical_Operator_out3533_out1;

  out910 <= Logical_Operator_out3534_out1;

  out911 <= Logical_Operator_out3535_out1;

  out912 <= Logical_Operator_out3536_out1;

  out913 <= Logical_Operator_out3537_out1;

  out914 <= Logical_Operator_out3538_out1;

  out915 <= Logical_Operator_out3539_out1;

  out916 <= Logical_Operator_out3540_out1;

  out917 <= Logical_Operator_out3541_out1;

  out918 <= Logical_Operator_out3542_out1;

  out919 <= Logical_Operator_out3543_out1;

  out920 <= Logical_Operator_out3544_out1;

  out921 <= Logical_Operator_out3545_out1;

  out922 <= Logical_Operator_out3546_out1;

  out923 <= Logical_Operator_out3547_out1;

  out924 <= Logical_Operator_out3548_out1;

  out925 <= Logical_Operator_out3549_out1;

  out926 <= Logical_Operator_out3550_out1;

  out927 <= Logical_Operator_out3551_out1;

  out928 <= Logical_Operator_out3552_out1;

  out929 <= Logical_Operator_out3553_out1;

  out930 <= Logical_Operator_out3554_out1;

  out931 <= Logical_Operator_out3555_out1;

  out932 <= Logical_Operator_out3556_out1;

  out933 <= Logical_Operator_out3557_out1;

  out934 <= Logical_Operator_out3558_out1;

  out935 <= Logical_Operator_out3559_out1;

  out936 <= Logical_Operator_out3560_out1;

  out937 <= Logical_Operator_out3561_out1;

  out938 <= Logical_Operator_out3562_out1;

  out939 <= Logical_Operator_out3563_out1;

  out940 <= Logical_Operator_out3564_out1;

  out941 <= Logical_Operator_out3565_out1;

  out942 <= Logical_Operator_out3566_out1;

  out943 <= Logical_Operator_out3567_out1;

  out944 <= Logical_Operator_out3568_out1;

  out945 <= Logical_Operator_out3569_out1;

  out946 <= Logical_Operator_out3570_out1;

  out947 <= Logical_Operator_out3571_out1;

  out948 <= Logical_Operator_out3572_out1;

  out949 <= Logical_Operator_out3573_out1;

  out950 <= Logical_Operator_out3574_out1;

  out951 <= Logical_Operator_out3575_out1;

  out952 <= Logical_Operator_out3576_out1;

  out953 <= Logical_Operator_out3577_out1;

  out954 <= Logical_Operator_out3578_out1;

  out955 <= Logical_Operator_out3579_out1;

  out956 <= Logical_Operator_out3580_out1;

  out957 <= Logical_Operator_out3581_out1;

  out958 <= Logical_Operator_out3582_out1;

  out959 <= Logical_Operator_out3583_out1;

  out960 <= Logical_Operator_out3584_out1;

  out961 <= Logical_Operator_out3041_out1;

  out962 <= Logical_Operator_out3042_out1;

  out963 <= Logical_Operator_out3043_out1;

  out964 <= Logical_Operator_out3044_out1;

  out965 <= Logical_Operator_out3045_out1;

  out966 <= Logical_Operator_out3046_out1;

  out967 <= Logical_Operator_out3047_out1;

  out968 <= Logical_Operator_out3048_out1;

  out969 <= Logical_Operator_out3049_out1;

  out970 <= Logical_Operator_out3050_out1;

  out971 <= Logical_Operator_out3051_out1;

  out972 <= Logical_Operator_out3052_out1;

  out973 <= Logical_Operator_out3053_out1;

  out974 <= Logical_Operator_out3054_out1;

  out975 <= Logical_Operator_out3055_out1;

  out976 <= Logical_Operator_out3056_out1;

  out977 <= Logical_Operator_out3057_out1;

  out978 <= Logical_Operator_out3058_out1;

  out979 <= Logical_Operator_out3059_out1;

  out980 <= Logical_Operator_out3060_out1;

  out981 <= Logical_Operator_out3061_out1;

  out982 <= Logical_Operator_out3062_out1;

  out983 <= Logical_Operator_out3063_out1;

  out984 <= Logical_Operator_out3064_out1;

  out985 <= Logical_Operator_out3065_out1;

  out986 <= Logical_Operator_out3066_out1;

  out987 <= Logical_Operator_out3067_out1;

  out988 <= Logical_Operator_out3068_out1;

  out989 <= Logical_Operator_out3069_out1;

  out990 <= Logical_Operator_out3070_out1;

  out991 <= Logical_Operator_out3071_out1;

  out992 <= Logical_Operator_out3072_out1;

  out993 <= Logical_Operator_out2545_out1;

  out994 <= Logical_Operator_out2546_out1;

  out995 <= Logical_Operator_out2547_out1;

  out996 <= Logical_Operator_out2548_out1;

  out997 <= Logical_Operator_out2549_out1;

  out998 <= Logical_Operator_out2550_out1;

  out999 <= Logical_Operator_out2551_out1;

  out1000 <= Logical_Operator_out2552_out1;

  out1001 <= Logical_Operator_out2553_out1;

  out1002 <= Logical_Operator_out2554_out1;

  out1003 <= Logical_Operator_out2555_out1;

  out1004 <= Logical_Operator_out2556_out1;

  out1005 <= Logical_Operator_out2557_out1;

  out1006 <= Logical_Operator_out2558_out1;

  out1007 <= Logical_Operator_out2559_out1;

  out1008 <= Logical_Operator_out2560_out1;

  out1009 <= Logical_Operator_out2041_out1;

  out1010 <= Logical_Operator_out2042_out1;

  out1011 <= Logical_Operator_out2043_out1;

  out1012 <= Logical_Operator_out2044_out1;

  out1013 <= Logical_Operator_out2045_out1;

  out1014 <= Logical_Operator_out2046_out1;

  out1015 <= Logical_Operator_out2047_out1;

  out1016 <= Logical_Operator_out2048_out1;

  out1017 <= Logical_Operator_out1533_out1;

  out1018 <= Logical_Operator_out1534_out1;

  out1019 <= Logical_Operator_out1535_out1;

  out1020 <= Logical_Operator_out1536_out1;

  out1021 <= Logical_Operator_out1023_out1;

  out1022 <= Logical_Operator_out1024_out1;

  out1023 <= Logical_Operator_out512_out1;

  out1024 <= in1024;

END rtl;
