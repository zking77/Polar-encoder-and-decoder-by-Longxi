LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY encoderN2048 IS
PORT( 
	in1                               :   IN    std_logic;
	in2                               :   IN    std_logic;
	in3                               :   IN    std_logic;
	in4                               :   IN    std_logic;
	in5                               :   IN    std_logic;
	in6                               :   IN    std_logic;
	in7                               :   IN    std_logic;
	in8                               :   IN    std_logic;
	in9                               :   IN    std_logic;
	in10                               :   IN    std_logic;
	in11                               :   IN    std_logic;
	in12                               :   IN    std_logic;
	in13                               :   IN    std_logic;
	in14                               :   IN    std_logic;
	in15                               :   IN    std_logic;
	in16                               :   IN    std_logic;
	in17                               :   IN    std_logic;
	in18                               :   IN    std_logic;
	in19                               :   IN    std_logic;
	in20                               :   IN    std_logic;
	in21                               :   IN    std_logic;
	in22                               :   IN    std_logic;
	in23                               :   IN    std_logic;
	in24                               :   IN    std_logic;
	in25                               :   IN    std_logic;
	in26                               :   IN    std_logic;
	in27                               :   IN    std_logic;
	in28                               :   IN    std_logic;
	in29                               :   IN    std_logic;
	in30                               :   IN    std_logic;
	in31                               :   IN    std_logic;
	in32                               :   IN    std_logic;
	in33                               :   IN    std_logic;
	in34                               :   IN    std_logic;
	in35                               :   IN    std_logic;
	in36                               :   IN    std_logic;
	in37                               :   IN    std_logic;
	in38                               :   IN    std_logic;
	in39                               :   IN    std_logic;
	in40                               :   IN    std_logic;
	in41                               :   IN    std_logic;
	in42                               :   IN    std_logic;
	in43                               :   IN    std_logic;
	in44                               :   IN    std_logic;
	in45                               :   IN    std_logic;
	in46                               :   IN    std_logic;
	in47                               :   IN    std_logic;
	in48                               :   IN    std_logic;
	in49                               :   IN    std_logic;
	in50                               :   IN    std_logic;
	in51                               :   IN    std_logic;
	in52                               :   IN    std_logic;
	in53                               :   IN    std_logic;
	in54                               :   IN    std_logic;
	in55                               :   IN    std_logic;
	in56                               :   IN    std_logic;
	in57                               :   IN    std_logic;
	in58                               :   IN    std_logic;
	in59                               :   IN    std_logic;
	in60                               :   IN    std_logic;
	in61                               :   IN    std_logic;
	in62                               :   IN    std_logic;
	in63                               :   IN    std_logic;
	in64                               :   IN    std_logic;
	in65                               :   IN    std_logic;
	in66                               :   IN    std_logic;
	in67                               :   IN    std_logic;
	in68                               :   IN    std_logic;
	in69                               :   IN    std_logic;
	in70                               :   IN    std_logic;
	in71                               :   IN    std_logic;
	in72                               :   IN    std_logic;
	in73                               :   IN    std_logic;
	in74                               :   IN    std_logic;
	in75                               :   IN    std_logic;
	in76                               :   IN    std_logic;
	in77                               :   IN    std_logic;
	in78                               :   IN    std_logic;
	in79                               :   IN    std_logic;
	in80                               :   IN    std_logic;
	in81                               :   IN    std_logic;
	in82                               :   IN    std_logic;
	in83                               :   IN    std_logic;
	in84                               :   IN    std_logic;
	in85                               :   IN    std_logic;
	in86                               :   IN    std_logic;
	in87                               :   IN    std_logic;
	in88                               :   IN    std_logic;
	in89                               :   IN    std_logic;
	in90                               :   IN    std_logic;
	in91                               :   IN    std_logic;
	in92                               :   IN    std_logic;
	in93                               :   IN    std_logic;
	in94                               :   IN    std_logic;
	in95                               :   IN    std_logic;
	in96                               :   IN    std_logic;
	in97                               :   IN    std_logic;
	in98                               :   IN    std_logic;
	in99                               :   IN    std_logic;
	in100                               :   IN    std_logic;
	in101                               :   IN    std_logic;
	in102                               :   IN    std_logic;
	in103                               :   IN    std_logic;
	in104                               :   IN    std_logic;
	in105                               :   IN    std_logic;
	in106                               :   IN    std_logic;
	in107                               :   IN    std_logic;
	in108                               :   IN    std_logic;
	in109                               :   IN    std_logic;
	in110                               :   IN    std_logic;
	in111                               :   IN    std_logic;
	in112                               :   IN    std_logic;
	in113                               :   IN    std_logic;
	in114                               :   IN    std_logic;
	in115                               :   IN    std_logic;
	in116                               :   IN    std_logic;
	in117                               :   IN    std_logic;
	in118                               :   IN    std_logic;
	in119                               :   IN    std_logic;
	in120                               :   IN    std_logic;
	in121                               :   IN    std_logic;
	in122                               :   IN    std_logic;
	in123                               :   IN    std_logic;
	in124                               :   IN    std_logic;
	in125                               :   IN    std_logic;
	in126                               :   IN    std_logic;
	in127                               :   IN    std_logic;
	in128                               :   IN    std_logic;
	in129                               :   IN    std_logic;
	in130                               :   IN    std_logic;
	in131                               :   IN    std_logic;
	in132                               :   IN    std_logic;
	in133                               :   IN    std_logic;
	in134                               :   IN    std_logic;
	in135                               :   IN    std_logic;
	in136                               :   IN    std_logic;
	in137                               :   IN    std_logic;
	in138                               :   IN    std_logic;
	in139                               :   IN    std_logic;
	in140                               :   IN    std_logic;
	in141                               :   IN    std_logic;
	in142                               :   IN    std_logic;
	in143                               :   IN    std_logic;
	in144                               :   IN    std_logic;
	in145                               :   IN    std_logic;
	in146                               :   IN    std_logic;
	in147                               :   IN    std_logic;
	in148                               :   IN    std_logic;
	in149                               :   IN    std_logic;
	in150                               :   IN    std_logic;
	in151                               :   IN    std_logic;
	in152                               :   IN    std_logic;
	in153                               :   IN    std_logic;
	in154                               :   IN    std_logic;
	in155                               :   IN    std_logic;
	in156                               :   IN    std_logic;
	in157                               :   IN    std_logic;
	in158                               :   IN    std_logic;
	in159                               :   IN    std_logic;
	in160                               :   IN    std_logic;
	in161                               :   IN    std_logic;
	in162                               :   IN    std_logic;
	in163                               :   IN    std_logic;
	in164                               :   IN    std_logic;
	in165                               :   IN    std_logic;
	in166                               :   IN    std_logic;
	in167                               :   IN    std_logic;
	in168                               :   IN    std_logic;
	in169                               :   IN    std_logic;
	in170                               :   IN    std_logic;
	in171                               :   IN    std_logic;
	in172                               :   IN    std_logic;
	in173                               :   IN    std_logic;
	in174                               :   IN    std_logic;
	in175                               :   IN    std_logic;
	in176                               :   IN    std_logic;
	in177                               :   IN    std_logic;
	in178                               :   IN    std_logic;
	in179                               :   IN    std_logic;
	in180                               :   IN    std_logic;
	in181                               :   IN    std_logic;
	in182                               :   IN    std_logic;
	in183                               :   IN    std_logic;
	in184                               :   IN    std_logic;
	in185                               :   IN    std_logic;
	in186                               :   IN    std_logic;
	in187                               :   IN    std_logic;
	in188                               :   IN    std_logic;
	in189                               :   IN    std_logic;
	in190                               :   IN    std_logic;
	in191                               :   IN    std_logic;
	in192                               :   IN    std_logic;
	in193                               :   IN    std_logic;
	in194                               :   IN    std_logic;
	in195                               :   IN    std_logic;
	in196                               :   IN    std_logic;
	in197                               :   IN    std_logic;
	in198                               :   IN    std_logic;
	in199                               :   IN    std_logic;
	in200                               :   IN    std_logic;
	in201                               :   IN    std_logic;
	in202                               :   IN    std_logic;
	in203                               :   IN    std_logic;
	in204                               :   IN    std_logic;
	in205                               :   IN    std_logic;
	in206                               :   IN    std_logic;
	in207                               :   IN    std_logic;
	in208                               :   IN    std_logic;
	in209                               :   IN    std_logic;
	in210                               :   IN    std_logic;
	in211                               :   IN    std_logic;
	in212                               :   IN    std_logic;
	in213                               :   IN    std_logic;
	in214                               :   IN    std_logic;
	in215                               :   IN    std_logic;
	in216                               :   IN    std_logic;
	in217                               :   IN    std_logic;
	in218                               :   IN    std_logic;
	in219                               :   IN    std_logic;
	in220                               :   IN    std_logic;
	in221                               :   IN    std_logic;
	in222                               :   IN    std_logic;
	in223                               :   IN    std_logic;
	in224                               :   IN    std_logic;
	in225                               :   IN    std_logic;
	in226                               :   IN    std_logic;
	in227                               :   IN    std_logic;
	in228                               :   IN    std_logic;
	in229                               :   IN    std_logic;
	in230                               :   IN    std_logic;
	in231                               :   IN    std_logic;
	in232                               :   IN    std_logic;
	in233                               :   IN    std_logic;
	in234                               :   IN    std_logic;
	in235                               :   IN    std_logic;
	in236                               :   IN    std_logic;
	in237                               :   IN    std_logic;
	in238                               :   IN    std_logic;
	in239                               :   IN    std_logic;
	in240                               :   IN    std_logic;
	in241                               :   IN    std_logic;
	in242                               :   IN    std_logic;
	in243                               :   IN    std_logic;
	in244                               :   IN    std_logic;
	in245                               :   IN    std_logic;
	in246                               :   IN    std_logic;
	in247                               :   IN    std_logic;
	in248                               :   IN    std_logic;
	in249                               :   IN    std_logic;
	in250                               :   IN    std_logic;
	in251                               :   IN    std_logic;
	in252                               :   IN    std_logic;
	in253                               :   IN    std_logic;
	in254                               :   IN    std_logic;
	in255                               :   IN    std_logic;
	in256                               :   IN    std_logic;
	in257                               :   IN    std_logic;
	in258                               :   IN    std_logic;
	in259                               :   IN    std_logic;
	in260                               :   IN    std_logic;
	in261                               :   IN    std_logic;
	in262                               :   IN    std_logic;
	in263                               :   IN    std_logic;
	in264                               :   IN    std_logic;
	in265                               :   IN    std_logic;
	in266                               :   IN    std_logic;
	in267                               :   IN    std_logic;
	in268                               :   IN    std_logic;
	in269                               :   IN    std_logic;
	in270                               :   IN    std_logic;
	in271                               :   IN    std_logic;
	in272                               :   IN    std_logic;
	in273                               :   IN    std_logic;
	in274                               :   IN    std_logic;
	in275                               :   IN    std_logic;
	in276                               :   IN    std_logic;
	in277                               :   IN    std_logic;
	in278                               :   IN    std_logic;
	in279                               :   IN    std_logic;
	in280                               :   IN    std_logic;
	in281                               :   IN    std_logic;
	in282                               :   IN    std_logic;
	in283                               :   IN    std_logic;
	in284                               :   IN    std_logic;
	in285                               :   IN    std_logic;
	in286                               :   IN    std_logic;
	in287                               :   IN    std_logic;
	in288                               :   IN    std_logic;
	in289                               :   IN    std_logic;
	in290                               :   IN    std_logic;
	in291                               :   IN    std_logic;
	in292                               :   IN    std_logic;
	in293                               :   IN    std_logic;
	in294                               :   IN    std_logic;
	in295                               :   IN    std_logic;
	in296                               :   IN    std_logic;
	in297                               :   IN    std_logic;
	in298                               :   IN    std_logic;
	in299                               :   IN    std_logic;
	in300                               :   IN    std_logic;
	in301                               :   IN    std_logic;
	in302                               :   IN    std_logic;
	in303                               :   IN    std_logic;
	in304                               :   IN    std_logic;
	in305                               :   IN    std_logic;
	in306                               :   IN    std_logic;
	in307                               :   IN    std_logic;
	in308                               :   IN    std_logic;
	in309                               :   IN    std_logic;
	in310                               :   IN    std_logic;
	in311                               :   IN    std_logic;
	in312                               :   IN    std_logic;
	in313                               :   IN    std_logic;
	in314                               :   IN    std_logic;
	in315                               :   IN    std_logic;
	in316                               :   IN    std_logic;
	in317                               :   IN    std_logic;
	in318                               :   IN    std_logic;
	in319                               :   IN    std_logic;
	in320                               :   IN    std_logic;
	in321                               :   IN    std_logic;
	in322                               :   IN    std_logic;
	in323                               :   IN    std_logic;
	in324                               :   IN    std_logic;
	in325                               :   IN    std_logic;
	in326                               :   IN    std_logic;
	in327                               :   IN    std_logic;
	in328                               :   IN    std_logic;
	in329                               :   IN    std_logic;
	in330                               :   IN    std_logic;
	in331                               :   IN    std_logic;
	in332                               :   IN    std_logic;
	in333                               :   IN    std_logic;
	in334                               :   IN    std_logic;
	in335                               :   IN    std_logic;
	in336                               :   IN    std_logic;
	in337                               :   IN    std_logic;
	in338                               :   IN    std_logic;
	in339                               :   IN    std_logic;
	in340                               :   IN    std_logic;
	in341                               :   IN    std_logic;
	in342                               :   IN    std_logic;
	in343                               :   IN    std_logic;
	in344                               :   IN    std_logic;
	in345                               :   IN    std_logic;
	in346                               :   IN    std_logic;
	in347                               :   IN    std_logic;
	in348                               :   IN    std_logic;
	in349                               :   IN    std_logic;
	in350                               :   IN    std_logic;
	in351                               :   IN    std_logic;
	in352                               :   IN    std_logic;
	in353                               :   IN    std_logic;
	in354                               :   IN    std_logic;
	in355                               :   IN    std_logic;
	in356                               :   IN    std_logic;
	in357                               :   IN    std_logic;
	in358                               :   IN    std_logic;
	in359                               :   IN    std_logic;
	in360                               :   IN    std_logic;
	in361                               :   IN    std_logic;
	in362                               :   IN    std_logic;
	in363                               :   IN    std_logic;
	in364                               :   IN    std_logic;
	in365                               :   IN    std_logic;
	in366                               :   IN    std_logic;
	in367                               :   IN    std_logic;
	in368                               :   IN    std_logic;
	in369                               :   IN    std_logic;
	in370                               :   IN    std_logic;
	in371                               :   IN    std_logic;
	in372                               :   IN    std_logic;
	in373                               :   IN    std_logic;
	in374                               :   IN    std_logic;
	in375                               :   IN    std_logic;
	in376                               :   IN    std_logic;
	in377                               :   IN    std_logic;
	in378                               :   IN    std_logic;
	in379                               :   IN    std_logic;
	in380                               :   IN    std_logic;
	in381                               :   IN    std_logic;
	in382                               :   IN    std_logic;
	in383                               :   IN    std_logic;
	in384                               :   IN    std_logic;
	in385                               :   IN    std_logic;
	in386                               :   IN    std_logic;
	in387                               :   IN    std_logic;
	in388                               :   IN    std_logic;
	in389                               :   IN    std_logic;
	in390                               :   IN    std_logic;
	in391                               :   IN    std_logic;
	in392                               :   IN    std_logic;
	in393                               :   IN    std_logic;
	in394                               :   IN    std_logic;
	in395                               :   IN    std_logic;
	in396                               :   IN    std_logic;
	in397                               :   IN    std_logic;
	in398                               :   IN    std_logic;
	in399                               :   IN    std_logic;
	in400                               :   IN    std_logic;
	in401                               :   IN    std_logic;
	in402                               :   IN    std_logic;
	in403                               :   IN    std_logic;
	in404                               :   IN    std_logic;
	in405                               :   IN    std_logic;
	in406                               :   IN    std_logic;
	in407                               :   IN    std_logic;
	in408                               :   IN    std_logic;
	in409                               :   IN    std_logic;
	in410                               :   IN    std_logic;
	in411                               :   IN    std_logic;
	in412                               :   IN    std_logic;
	in413                               :   IN    std_logic;
	in414                               :   IN    std_logic;
	in415                               :   IN    std_logic;
	in416                               :   IN    std_logic;
	in417                               :   IN    std_logic;
	in418                               :   IN    std_logic;
	in419                               :   IN    std_logic;
	in420                               :   IN    std_logic;
	in421                               :   IN    std_logic;
	in422                               :   IN    std_logic;
	in423                               :   IN    std_logic;
	in424                               :   IN    std_logic;
	in425                               :   IN    std_logic;
	in426                               :   IN    std_logic;
	in427                               :   IN    std_logic;
	in428                               :   IN    std_logic;
	in429                               :   IN    std_logic;
	in430                               :   IN    std_logic;
	in431                               :   IN    std_logic;
	in432                               :   IN    std_logic;
	in433                               :   IN    std_logic;
	in434                               :   IN    std_logic;
	in435                               :   IN    std_logic;
	in436                               :   IN    std_logic;
	in437                               :   IN    std_logic;
	in438                               :   IN    std_logic;
	in439                               :   IN    std_logic;
	in440                               :   IN    std_logic;
	in441                               :   IN    std_logic;
	in442                               :   IN    std_logic;
	in443                               :   IN    std_logic;
	in444                               :   IN    std_logic;
	in445                               :   IN    std_logic;
	in446                               :   IN    std_logic;
	in447                               :   IN    std_logic;
	in448                               :   IN    std_logic;
	in449                               :   IN    std_logic;
	in450                               :   IN    std_logic;
	in451                               :   IN    std_logic;
	in452                               :   IN    std_logic;
	in453                               :   IN    std_logic;
	in454                               :   IN    std_logic;
	in455                               :   IN    std_logic;
	in456                               :   IN    std_logic;
	in457                               :   IN    std_logic;
	in458                               :   IN    std_logic;
	in459                               :   IN    std_logic;
	in460                               :   IN    std_logic;
	in461                               :   IN    std_logic;
	in462                               :   IN    std_logic;
	in463                               :   IN    std_logic;
	in464                               :   IN    std_logic;
	in465                               :   IN    std_logic;
	in466                               :   IN    std_logic;
	in467                               :   IN    std_logic;
	in468                               :   IN    std_logic;
	in469                               :   IN    std_logic;
	in470                               :   IN    std_logic;
	in471                               :   IN    std_logic;
	in472                               :   IN    std_logic;
	in473                               :   IN    std_logic;
	in474                               :   IN    std_logic;
	in475                               :   IN    std_logic;
	in476                               :   IN    std_logic;
	in477                               :   IN    std_logic;
	in478                               :   IN    std_logic;
	in479                               :   IN    std_logic;
	in480                               :   IN    std_logic;
	in481                               :   IN    std_logic;
	in482                               :   IN    std_logic;
	in483                               :   IN    std_logic;
	in484                               :   IN    std_logic;
	in485                               :   IN    std_logic;
	in486                               :   IN    std_logic;
	in487                               :   IN    std_logic;
	in488                               :   IN    std_logic;
	in489                               :   IN    std_logic;
	in490                               :   IN    std_logic;
	in491                               :   IN    std_logic;
	in492                               :   IN    std_logic;
	in493                               :   IN    std_logic;
	in494                               :   IN    std_logic;
	in495                               :   IN    std_logic;
	in496                               :   IN    std_logic;
	in497                               :   IN    std_logic;
	in498                               :   IN    std_logic;
	in499                               :   IN    std_logic;
	in500                               :   IN    std_logic;
	in501                               :   IN    std_logic;
	in502                               :   IN    std_logic;
	in503                               :   IN    std_logic;
	in504                               :   IN    std_logic;
	in505                               :   IN    std_logic;
	in506                               :   IN    std_logic;
	in507                               :   IN    std_logic;
	in508                               :   IN    std_logic;
	in509                               :   IN    std_logic;
	in510                               :   IN    std_logic;
	in511                               :   IN    std_logic;
	in512                               :   IN    std_logic;
	in513                               :   IN    std_logic;
	in514                               :   IN    std_logic;
	in515                               :   IN    std_logic;
	in516                               :   IN    std_logic;
	in517                               :   IN    std_logic;
	in518                               :   IN    std_logic;
	in519                               :   IN    std_logic;
	in520                               :   IN    std_logic;
	in521                               :   IN    std_logic;
	in522                               :   IN    std_logic;
	in523                               :   IN    std_logic;
	in524                               :   IN    std_logic;
	in525                               :   IN    std_logic;
	in526                               :   IN    std_logic;
	in527                               :   IN    std_logic;
	in528                               :   IN    std_logic;
	in529                               :   IN    std_logic;
	in530                               :   IN    std_logic;
	in531                               :   IN    std_logic;
	in532                               :   IN    std_logic;
	in533                               :   IN    std_logic;
	in534                               :   IN    std_logic;
	in535                               :   IN    std_logic;
	in536                               :   IN    std_logic;
	in537                               :   IN    std_logic;
	in538                               :   IN    std_logic;
	in539                               :   IN    std_logic;
	in540                               :   IN    std_logic;
	in541                               :   IN    std_logic;
	in542                               :   IN    std_logic;
	in543                               :   IN    std_logic;
	in544                               :   IN    std_logic;
	in545                               :   IN    std_logic;
	in546                               :   IN    std_logic;
	in547                               :   IN    std_logic;
	in548                               :   IN    std_logic;
	in549                               :   IN    std_logic;
	in550                               :   IN    std_logic;
	in551                               :   IN    std_logic;
	in552                               :   IN    std_logic;
	in553                               :   IN    std_logic;
	in554                               :   IN    std_logic;
	in555                               :   IN    std_logic;
	in556                               :   IN    std_logic;
	in557                               :   IN    std_logic;
	in558                               :   IN    std_logic;
	in559                               :   IN    std_logic;
	in560                               :   IN    std_logic;
	in561                               :   IN    std_logic;
	in562                               :   IN    std_logic;
	in563                               :   IN    std_logic;
	in564                               :   IN    std_logic;
	in565                               :   IN    std_logic;
	in566                               :   IN    std_logic;
	in567                               :   IN    std_logic;
	in568                               :   IN    std_logic;
	in569                               :   IN    std_logic;
	in570                               :   IN    std_logic;
	in571                               :   IN    std_logic;
	in572                               :   IN    std_logic;
	in573                               :   IN    std_logic;
	in574                               :   IN    std_logic;
	in575                               :   IN    std_logic;
	in576                               :   IN    std_logic;
	in577                               :   IN    std_logic;
	in578                               :   IN    std_logic;
	in579                               :   IN    std_logic;
	in580                               :   IN    std_logic;
	in581                               :   IN    std_logic;
	in582                               :   IN    std_logic;
	in583                               :   IN    std_logic;
	in584                               :   IN    std_logic;
	in585                               :   IN    std_logic;
	in586                               :   IN    std_logic;
	in587                               :   IN    std_logic;
	in588                               :   IN    std_logic;
	in589                               :   IN    std_logic;
	in590                               :   IN    std_logic;
	in591                               :   IN    std_logic;
	in592                               :   IN    std_logic;
	in593                               :   IN    std_logic;
	in594                               :   IN    std_logic;
	in595                               :   IN    std_logic;
	in596                               :   IN    std_logic;
	in597                               :   IN    std_logic;
	in598                               :   IN    std_logic;
	in599                               :   IN    std_logic;
	in600                               :   IN    std_logic;
	in601                               :   IN    std_logic;
	in602                               :   IN    std_logic;
	in603                               :   IN    std_logic;
	in604                               :   IN    std_logic;
	in605                               :   IN    std_logic;
	in606                               :   IN    std_logic;
	in607                               :   IN    std_logic;
	in608                               :   IN    std_logic;
	in609                               :   IN    std_logic;
	in610                               :   IN    std_logic;
	in611                               :   IN    std_logic;
	in612                               :   IN    std_logic;
	in613                               :   IN    std_logic;
	in614                               :   IN    std_logic;
	in615                               :   IN    std_logic;
	in616                               :   IN    std_logic;
	in617                               :   IN    std_logic;
	in618                               :   IN    std_logic;
	in619                               :   IN    std_logic;
	in620                               :   IN    std_logic;
	in621                               :   IN    std_logic;
	in622                               :   IN    std_logic;
	in623                               :   IN    std_logic;
	in624                               :   IN    std_logic;
	in625                               :   IN    std_logic;
	in626                               :   IN    std_logic;
	in627                               :   IN    std_logic;
	in628                               :   IN    std_logic;
	in629                               :   IN    std_logic;
	in630                               :   IN    std_logic;
	in631                               :   IN    std_logic;
	in632                               :   IN    std_logic;
	in633                               :   IN    std_logic;
	in634                               :   IN    std_logic;
	in635                               :   IN    std_logic;
	in636                               :   IN    std_logic;
	in637                               :   IN    std_logic;
	in638                               :   IN    std_logic;
	in639                               :   IN    std_logic;
	in640                               :   IN    std_logic;
	in641                               :   IN    std_logic;
	in642                               :   IN    std_logic;
	in643                               :   IN    std_logic;
	in644                               :   IN    std_logic;
	in645                               :   IN    std_logic;
	in646                               :   IN    std_logic;
	in647                               :   IN    std_logic;
	in648                               :   IN    std_logic;
	in649                               :   IN    std_logic;
	in650                               :   IN    std_logic;
	in651                               :   IN    std_logic;
	in652                               :   IN    std_logic;
	in653                               :   IN    std_logic;
	in654                               :   IN    std_logic;
	in655                               :   IN    std_logic;
	in656                               :   IN    std_logic;
	in657                               :   IN    std_logic;
	in658                               :   IN    std_logic;
	in659                               :   IN    std_logic;
	in660                               :   IN    std_logic;
	in661                               :   IN    std_logic;
	in662                               :   IN    std_logic;
	in663                               :   IN    std_logic;
	in664                               :   IN    std_logic;
	in665                               :   IN    std_logic;
	in666                               :   IN    std_logic;
	in667                               :   IN    std_logic;
	in668                               :   IN    std_logic;
	in669                               :   IN    std_logic;
	in670                               :   IN    std_logic;
	in671                               :   IN    std_logic;
	in672                               :   IN    std_logic;
	in673                               :   IN    std_logic;
	in674                               :   IN    std_logic;
	in675                               :   IN    std_logic;
	in676                               :   IN    std_logic;
	in677                               :   IN    std_logic;
	in678                               :   IN    std_logic;
	in679                               :   IN    std_logic;
	in680                               :   IN    std_logic;
	in681                               :   IN    std_logic;
	in682                               :   IN    std_logic;
	in683                               :   IN    std_logic;
	in684                               :   IN    std_logic;
	in685                               :   IN    std_logic;
	in686                               :   IN    std_logic;
	in687                               :   IN    std_logic;
	in688                               :   IN    std_logic;
	in689                               :   IN    std_logic;
	in690                               :   IN    std_logic;
	in691                               :   IN    std_logic;
	in692                               :   IN    std_logic;
	in693                               :   IN    std_logic;
	in694                               :   IN    std_logic;
	in695                               :   IN    std_logic;
	in696                               :   IN    std_logic;
	in697                               :   IN    std_logic;
	in698                               :   IN    std_logic;
	in699                               :   IN    std_logic;
	in700                               :   IN    std_logic;
	in701                               :   IN    std_logic;
	in702                               :   IN    std_logic;
	in703                               :   IN    std_logic;
	in704                               :   IN    std_logic;
	in705                               :   IN    std_logic;
	in706                               :   IN    std_logic;
	in707                               :   IN    std_logic;
	in708                               :   IN    std_logic;
	in709                               :   IN    std_logic;
	in710                               :   IN    std_logic;
	in711                               :   IN    std_logic;
	in712                               :   IN    std_logic;
	in713                               :   IN    std_logic;
	in714                               :   IN    std_logic;
	in715                               :   IN    std_logic;
	in716                               :   IN    std_logic;
	in717                               :   IN    std_logic;
	in718                               :   IN    std_logic;
	in719                               :   IN    std_logic;
	in720                               :   IN    std_logic;
	in721                               :   IN    std_logic;
	in722                               :   IN    std_logic;
	in723                               :   IN    std_logic;
	in724                               :   IN    std_logic;
	in725                               :   IN    std_logic;
	in726                               :   IN    std_logic;
	in727                               :   IN    std_logic;
	in728                               :   IN    std_logic;
	in729                               :   IN    std_logic;
	in730                               :   IN    std_logic;
	in731                               :   IN    std_logic;
	in732                               :   IN    std_logic;
	in733                               :   IN    std_logic;
	in734                               :   IN    std_logic;
	in735                               :   IN    std_logic;
	in736                               :   IN    std_logic;
	in737                               :   IN    std_logic;
	in738                               :   IN    std_logic;
	in739                               :   IN    std_logic;
	in740                               :   IN    std_logic;
	in741                               :   IN    std_logic;
	in742                               :   IN    std_logic;
	in743                               :   IN    std_logic;
	in744                               :   IN    std_logic;
	in745                               :   IN    std_logic;
	in746                               :   IN    std_logic;
	in747                               :   IN    std_logic;
	in748                               :   IN    std_logic;
	in749                               :   IN    std_logic;
	in750                               :   IN    std_logic;
	in751                               :   IN    std_logic;
	in752                               :   IN    std_logic;
	in753                               :   IN    std_logic;
	in754                               :   IN    std_logic;
	in755                               :   IN    std_logic;
	in756                               :   IN    std_logic;
	in757                               :   IN    std_logic;
	in758                               :   IN    std_logic;
	in759                               :   IN    std_logic;
	in760                               :   IN    std_logic;
	in761                               :   IN    std_logic;
	in762                               :   IN    std_logic;
	in763                               :   IN    std_logic;
	in764                               :   IN    std_logic;
	in765                               :   IN    std_logic;
	in766                               :   IN    std_logic;
	in767                               :   IN    std_logic;
	in768                               :   IN    std_logic;
	in769                               :   IN    std_logic;
	in770                               :   IN    std_logic;
	in771                               :   IN    std_logic;
	in772                               :   IN    std_logic;
	in773                               :   IN    std_logic;
	in774                               :   IN    std_logic;
	in775                               :   IN    std_logic;
	in776                               :   IN    std_logic;
	in777                               :   IN    std_logic;
	in778                               :   IN    std_logic;
	in779                               :   IN    std_logic;
	in780                               :   IN    std_logic;
	in781                               :   IN    std_logic;
	in782                               :   IN    std_logic;
	in783                               :   IN    std_logic;
	in784                               :   IN    std_logic;
	in785                               :   IN    std_logic;
	in786                               :   IN    std_logic;
	in787                               :   IN    std_logic;
	in788                               :   IN    std_logic;
	in789                               :   IN    std_logic;
	in790                               :   IN    std_logic;
	in791                               :   IN    std_logic;
	in792                               :   IN    std_logic;
	in793                               :   IN    std_logic;
	in794                               :   IN    std_logic;
	in795                               :   IN    std_logic;
	in796                               :   IN    std_logic;
	in797                               :   IN    std_logic;
	in798                               :   IN    std_logic;
	in799                               :   IN    std_logic;
	in800                               :   IN    std_logic;
	in801                               :   IN    std_logic;
	in802                               :   IN    std_logic;
	in803                               :   IN    std_logic;
	in804                               :   IN    std_logic;
	in805                               :   IN    std_logic;
	in806                               :   IN    std_logic;
	in807                               :   IN    std_logic;
	in808                               :   IN    std_logic;
	in809                               :   IN    std_logic;
	in810                               :   IN    std_logic;
	in811                               :   IN    std_logic;
	in812                               :   IN    std_logic;
	in813                               :   IN    std_logic;
	in814                               :   IN    std_logic;
	in815                               :   IN    std_logic;
	in816                               :   IN    std_logic;
	in817                               :   IN    std_logic;
	in818                               :   IN    std_logic;
	in819                               :   IN    std_logic;
	in820                               :   IN    std_logic;
	in821                               :   IN    std_logic;
	in822                               :   IN    std_logic;
	in823                               :   IN    std_logic;
	in824                               :   IN    std_logic;
	in825                               :   IN    std_logic;
	in826                               :   IN    std_logic;
	in827                               :   IN    std_logic;
	in828                               :   IN    std_logic;
	in829                               :   IN    std_logic;
	in830                               :   IN    std_logic;
	in831                               :   IN    std_logic;
	in832                               :   IN    std_logic;
	in833                               :   IN    std_logic;
	in834                               :   IN    std_logic;
	in835                               :   IN    std_logic;
	in836                               :   IN    std_logic;
	in837                               :   IN    std_logic;
	in838                               :   IN    std_logic;
	in839                               :   IN    std_logic;
	in840                               :   IN    std_logic;
	in841                               :   IN    std_logic;
	in842                               :   IN    std_logic;
	in843                               :   IN    std_logic;
	in844                               :   IN    std_logic;
	in845                               :   IN    std_logic;
	in846                               :   IN    std_logic;
	in847                               :   IN    std_logic;
	in848                               :   IN    std_logic;
	in849                               :   IN    std_logic;
	in850                               :   IN    std_logic;
	in851                               :   IN    std_logic;
	in852                               :   IN    std_logic;
	in853                               :   IN    std_logic;
	in854                               :   IN    std_logic;
	in855                               :   IN    std_logic;
	in856                               :   IN    std_logic;
	in857                               :   IN    std_logic;
	in858                               :   IN    std_logic;
	in859                               :   IN    std_logic;
	in860                               :   IN    std_logic;
	in861                               :   IN    std_logic;
	in862                               :   IN    std_logic;
	in863                               :   IN    std_logic;
	in864                               :   IN    std_logic;
	in865                               :   IN    std_logic;
	in866                               :   IN    std_logic;
	in867                               :   IN    std_logic;
	in868                               :   IN    std_logic;
	in869                               :   IN    std_logic;
	in870                               :   IN    std_logic;
	in871                               :   IN    std_logic;
	in872                               :   IN    std_logic;
	in873                               :   IN    std_logic;
	in874                               :   IN    std_logic;
	in875                               :   IN    std_logic;
	in876                               :   IN    std_logic;
	in877                               :   IN    std_logic;
	in878                               :   IN    std_logic;
	in879                               :   IN    std_logic;
	in880                               :   IN    std_logic;
	in881                               :   IN    std_logic;
	in882                               :   IN    std_logic;
	in883                               :   IN    std_logic;
	in884                               :   IN    std_logic;
	in885                               :   IN    std_logic;
	in886                               :   IN    std_logic;
	in887                               :   IN    std_logic;
	in888                               :   IN    std_logic;
	in889                               :   IN    std_logic;
	in890                               :   IN    std_logic;
	in891                               :   IN    std_logic;
	in892                               :   IN    std_logic;
	in893                               :   IN    std_logic;
	in894                               :   IN    std_logic;
	in895                               :   IN    std_logic;
	in896                               :   IN    std_logic;
	in897                               :   IN    std_logic;
	in898                               :   IN    std_logic;
	in899                               :   IN    std_logic;
	in900                               :   IN    std_logic;
	in901                               :   IN    std_logic;
	in902                               :   IN    std_logic;
	in903                               :   IN    std_logic;
	in904                               :   IN    std_logic;
	in905                               :   IN    std_logic;
	in906                               :   IN    std_logic;
	in907                               :   IN    std_logic;
	in908                               :   IN    std_logic;
	in909                               :   IN    std_logic;
	in910                               :   IN    std_logic;
	in911                               :   IN    std_logic;
	in912                               :   IN    std_logic;
	in913                               :   IN    std_logic;
	in914                               :   IN    std_logic;
	in915                               :   IN    std_logic;
	in916                               :   IN    std_logic;
	in917                               :   IN    std_logic;
	in918                               :   IN    std_logic;
	in919                               :   IN    std_logic;
	in920                               :   IN    std_logic;
	in921                               :   IN    std_logic;
	in922                               :   IN    std_logic;
	in923                               :   IN    std_logic;
	in924                               :   IN    std_logic;
	in925                               :   IN    std_logic;
	in926                               :   IN    std_logic;
	in927                               :   IN    std_logic;
	in928                               :   IN    std_logic;
	in929                               :   IN    std_logic;
	in930                               :   IN    std_logic;
	in931                               :   IN    std_logic;
	in932                               :   IN    std_logic;
	in933                               :   IN    std_logic;
	in934                               :   IN    std_logic;
	in935                               :   IN    std_logic;
	in936                               :   IN    std_logic;
	in937                               :   IN    std_logic;
	in938                               :   IN    std_logic;
	in939                               :   IN    std_logic;
	in940                               :   IN    std_logic;
	in941                               :   IN    std_logic;
	in942                               :   IN    std_logic;
	in943                               :   IN    std_logic;
	in944                               :   IN    std_logic;
	in945                               :   IN    std_logic;
	in946                               :   IN    std_logic;
	in947                               :   IN    std_logic;
	in948                               :   IN    std_logic;
	in949                               :   IN    std_logic;
	in950                               :   IN    std_logic;
	in951                               :   IN    std_logic;
	in952                               :   IN    std_logic;
	in953                               :   IN    std_logic;
	in954                               :   IN    std_logic;
	in955                               :   IN    std_logic;
	in956                               :   IN    std_logic;
	in957                               :   IN    std_logic;
	in958                               :   IN    std_logic;
	in959                               :   IN    std_logic;
	in960                               :   IN    std_logic;
	in961                               :   IN    std_logic;
	in962                               :   IN    std_logic;
	in963                               :   IN    std_logic;
	in964                               :   IN    std_logic;
	in965                               :   IN    std_logic;
	in966                               :   IN    std_logic;
	in967                               :   IN    std_logic;
	in968                               :   IN    std_logic;
	in969                               :   IN    std_logic;
	in970                               :   IN    std_logic;
	in971                               :   IN    std_logic;
	in972                               :   IN    std_logic;
	in973                               :   IN    std_logic;
	in974                               :   IN    std_logic;
	in975                               :   IN    std_logic;
	in976                               :   IN    std_logic;
	in977                               :   IN    std_logic;
	in978                               :   IN    std_logic;
	in979                               :   IN    std_logic;
	in980                               :   IN    std_logic;
	in981                               :   IN    std_logic;
	in982                               :   IN    std_logic;
	in983                               :   IN    std_logic;
	in984                               :   IN    std_logic;
	in985                               :   IN    std_logic;
	in986                               :   IN    std_logic;
	in987                               :   IN    std_logic;
	in988                               :   IN    std_logic;
	in989                               :   IN    std_logic;
	in990                               :   IN    std_logic;
	in991                               :   IN    std_logic;
	in992                               :   IN    std_logic;
	in993                               :   IN    std_logic;
	in994                               :   IN    std_logic;
	in995                               :   IN    std_logic;
	in996                               :   IN    std_logic;
	in997                               :   IN    std_logic;
	in998                               :   IN    std_logic;
	in999                               :   IN    std_logic;
	in1000                               :   IN    std_logic;
	in1001                               :   IN    std_logic;
	in1002                               :   IN    std_logic;
	in1003                               :   IN    std_logic;
	in1004                               :   IN    std_logic;
	in1005                               :   IN    std_logic;
	in1006                               :   IN    std_logic;
	in1007                               :   IN    std_logic;
	in1008                               :   IN    std_logic;
	in1009                               :   IN    std_logic;
	in1010                               :   IN    std_logic;
	in1011                               :   IN    std_logic;
	in1012                               :   IN    std_logic;
	in1013                               :   IN    std_logic;
	in1014                               :   IN    std_logic;
	in1015                               :   IN    std_logic;
	in1016                               :   IN    std_logic;
	in1017                               :   IN    std_logic;
	in1018                               :   IN    std_logic;
	in1019                               :   IN    std_logic;
	in1020                               :   IN    std_logic;
	in1021                               :   IN    std_logic;
	in1022                               :   IN    std_logic;
	in1023                               :   IN    std_logic;
	in1024                               :   IN    std_logic;
	in1025                               :   IN    std_logic;
	in1026                               :   IN    std_logic;
	in1027                               :   IN    std_logic;
	in1028                               :   IN    std_logic;
	in1029                               :   IN    std_logic;
	in1030                               :   IN    std_logic;
	in1031                               :   IN    std_logic;
	in1032                               :   IN    std_logic;
	in1033                               :   IN    std_logic;
	in1034                               :   IN    std_logic;
	in1035                               :   IN    std_logic;
	in1036                               :   IN    std_logic;
	in1037                               :   IN    std_logic;
	in1038                               :   IN    std_logic;
	in1039                               :   IN    std_logic;
	in1040                               :   IN    std_logic;
	in1041                               :   IN    std_logic;
	in1042                               :   IN    std_logic;
	in1043                               :   IN    std_logic;
	in1044                               :   IN    std_logic;
	in1045                               :   IN    std_logic;
	in1046                               :   IN    std_logic;
	in1047                               :   IN    std_logic;
	in1048                               :   IN    std_logic;
	in1049                               :   IN    std_logic;
	in1050                               :   IN    std_logic;
	in1051                               :   IN    std_logic;
	in1052                               :   IN    std_logic;
	in1053                               :   IN    std_logic;
	in1054                               :   IN    std_logic;
	in1055                               :   IN    std_logic;
	in1056                               :   IN    std_logic;
	in1057                               :   IN    std_logic;
	in1058                               :   IN    std_logic;
	in1059                               :   IN    std_logic;
	in1060                               :   IN    std_logic;
	in1061                               :   IN    std_logic;
	in1062                               :   IN    std_logic;
	in1063                               :   IN    std_logic;
	in1064                               :   IN    std_logic;
	in1065                               :   IN    std_logic;
	in1066                               :   IN    std_logic;
	in1067                               :   IN    std_logic;
	in1068                               :   IN    std_logic;
	in1069                               :   IN    std_logic;
	in1070                               :   IN    std_logic;
	in1071                               :   IN    std_logic;
	in1072                               :   IN    std_logic;
	in1073                               :   IN    std_logic;
	in1074                               :   IN    std_logic;
	in1075                               :   IN    std_logic;
	in1076                               :   IN    std_logic;
	in1077                               :   IN    std_logic;
	in1078                               :   IN    std_logic;
	in1079                               :   IN    std_logic;
	in1080                               :   IN    std_logic;
	in1081                               :   IN    std_logic;
	in1082                               :   IN    std_logic;
	in1083                               :   IN    std_logic;
	in1084                               :   IN    std_logic;
	in1085                               :   IN    std_logic;
	in1086                               :   IN    std_logic;
	in1087                               :   IN    std_logic;
	in1088                               :   IN    std_logic;
	in1089                               :   IN    std_logic;
	in1090                               :   IN    std_logic;
	in1091                               :   IN    std_logic;
	in1092                               :   IN    std_logic;
	in1093                               :   IN    std_logic;
	in1094                               :   IN    std_logic;
	in1095                               :   IN    std_logic;
	in1096                               :   IN    std_logic;
	in1097                               :   IN    std_logic;
	in1098                               :   IN    std_logic;
	in1099                               :   IN    std_logic;
	in1100                               :   IN    std_logic;
	in1101                               :   IN    std_logic;
	in1102                               :   IN    std_logic;
	in1103                               :   IN    std_logic;
	in1104                               :   IN    std_logic;
	in1105                               :   IN    std_logic;
	in1106                               :   IN    std_logic;
	in1107                               :   IN    std_logic;
	in1108                               :   IN    std_logic;
	in1109                               :   IN    std_logic;
	in1110                               :   IN    std_logic;
	in1111                               :   IN    std_logic;
	in1112                               :   IN    std_logic;
	in1113                               :   IN    std_logic;
	in1114                               :   IN    std_logic;
	in1115                               :   IN    std_logic;
	in1116                               :   IN    std_logic;
	in1117                               :   IN    std_logic;
	in1118                               :   IN    std_logic;
	in1119                               :   IN    std_logic;
	in1120                               :   IN    std_logic;
	in1121                               :   IN    std_logic;
	in1122                               :   IN    std_logic;
	in1123                               :   IN    std_logic;
	in1124                               :   IN    std_logic;
	in1125                               :   IN    std_logic;
	in1126                               :   IN    std_logic;
	in1127                               :   IN    std_logic;
	in1128                               :   IN    std_logic;
	in1129                               :   IN    std_logic;
	in1130                               :   IN    std_logic;
	in1131                               :   IN    std_logic;
	in1132                               :   IN    std_logic;
	in1133                               :   IN    std_logic;
	in1134                               :   IN    std_logic;
	in1135                               :   IN    std_logic;
	in1136                               :   IN    std_logic;
	in1137                               :   IN    std_logic;
	in1138                               :   IN    std_logic;
	in1139                               :   IN    std_logic;
	in1140                               :   IN    std_logic;
	in1141                               :   IN    std_logic;
	in1142                               :   IN    std_logic;
	in1143                               :   IN    std_logic;
	in1144                               :   IN    std_logic;
	in1145                               :   IN    std_logic;
	in1146                               :   IN    std_logic;
	in1147                               :   IN    std_logic;
	in1148                               :   IN    std_logic;
	in1149                               :   IN    std_logic;
	in1150                               :   IN    std_logic;
	in1151                               :   IN    std_logic;
	in1152                               :   IN    std_logic;
	in1153                               :   IN    std_logic;
	in1154                               :   IN    std_logic;
	in1155                               :   IN    std_logic;
	in1156                               :   IN    std_logic;
	in1157                               :   IN    std_logic;
	in1158                               :   IN    std_logic;
	in1159                               :   IN    std_logic;
	in1160                               :   IN    std_logic;
	in1161                               :   IN    std_logic;
	in1162                               :   IN    std_logic;
	in1163                               :   IN    std_logic;
	in1164                               :   IN    std_logic;
	in1165                               :   IN    std_logic;
	in1166                               :   IN    std_logic;
	in1167                               :   IN    std_logic;
	in1168                               :   IN    std_logic;
	in1169                               :   IN    std_logic;
	in1170                               :   IN    std_logic;
	in1171                               :   IN    std_logic;
	in1172                               :   IN    std_logic;
	in1173                               :   IN    std_logic;
	in1174                               :   IN    std_logic;
	in1175                               :   IN    std_logic;
	in1176                               :   IN    std_logic;
	in1177                               :   IN    std_logic;
	in1178                               :   IN    std_logic;
	in1179                               :   IN    std_logic;
	in1180                               :   IN    std_logic;
	in1181                               :   IN    std_logic;
	in1182                               :   IN    std_logic;
	in1183                               :   IN    std_logic;
	in1184                               :   IN    std_logic;
	in1185                               :   IN    std_logic;
	in1186                               :   IN    std_logic;
	in1187                               :   IN    std_logic;
	in1188                               :   IN    std_logic;
	in1189                               :   IN    std_logic;
	in1190                               :   IN    std_logic;
	in1191                               :   IN    std_logic;
	in1192                               :   IN    std_logic;
	in1193                               :   IN    std_logic;
	in1194                               :   IN    std_logic;
	in1195                               :   IN    std_logic;
	in1196                               :   IN    std_logic;
	in1197                               :   IN    std_logic;
	in1198                               :   IN    std_logic;
	in1199                               :   IN    std_logic;
	in1200                               :   IN    std_logic;
	in1201                               :   IN    std_logic;
	in1202                               :   IN    std_logic;
	in1203                               :   IN    std_logic;
	in1204                               :   IN    std_logic;
	in1205                               :   IN    std_logic;
	in1206                               :   IN    std_logic;
	in1207                               :   IN    std_logic;
	in1208                               :   IN    std_logic;
	in1209                               :   IN    std_logic;
	in1210                               :   IN    std_logic;
	in1211                               :   IN    std_logic;
	in1212                               :   IN    std_logic;
	in1213                               :   IN    std_logic;
	in1214                               :   IN    std_logic;
	in1215                               :   IN    std_logic;
	in1216                               :   IN    std_logic;
	in1217                               :   IN    std_logic;
	in1218                               :   IN    std_logic;
	in1219                               :   IN    std_logic;
	in1220                               :   IN    std_logic;
	in1221                               :   IN    std_logic;
	in1222                               :   IN    std_logic;
	in1223                               :   IN    std_logic;
	in1224                               :   IN    std_logic;
	in1225                               :   IN    std_logic;
	in1226                               :   IN    std_logic;
	in1227                               :   IN    std_logic;
	in1228                               :   IN    std_logic;
	in1229                               :   IN    std_logic;
	in1230                               :   IN    std_logic;
	in1231                               :   IN    std_logic;
	in1232                               :   IN    std_logic;
	in1233                               :   IN    std_logic;
	in1234                               :   IN    std_logic;
	in1235                               :   IN    std_logic;
	in1236                               :   IN    std_logic;
	in1237                               :   IN    std_logic;
	in1238                               :   IN    std_logic;
	in1239                               :   IN    std_logic;
	in1240                               :   IN    std_logic;
	in1241                               :   IN    std_logic;
	in1242                               :   IN    std_logic;
	in1243                               :   IN    std_logic;
	in1244                               :   IN    std_logic;
	in1245                               :   IN    std_logic;
	in1246                               :   IN    std_logic;
	in1247                               :   IN    std_logic;
	in1248                               :   IN    std_logic;
	in1249                               :   IN    std_logic;
	in1250                               :   IN    std_logic;
	in1251                               :   IN    std_logic;
	in1252                               :   IN    std_logic;
	in1253                               :   IN    std_logic;
	in1254                               :   IN    std_logic;
	in1255                               :   IN    std_logic;
	in1256                               :   IN    std_logic;
	in1257                               :   IN    std_logic;
	in1258                               :   IN    std_logic;
	in1259                               :   IN    std_logic;
	in1260                               :   IN    std_logic;
	in1261                               :   IN    std_logic;
	in1262                               :   IN    std_logic;
	in1263                               :   IN    std_logic;
	in1264                               :   IN    std_logic;
	in1265                               :   IN    std_logic;
	in1266                               :   IN    std_logic;
	in1267                               :   IN    std_logic;
	in1268                               :   IN    std_logic;
	in1269                               :   IN    std_logic;
	in1270                               :   IN    std_logic;
	in1271                               :   IN    std_logic;
	in1272                               :   IN    std_logic;
	in1273                               :   IN    std_logic;
	in1274                               :   IN    std_logic;
	in1275                               :   IN    std_logic;
	in1276                               :   IN    std_logic;
	in1277                               :   IN    std_logic;
	in1278                               :   IN    std_logic;
	in1279                               :   IN    std_logic;
	in1280                               :   IN    std_logic;
	in1281                               :   IN    std_logic;
	in1282                               :   IN    std_logic;
	in1283                               :   IN    std_logic;
	in1284                               :   IN    std_logic;
	in1285                               :   IN    std_logic;
	in1286                               :   IN    std_logic;
	in1287                               :   IN    std_logic;
	in1288                               :   IN    std_logic;
	in1289                               :   IN    std_logic;
	in1290                               :   IN    std_logic;
	in1291                               :   IN    std_logic;
	in1292                               :   IN    std_logic;
	in1293                               :   IN    std_logic;
	in1294                               :   IN    std_logic;
	in1295                               :   IN    std_logic;
	in1296                               :   IN    std_logic;
	in1297                               :   IN    std_logic;
	in1298                               :   IN    std_logic;
	in1299                               :   IN    std_logic;
	in1300                               :   IN    std_logic;
	in1301                               :   IN    std_logic;
	in1302                               :   IN    std_logic;
	in1303                               :   IN    std_logic;
	in1304                               :   IN    std_logic;
	in1305                               :   IN    std_logic;
	in1306                               :   IN    std_logic;
	in1307                               :   IN    std_logic;
	in1308                               :   IN    std_logic;
	in1309                               :   IN    std_logic;
	in1310                               :   IN    std_logic;
	in1311                               :   IN    std_logic;
	in1312                               :   IN    std_logic;
	in1313                               :   IN    std_logic;
	in1314                               :   IN    std_logic;
	in1315                               :   IN    std_logic;
	in1316                               :   IN    std_logic;
	in1317                               :   IN    std_logic;
	in1318                               :   IN    std_logic;
	in1319                               :   IN    std_logic;
	in1320                               :   IN    std_logic;
	in1321                               :   IN    std_logic;
	in1322                               :   IN    std_logic;
	in1323                               :   IN    std_logic;
	in1324                               :   IN    std_logic;
	in1325                               :   IN    std_logic;
	in1326                               :   IN    std_logic;
	in1327                               :   IN    std_logic;
	in1328                               :   IN    std_logic;
	in1329                               :   IN    std_logic;
	in1330                               :   IN    std_logic;
	in1331                               :   IN    std_logic;
	in1332                               :   IN    std_logic;
	in1333                               :   IN    std_logic;
	in1334                               :   IN    std_logic;
	in1335                               :   IN    std_logic;
	in1336                               :   IN    std_logic;
	in1337                               :   IN    std_logic;
	in1338                               :   IN    std_logic;
	in1339                               :   IN    std_logic;
	in1340                               :   IN    std_logic;
	in1341                               :   IN    std_logic;
	in1342                               :   IN    std_logic;
	in1343                               :   IN    std_logic;
	in1344                               :   IN    std_logic;
	in1345                               :   IN    std_logic;
	in1346                               :   IN    std_logic;
	in1347                               :   IN    std_logic;
	in1348                               :   IN    std_logic;
	in1349                               :   IN    std_logic;
	in1350                               :   IN    std_logic;
	in1351                               :   IN    std_logic;
	in1352                               :   IN    std_logic;
	in1353                               :   IN    std_logic;
	in1354                               :   IN    std_logic;
	in1355                               :   IN    std_logic;
	in1356                               :   IN    std_logic;
	in1357                               :   IN    std_logic;
	in1358                               :   IN    std_logic;
	in1359                               :   IN    std_logic;
	in1360                               :   IN    std_logic;
	in1361                               :   IN    std_logic;
	in1362                               :   IN    std_logic;
	in1363                               :   IN    std_logic;
	in1364                               :   IN    std_logic;
	in1365                               :   IN    std_logic;
	in1366                               :   IN    std_logic;
	in1367                               :   IN    std_logic;
	in1368                               :   IN    std_logic;
	in1369                               :   IN    std_logic;
	in1370                               :   IN    std_logic;
	in1371                               :   IN    std_logic;
	in1372                               :   IN    std_logic;
	in1373                               :   IN    std_logic;
	in1374                               :   IN    std_logic;
	in1375                               :   IN    std_logic;
	in1376                               :   IN    std_logic;
	in1377                               :   IN    std_logic;
	in1378                               :   IN    std_logic;
	in1379                               :   IN    std_logic;
	in1380                               :   IN    std_logic;
	in1381                               :   IN    std_logic;
	in1382                               :   IN    std_logic;
	in1383                               :   IN    std_logic;
	in1384                               :   IN    std_logic;
	in1385                               :   IN    std_logic;
	in1386                               :   IN    std_logic;
	in1387                               :   IN    std_logic;
	in1388                               :   IN    std_logic;
	in1389                               :   IN    std_logic;
	in1390                               :   IN    std_logic;
	in1391                               :   IN    std_logic;
	in1392                               :   IN    std_logic;
	in1393                               :   IN    std_logic;
	in1394                               :   IN    std_logic;
	in1395                               :   IN    std_logic;
	in1396                               :   IN    std_logic;
	in1397                               :   IN    std_logic;
	in1398                               :   IN    std_logic;
	in1399                               :   IN    std_logic;
	in1400                               :   IN    std_logic;
	in1401                               :   IN    std_logic;
	in1402                               :   IN    std_logic;
	in1403                               :   IN    std_logic;
	in1404                               :   IN    std_logic;
	in1405                               :   IN    std_logic;
	in1406                               :   IN    std_logic;
	in1407                               :   IN    std_logic;
	in1408                               :   IN    std_logic;
	in1409                               :   IN    std_logic;
	in1410                               :   IN    std_logic;
	in1411                               :   IN    std_logic;
	in1412                               :   IN    std_logic;
	in1413                               :   IN    std_logic;
	in1414                               :   IN    std_logic;
	in1415                               :   IN    std_logic;
	in1416                               :   IN    std_logic;
	in1417                               :   IN    std_logic;
	in1418                               :   IN    std_logic;
	in1419                               :   IN    std_logic;
	in1420                               :   IN    std_logic;
	in1421                               :   IN    std_logic;
	in1422                               :   IN    std_logic;
	in1423                               :   IN    std_logic;
	in1424                               :   IN    std_logic;
	in1425                               :   IN    std_logic;
	in1426                               :   IN    std_logic;
	in1427                               :   IN    std_logic;
	in1428                               :   IN    std_logic;
	in1429                               :   IN    std_logic;
	in1430                               :   IN    std_logic;
	in1431                               :   IN    std_logic;
	in1432                               :   IN    std_logic;
	in1433                               :   IN    std_logic;
	in1434                               :   IN    std_logic;
	in1435                               :   IN    std_logic;
	in1436                               :   IN    std_logic;
	in1437                               :   IN    std_logic;
	in1438                               :   IN    std_logic;
	in1439                               :   IN    std_logic;
	in1440                               :   IN    std_logic;
	in1441                               :   IN    std_logic;
	in1442                               :   IN    std_logic;
	in1443                               :   IN    std_logic;
	in1444                               :   IN    std_logic;
	in1445                               :   IN    std_logic;
	in1446                               :   IN    std_logic;
	in1447                               :   IN    std_logic;
	in1448                               :   IN    std_logic;
	in1449                               :   IN    std_logic;
	in1450                               :   IN    std_logic;
	in1451                               :   IN    std_logic;
	in1452                               :   IN    std_logic;
	in1453                               :   IN    std_logic;
	in1454                               :   IN    std_logic;
	in1455                               :   IN    std_logic;
	in1456                               :   IN    std_logic;
	in1457                               :   IN    std_logic;
	in1458                               :   IN    std_logic;
	in1459                               :   IN    std_logic;
	in1460                               :   IN    std_logic;
	in1461                               :   IN    std_logic;
	in1462                               :   IN    std_logic;
	in1463                               :   IN    std_logic;
	in1464                               :   IN    std_logic;
	in1465                               :   IN    std_logic;
	in1466                               :   IN    std_logic;
	in1467                               :   IN    std_logic;
	in1468                               :   IN    std_logic;
	in1469                               :   IN    std_logic;
	in1470                               :   IN    std_logic;
	in1471                               :   IN    std_logic;
	in1472                               :   IN    std_logic;
	in1473                               :   IN    std_logic;
	in1474                               :   IN    std_logic;
	in1475                               :   IN    std_logic;
	in1476                               :   IN    std_logic;
	in1477                               :   IN    std_logic;
	in1478                               :   IN    std_logic;
	in1479                               :   IN    std_logic;
	in1480                               :   IN    std_logic;
	in1481                               :   IN    std_logic;
	in1482                               :   IN    std_logic;
	in1483                               :   IN    std_logic;
	in1484                               :   IN    std_logic;
	in1485                               :   IN    std_logic;
	in1486                               :   IN    std_logic;
	in1487                               :   IN    std_logic;
	in1488                               :   IN    std_logic;
	in1489                               :   IN    std_logic;
	in1490                               :   IN    std_logic;
	in1491                               :   IN    std_logic;
	in1492                               :   IN    std_logic;
	in1493                               :   IN    std_logic;
	in1494                               :   IN    std_logic;
	in1495                               :   IN    std_logic;
	in1496                               :   IN    std_logic;
	in1497                               :   IN    std_logic;
	in1498                               :   IN    std_logic;
	in1499                               :   IN    std_logic;
	in1500                               :   IN    std_logic;
	in1501                               :   IN    std_logic;
	in1502                               :   IN    std_logic;
	in1503                               :   IN    std_logic;
	in1504                               :   IN    std_logic;
	in1505                               :   IN    std_logic;
	in1506                               :   IN    std_logic;
	in1507                               :   IN    std_logic;
	in1508                               :   IN    std_logic;
	in1509                               :   IN    std_logic;
	in1510                               :   IN    std_logic;
	in1511                               :   IN    std_logic;
	in1512                               :   IN    std_logic;
	in1513                               :   IN    std_logic;
	in1514                               :   IN    std_logic;
	in1515                               :   IN    std_logic;
	in1516                               :   IN    std_logic;
	in1517                               :   IN    std_logic;
	in1518                               :   IN    std_logic;
	in1519                               :   IN    std_logic;
	in1520                               :   IN    std_logic;
	in1521                               :   IN    std_logic;
	in1522                               :   IN    std_logic;
	in1523                               :   IN    std_logic;
	in1524                               :   IN    std_logic;
	in1525                               :   IN    std_logic;
	in1526                               :   IN    std_logic;
	in1527                               :   IN    std_logic;
	in1528                               :   IN    std_logic;
	in1529                               :   IN    std_logic;
	in1530                               :   IN    std_logic;
	in1531                               :   IN    std_logic;
	in1532                               :   IN    std_logic;
	in1533                               :   IN    std_logic;
	in1534                               :   IN    std_logic;
	in1535                               :   IN    std_logic;
	in1536                               :   IN    std_logic;
	in1537                               :   IN    std_logic;
	in1538                               :   IN    std_logic;
	in1539                               :   IN    std_logic;
	in1540                               :   IN    std_logic;
	in1541                               :   IN    std_logic;
	in1542                               :   IN    std_logic;
	in1543                               :   IN    std_logic;
	in1544                               :   IN    std_logic;
	in1545                               :   IN    std_logic;
	in1546                               :   IN    std_logic;
	in1547                               :   IN    std_logic;
	in1548                               :   IN    std_logic;
	in1549                               :   IN    std_logic;
	in1550                               :   IN    std_logic;
	in1551                               :   IN    std_logic;
	in1552                               :   IN    std_logic;
	in1553                               :   IN    std_logic;
	in1554                               :   IN    std_logic;
	in1555                               :   IN    std_logic;
	in1556                               :   IN    std_logic;
	in1557                               :   IN    std_logic;
	in1558                               :   IN    std_logic;
	in1559                               :   IN    std_logic;
	in1560                               :   IN    std_logic;
	in1561                               :   IN    std_logic;
	in1562                               :   IN    std_logic;
	in1563                               :   IN    std_logic;
	in1564                               :   IN    std_logic;
	in1565                               :   IN    std_logic;
	in1566                               :   IN    std_logic;
	in1567                               :   IN    std_logic;
	in1568                               :   IN    std_logic;
	in1569                               :   IN    std_logic;
	in1570                               :   IN    std_logic;
	in1571                               :   IN    std_logic;
	in1572                               :   IN    std_logic;
	in1573                               :   IN    std_logic;
	in1574                               :   IN    std_logic;
	in1575                               :   IN    std_logic;
	in1576                               :   IN    std_logic;
	in1577                               :   IN    std_logic;
	in1578                               :   IN    std_logic;
	in1579                               :   IN    std_logic;
	in1580                               :   IN    std_logic;
	in1581                               :   IN    std_logic;
	in1582                               :   IN    std_logic;
	in1583                               :   IN    std_logic;
	in1584                               :   IN    std_logic;
	in1585                               :   IN    std_logic;
	in1586                               :   IN    std_logic;
	in1587                               :   IN    std_logic;
	in1588                               :   IN    std_logic;
	in1589                               :   IN    std_logic;
	in1590                               :   IN    std_logic;
	in1591                               :   IN    std_logic;
	in1592                               :   IN    std_logic;
	in1593                               :   IN    std_logic;
	in1594                               :   IN    std_logic;
	in1595                               :   IN    std_logic;
	in1596                               :   IN    std_logic;
	in1597                               :   IN    std_logic;
	in1598                               :   IN    std_logic;
	in1599                               :   IN    std_logic;
	in1600                               :   IN    std_logic;
	in1601                               :   IN    std_logic;
	in1602                               :   IN    std_logic;
	in1603                               :   IN    std_logic;
	in1604                               :   IN    std_logic;
	in1605                               :   IN    std_logic;
	in1606                               :   IN    std_logic;
	in1607                               :   IN    std_logic;
	in1608                               :   IN    std_logic;
	in1609                               :   IN    std_logic;
	in1610                               :   IN    std_logic;
	in1611                               :   IN    std_logic;
	in1612                               :   IN    std_logic;
	in1613                               :   IN    std_logic;
	in1614                               :   IN    std_logic;
	in1615                               :   IN    std_logic;
	in1616                               :   IN    std_logic;
	in1617                               :   IN    std_logic;
	in1618                               :   IN    std_logic;
	in1619                               :   IN    std_logic;
	in1620                               :   IN    std_logic;
	in1621                               :   IN    std_logic;
	in1622                               :   IN    std_logic;
	in1623                               :   IN    std_logic;
	in1624                               :   IN    std_logic;
	in1625                               :   IN    std_logic;
	in1626                               :   IN    std_logic;
	in1627                               :   IN    std_logic;
	in1628                               :   IN    std_logic;
	in1629                               :   IN    std_logic;
	in1630                               :   IN    std_logic;
	in1631                               :   IN    std_logic;
	in1632                               :   IN    std_logic;
	in1633                               :   IN    std_logic;
	in1634                               :   IN    std_logic;
	in1635                               :   IN    std_logic;
	in1636                               :   IN    std_logic;
	in1637                               :   IN    std_logic;
	in1638                               :   IN    std_logic;
	in1639                               :   IN    std_logic;
	in1640                               :   IN    std_logic;
	in1641                               :   IN    std_logic;
	in1642                               :   IN    std_logic;
	in1643                               :   IN    std_logic;
	in1644                               :   IN    std_logic;
	in1645                               :   IN    std_logic;
	in1646                               :   IN    std_logic;
	in1647                               :   IN    std_logic;
	in1648                               :   IN    std_logic;
	in1649                               :   IN    std_logic;
	in1650                               :   IN    std_logic;
	in1651                               :   IN    std_logic;
	in1652                               :   IN    std_logic;
	in1653                               :   IN    std_logic;
	in1654                               :   IN    std_logic;
	in1655                               :   IN    std_logic;
	in1656                               :   IN    std_logic;
	in1657                               :   IN    std_logic;
	in1658                               :   IN    std_logic;
	in1659                               :   IN    std_logic;
	in1660                               :   IN    std_logic;
	in1661                               :   IN    std_logic;
	in1662                               :   IN    std_logic;
	in1663                               :   IN    std_logic;
	in1664                               :   IN    std_logic;
	in1665                               :   IN    std_logic;
	in1666                               :   IN    std_logic;
	in1667                               :   IN    std_logic;
	in1668                               :   IN    std_logic;
	in1669                               :   IN    std_logic;
	in1670                               :   IN    std_logic;
	in1671                               :   IN    std_logic;
	in1672                               :   IN    std_logic;
	in1673                               :   IN    std_logic;
	in1674                               :   IN    std_logic;
	in1675                               :   IN    std_logic;
	in1676                               :   IN    std_logic;
	in1677                               :   IN    std_logic;
	in1678                               :   IN    std_logic;
	in1679                               :   IN    std_logic;
	in1680                               :   IN    std_logic;
	in1681                               :   IN    std_logic;
	in1682                               :   IN    std_logic;
	in1683                               :   IN    std_logic;
	in1684                               :   IN    std_logic;
	in1685                               :   IN    std_logic;
	in1686                               :   IN    std_logic;
	in1687                               :   IN    std_logic;
	in1688                               :   IN    std_logic;
	in1689                               :   IN    std_logic;
	in1690                               :   IN    std_logic;
	in1691                               :   IN    std_logic;
	in1692                               :   IN    std_logic;
	in1693                               :   IN    std_logic;
	in1694                               :   IN    std_logic;
	in1695                               :   IN    std_logic;
	in1696                               :   IN    std_logic;
	in1697                               :   IN    std_logic;
	in1698                               :   IN    std_logic;
	in1699                               :   IN    std_logic;
	in1700                               :   IN    std_logic;
	in1701                               :   IN    std_logic;
	in1702                               :   IN    std_logic;
	in1703                               :   IN    std_logic;
	in1704                               :   IN    std_logic;
	in1705                               :   IN    std_logic;
	in1706                               :   IN    std_logic;
	in1707                               :   IN    std_logic;
	in1708                               :   IN    std_logic;
	in1709                               :   IN    std_logic;
	in1710                               :   IN    std_logic;
	in1711                               :   IN    std_logic;
	in1712                               :   IN    std_logic;
	in1713                               :   IN    std_logic;
	in1714                               :   IN    std_logic;
	in1715                               :   IN    std_logic;
	in1716                               :   IN    std_logic;
	in1717                               :   IN    std_logic;
	in1718                               :   IN    std_logic;
	in1719                               :   IN    std_logic;
	in1720                               :   IN    std_logic;
	in1721                               :   IN    std_logic;
	in1722                               :   IN    std_logic;
	in1723                               :   IN    std_logic;
	in1724                               :   IN    std_logic;
	in1725                               :   IN    std_logic;
	in1726                               :   IN    std_logic;
	in1727                               :   IN    std_logic;
	in1728                               :   IN    std_logic;
	in1729                               :   IN    std_logic;
	in1730                               :   IN    std_logic;
	in1731                               :   IN    std_logic;
	in1732                               :   IN    std_logic;
	in1733                               :   IN    std_logic;
	in1734                               :   IN    std_logic;
	in1735                               :   IN    std_logic;
	in1736                               :   IN    std_logic;
	in1737                               :   IN    std_logic;
	in1738                               :   IN    std_logic;
	in1739                               :   IN    std_logic;
	in1740                               :   IN    std_logic;
	in1741                               :   IN    std_logic;
	in1742                               :   IN    std_logic;
	in1743                               :   IN    std_logic;
	in1744                               :   IN    std_logic;
	in1745                               :   IN    std_logic;
	in1746                               :   IN    std_logic;
	in1747                               :   IN    std_logic;
	in1748                               :   IN    std_logic;
	in1749                               :   IN    std_logic;
	in1750                               :   IN    std_logic;
	in1751                               :   IN    std_logic;
	in1752                               :   IN    std_logic;
	in1753                               :   IN    std_logic;
	in1754                               :   IN    std_logic;
	in1755                               :   IN    std_logic;
	in1756                               :   IN    std_logic;
	in1757                               :   IN    std_logic;
	in1758                               :   IN    std_logic;
	in1759                               :   IN    std_logic;
	in1760                               :   IN    std_logic;
	in1761                               :   IN    std_logic;
	in1762                               :   IN    std_logic;
	in1763                               :   IN    std_logic;
	in1764                               :   IN    std_logic;
	in1765                               :   IN    std_logic;
	in1766                               :   IN    std_logic;
	in1767                               :   IN    std_logic;
	in1768                               :   IN    std_logic;
	in1769                               :   IN    std_logic;
	in1770                               :   IN    std_logic;
	in1771                               :   IN    std_logic;
	in1772                               :   IN    std_logic;
	in1773                               :   IN    std_logic;
	in1774                               :   IN    std_logic;
	in1775                               :   IN    std_logic;
	in1776                               :   IN    std_logic;
	in1777                               :   IN    std_logic;
	in1778                               :   IN    std_logic;
	in1779                               :   IN    std_logic;
	in1780                               :   IN    std_logic;
	in1781                               :   IN    std_logic;
	in1782                               :   IN    std_logic;
	in1783                               :   IN    std_logic;
	in1784                               :   IN    std_logic;
	in1785                               :   IN    std_logic;
	in1786                               :   IN    std_logic;
	in1787                               :   IN    std_logic;
	in1788                               :   IN    std_logic;
	in1789                               :   IN    std_logic;
	in1790                               :   IN    std_logic;
	in1791                               :   IN    std_logic;
	in1792                               :   IN    std_logic;
	in1793                               :   IN    std_logic;
	in1794                               :   IN    std_logic;
	in1795                               :   IN    std_logic;
	in1796                               :   IN    std_logic;
	in1797                               :   IN    std_logic;
	in1798                               :   IN    std_logic;
	in1799                               :   IN    std_logic;
	in1800                               :   IN    std_logic;
	in1801                               :   IN    std_logic;
	in1802                               :   IN    std_logic;
	in1803                               :   IN    std_logic;
	in1804                               :   IN    std_logic;
	in1805                               :   IN    std_logic;
	in1806                               :   IN    std_logic;
	in1807                               :   IN    std_logic;
	in1808                               :   IN    std_logic;
	in1809                               :   IN    std_logic;
	in1810                               :   IN    std_logic;
	in1811                               :   IN    std_logic;
	in1812                               :   IN    std_logic;
	in1813                               :   IN    std_logic;
	in1814                               :   IN    std_logic;
	in1815                               :   IN    std_logic;
	in1816                               :   IN    std_logic;
	in1817                               :   IN    std_logic;
	in1818                               :   IN    std_logic;
	in1819                               :   IN    std_logic;
	in1820                               :   IN    std_logic;
	in1821                               :   IN    std_logic;
	in1822                               :   IN    std_logic;
	in1823                               :   IN    std_logic;
	in1824                               :   IN    std_logic;
	in1825                               :   IN    std_logic;
	in1826                               :   IN    std_logic;
	in1827                               :   IN    std_logic;
	in1828                               :   IN    std_logic;
	in1829                               :   IN    std_logic;
	in1830                               :   IN    std_logic;
	in1831                               :   IN    std_logic;
	in1832                               :   IN    std_logic;
	in1833                               :   IN    std_logic;
	in1834                               :   IN    std_logic;
	in1835                               :   IN    std_logic;
	in1836                               :   IN    std_logic;
	in1837                               :   IN    std_logic;
	in1838                               :   IN    std_logic;
	in1839                               :   IN    std_logic;
	in1840                               :   IN    std_logic;
	in1841                               :   IN    std_logic;
	in1842                               :   IN    std_logic;
	in1843                               :   IN    std_logic;
	in1844                               :   IN    std_logic;
	in1845                               :   IN    std_logic;
	in1846                               :   IN    std_logic;
	in1847                               :   IN    std_logic;
	in1848                               :   IN    std_logic;
	in1849                               :   IN    std_logic;
	in1850                               :   IN    std_logic;
	in1851                               :   IN    std_logic;
	in1852                               :   IN    std_logic;
	in1853                               :   IN    std_logic;
	in1854                               :   IN    std_logic;
	in1855                               :   IN    std_logic;
	in1856                               :   IN    std_logic;
	in1857                               :   IN    std_logic;
	in1858                               :   IN    std_logic;
	in1859                               :   IN    std_logic;
	in1860                               :   IN    std_logic;
	in1861                               :   IN    std_logic;
	in1862                               :   IN    std_logic;
	in1863                               :   IN    std_logic;
	in1864                               :   IN    std_logic;
	in1865                               :   IN    std_logic;
	in1866                               :   IN    std_logic;
	in1867                               :   IN    std_logic;
	in1868                               :   IN    std_logic;
	in1869                               :   IN    std_logic;
	in1870                               :   IN    std_logic;
	in1871                               :   IN    std_logic;
	in1872                               :   IN    std_logic;
	in1873                               :   IN    std_logic;
	in1874                               :   IN    std_logic;
	in1875                               :   IN    std_logic;
	in1876                               :   IN    std_logic;
	in1877                               :   IN    std_logic;
	in1878                               :   IN    std_logic;
	in1879                               :   IN    std_logic;
	in1880                               :   IN    std_logic;
	in1881                               :   IN    std_logic;
	in1882                               :   IN    std_logic;
	in1883                               :   IN    std_logic;
	in1884                               :   IN    std_logic;
	in1885                               :   IN    std_logic;
	in1886                               :   IN    std_logic;
	in1887                               :   IN    std_logic;
	in1888                               :   IN    std_logic;
	in1889                               :   IN    std_logic;
	in1890                               :   IN    std_logic;
	in1891                               :   IN    std_logic;
	in1892                               :   IN    std_logic;
	in1893                               :   IN    std_logic;
	in1894                               :   IN    std_logic;
	in1895                               :   IN    std_logic;
	in1896                               :   IN    std_logic;
	in1897                               :   IN    std_logic;
	in1898                               :   IN    std_logic;
	in1899                               :   IN    std_logic;
	in1900                               :   IN    std_logic;
	in1901                               :   IN    std_logic;
	in1902                               :   IN    std_logic;
	in1903                               :   IN    std_logic;
	in1904                               :   IN    std_logic;
	in1905                               :   IN    std_logic;
	in1906                               :   IN    std_logic;
	in1907                               :   IN    std_logic;
	in1908                               :   IN    std_logic;
	in1909                               :   IN    std_logic;
	in1910                               :   IN    std_logic;
	in1911                               :   IN    std_logic;
	in1912                               :   IN    std_logic;
	in1913                               :   IN    std_logic;
	in1914                               :   IN    std_logic;
	in1915                               :   IN    std_logic;
	in1916                               :   IN    std_logic;
	in1917                               :   IN    std_logic;
	in1918                               :   IN    std_logic;
	in1919                               :   IN    std_logic;
	in1920                               :   IN    std_logic;
	in1921                               :   IN    std_logic;
	in1922                               :   IN    std_logic;
	in1923                               :   IN    std_logic;
	in1924                               :   IN    std_logic;
	in1925                               :   IN    std_logic;
	in1926                               :   IN    std_logic;
	in1927                               :   IN    std_logic;
	in1928                               :   IN    std_logic;
	in1929                               :   IN    std_logic;
	in1930                               :   IN    std_logic;
	in1931                               :   IN    std_logic;
	in1932                               :   IN    std_logic;
	in1933                               :   IN    std_logic;
	in1934                               :   IN    std_logic;
	in1935                               :   IN    std_logic;
	in1936                               :   IN    std_logic;
	in1937                               :   IN    std_logic;
	in1938                               :   IN    std_logic;
	in1939                               :   IN    std_logic;
	in1940                               :   IN    std_logic;
	in1941                               :   IN    std_logic;
	in1942                               :   IN    std_logic;
	in1943                               :   IN    std_logic;
	in1944                               :   IN    std_logic;
	in1945                               :   IN    std_logic;
	in1946                               :   IN    std_logic;
	in1947                               :   IN    std_logic;
	in1948                               :   IN    std_logic;
	in1949                               :   IN    std_logic;
	in1950                               :   IN    std_logic;
	in1951                               :   IN    std_logic;
	in1952                               :   IN    std_logic;
	in1953                               :   IN    std_logic;
	in1954                               :   IN    std_logic;
	in1955                               :   IN    std_logic;
	in1956                               :   IN    std_logic;
	in1957                               :   IN    std_logic;
	in1958                               :   IN    std_logic;
	in1959                               :   IN    std_logic;
	in1960                               :   IN    std_logic;
	in1961                               :   IN    std_logic;
	in1962                               :   IN    std_logic;
	in1963                               :   IN    std_logic;
	in1964                               :   IN    std_logic;
	in1965                               :   IN    std_logic;
	in1966                               :   IN    std_logic;
	in1967                               :   IN    std_logic;
	in1968                               :   IN    std_logic;
	in1969                               :   IN    std_logic;
	in1970                               :   IN    std_logic;
	in1971                               :   IN    std_logic;
	in1972                               :   IN    std_logic;
	in1973                               :   IN    std_logic;
	in1974                               :   IN    std_logic;
	in1975                               :   IN    std_logic;
	in1976                               :   IN    std_logic;
	in1977                               :   IN    std_logic;
	in1978                               :   IN    std_logic;
	in1979                               :   IN    std_logic;
	in1980                               :   IN    std_logic;
	in1981                               :   IN    std_logic;
	in1982                               :   IN    std_logic;
	in1983                               :   IN    std_logic;
	in1984                               :   IN    std_logic;
	in1985                               :   IN    std_logic;
	in1986                               :   IN    std_logic;
	in1987                               :   IN    std_logic;
	in1988                               :   IN    std_logic;
	in1989                               :   IN    std_logic;
	in1990                               :   IN    std_logic;
	in1991                               :   IN    std_logic;
	in1992                               :   IN    std_logic;
	in1993                               :   IN    std_logic;
	in1994                               :   IN    std_logic;
	in1995                               :   IN    std_logic;
	in1996                               :   IN    std_logic;
	in1997                               :   IN    std_logic;
	in1998                               :   IN    std_logic;
	in1999                               :   IN    std_logic;
	in2000                               :   IN    std_logic;
	in2001                               :   IN    std_logic;
	in2002                               :   IN    std_logic;
	in2003                               :   IN    std_logic;
	in2004                               :   IN    std_logic;
	in2005                               :   IN    std_logic;
	in2006                               :   IN    std_logic;
	in2007                               :   IN    std_logic;
	in2008                               :   IN    std_logic;
	in2009                               :   IN    std_logic;
	in2010                               :   IN    std_logic;
	in2011                               :   IN    std_logic;
	in2012                               :   IN    std_logic;
	in2013                               :   IN    std_logic;
	in2014                               :   IN    std_logic;
	in2015                               :   IN    std_logic;
	in2016                               :   IN    std_logic;
	in2017                               :   IN    std_logic;
	in2018                               :   IN    std_logic;
	in2019                               :   IN    std_logic;
	in2020                               :   IN    std_logic;
	in2021                               :   IN    std_logic;
	in2022                               :   IN    std_logic;
	in2023                               :   IN    std_logic;
	in2024                               :   IN    std_logic;
	in2025                               :   IN    std_logic;
	in2026                               :   IN    std_logic;
	in2027                               :   IN    std_logic;
	in2028                               :   IN    std_logic;
	in2029                               :   IN    std_logic;
	in2030                               :   IN    std_logic;
	in2031                               :   IN    std_logic;
	in2032                               :   IN    std_logic;
	in2033                               :   IN    std_logic;
	in2034                               :   IN    std_logic;
	in2035                               :   IN    std_logic;
	in2036                               :   IN    std_logic;
	in2037                               :   IN    std_logic;
	in2038                               :   IN    std_logic;
	in2039                               :   IN    std_logic;
	in2040                               :   IN    std_logic;
	in2041                               :   IN    std_logic;
	in2042                               :   IN    std_logic;
	in2043                               :   IN    std_logic;
	in2044                               :   IN    std_logic;
	in2045                               :   IN    std_logic;
	in2046                               :   IN    std_logic;
	in2047                               :   IN    std_logic;
	in2048                               :   IN    std_logic;
	out1                               :   OUT    std_logic;
	out2                               :   OUT    std_logic;
	out3                               :   OUT    std_logic;
	out4                               :   OUT    std_logic;
	out5                               :   OUT    std_logic;
	out6                               :   OUT    std_logic;
	out7                               :   OUT    std_logic;
	out8                               :   OUT    std_logic;
	out9                               :   OUT    std_logic;
	out10                               :   OUT    std_logic;
	out11                               :   OUT    std_logic;
	out12                               :   OUT    std_logic;
	out13                               :   OUT    std_logic;
	out14                               :   OUT    std_logic;
	out15                               :   OUT    std_logic;
	out16                               :   OUT    std_logic;
	out17                               :   OUT    std_logic;
	out18                               :   OUT    std_logic;
	out19                               :   OUT    std_logic;
	out20                               :   OUT    std_logic;
	out21                               :   OUT    std_logic;
	out22                               :   OUT    std_logic;
	out23                               :   OUT    std_logic;
	out24                               :   OUT    std_logic;
	out25                               :   OUT    std_logic;
	out26                               :   OUT    std_logic;
	out27                               :   OUT    std_logic;
	out28                               :   OUT    std_logic;
	out29                               :   OUT    std_logic;
	out30                               :   OUT    std_logic;
	out31                               :   OUT    std_logic;
	out32                               :   OUT    std_logic;
	out33                               :   OUT    std_logic;
	out34                               :   OUT    std_logic;
	out35                               :   OUT    std_logic;
	out36                               :   OUT    std_logic;
	out37                               :   OUT    std_logic;
	out38                               :   OUT    std_logic;
	out39                               :   OUT    std_logic;
	out40                               :   OUT    std_logic;
	out41                               :   OUT    std_logic;
	out42                               :   OUT    std_logic;
	out43                               :   OUT    std_logic;
	out44                               :   OUT    std_logic;
	out45                               :   OUT    std_logic;
	out46                               :   OUT    std_logic;
	out47                               :   OUT    std_logic;
	out48                               :   OUT    std_logic;
	out49                               :   OUT    std_logic;
	out50                               :   OUT    std_logic;
	out51                               :   OUT    std_logic;
	out52                               :   OUT    std_logic;
	out53                               :   OUT    std_logic;
	out54                               :   OUT    std_logic;
	out55                               :   OUT    std_logic;
	out56                               :   OUT    std_logic;
	out57                               :   OUT    std_logic;
	out58                               :   OUT    std_logic;
	out59                               :   OUT    std_logic;
	out60                               :   OUT    std_logic;
	out61                               :   OUT    std_logic;
	out62                               :   OUT    std_logic;
	out63                               :   OUT    std_logic;
	out64                               :   OUT    std_logic;
	out65                               :   OUT    std_logic;
	out66                               :   OUT    std_logic;
	out67                               :   OUT    std_logic;
	out68                               :   OUT    std_logic;
	out69                               :   OUT    std_logic;
	out70                               :   OUT    std_logic;
	out71                               :   OUT    std_logic;
	out72                               :   OUT    std_logic;
	out73                               :   OUT    std_logic;
	out74                               :   OUT    std_logic;
	out75                               :   OUT    std_logic;
	out76                               :   OUT    std_logic;
	out77                               :   OUT    std_logic;
	out78                               :   OUT    std_logic;
	out79                               :   OUT    std_logic;
	out80                               :   OUT    std_logic;
	out81                               :   OUT    std_logic;
	out82                               :   OUT    std_logic;
	out83                               :   OUT    std_logic;
	out84                               :   OUT    std_logic;
	out85                               :   OUT    std_logic;
	out86                               :   OUT    std_logic;
	out87                               :   OUT    std_logic;
	out88                               :   OUT    std_logic;
	out89                               :   OUT    std_logic;
	out90                               :   OUT    std_logic;
	out91                               :   OUT    std_logic;
	out92                               :   OUT    std_logic;
	out93                               :   OUT    std_logic;
	out94                               :   OUT    std_logic;
	out95                               :   OUT    std_logic;
	out96                               :   OUT    std_logic;
	out97                               :   OUT    std_logic;
	out98                               :   OUT    std_logic;
	out99                               :   OUT    std_logic;
	out100                               :   OUT    std_logic;
	out101                               :   OUT    std_logic;
	out102                               :   OUT    std_logic;
	out103                               :   OUT    std_logic;
	out104                               :   OUT    std_logic;
	out105                               :   OUT    std_logic;
	out106                               :   OUT    std_logic;
	out107                               :   OUT    std_logic;
	out108                               :   OUT    std_logic;
	out109                               :   OUT    std_logic;
	out110                               :   OUT    std_logic;
	out111                               :   OUT    std_logic;
	out112                               :   OUT    std_logic;
	out113                               :   OUT    std_logic;
	out114                               :   OUT    std_logic;
	out115                               :   OUT    std_logic;
	out116                               :   OUT    std_logic;
	out117                               :   OUT    std_logic;
	out118                               :   OUT    std_logic;
	out119                               :   OUT    std_logic;
	out120                               :   OUT    std_logic;
	out121                               :   OUT    std_logic;
	out122                               :   OUT    std_logic;
	out123                               :   OUT    std_logic;
	out124                               :   OUT    std_logic;
	out125                               :   OUT    std_logic;
	out126                               :   OUT    std_logic;
	out127                               :   OUT    std_logic;
	out128                               :   OUT    std_logic;
	out129                               :   OUT    std_logic;
	out130                               :   OUT    std_logic;
	out131                               :   OUT    std_logic;
	out132                               :   OUT    std_logic;
	out133                               :   OUT    std_logic;
	out134                               :   OUT    std_logic;
	out135                               :   OUT    std_logic;
	out136                               :   OUT    std_logic;
	out137                               :   OUT    std_logic;
	out138                               :   OUT    std_logic;
	out139                               :   OUT    std_logic;
	out140                               :   OUT    std_logic;
	out141                               :   OUT    std_logic;
	out142                               :   OUT    std_logic;
	out143                               :   OUT    std_logic;
	out144                               :   OUT    std_logic;
	out145                               :   OUT    std_logic;
	out146                               :   OUT    std_logic;
	out147                               :   OUT    std_logic;
	out148                               :   OUT    std_logic;
	out149                               :   OUT    std_logic;
	out150                               :   OUT    std_logic;
	out151                               :   OUT    std_logic;
	out152                               :   OUT    std_logic;
	out153                               :   OUT    std_logic;
	out154                               :   OUT    std_logic;
	out155                               :   OUT    std_logic;
	out156                               :   OUT    std_logic;
	out157                               :   OUT    std_logic;
	out158                               :   OUT    std_logic;
	out159                               :   OUT    std_logic;
	out160                               :   OUT    std_logic;
	out161                               :   OUT    std_logic;
	out162                               :   OUT    std_logic;
	out163                               :   OUT    std_logic;
	out164                               :   OUT    std_logic;
	out165                               :   OUT    std_logic;
	out166                               :   OUT    std_logic;
	out167                               :   OUT    std_logic;
	out168                               :   OUT    std_logic;
	out169                               :   OUT    std_logic;
	out170                               :   OUT    std_logic;
	out171                               :   OUT    std_logic;
	out172                               :   OUT    std_logic;
	out173                               :   OUT    std_logic;
	out174                               :   OUT    std_logic;
	out175                               :   OUT    std_logic;
	out176                               :   OUT    std_logic;
	out177                               :   OUT    std_logic;
	out178                               :   OUT    std_logic;
	out179                               :   OUT    std_logic;
	out180                               :   OUT    std_logic;
	out181                               :   OUT    std_logic;
	out182                               :   OUT    std_logic;
	out183                               :   OUT    std_logic;
	out184                               :   OUT    std_logic;
	out185                               :   OUT    std_logic;
	out186                               :   OUT    std_logic;
	out187                               :   OUT    std_logic;
	out188                               :   OUT    std_logic;
	out189                               :   OUT    std_logic;
	out190                               :   OUT    std_logic;
	out191                               :   OUT    std_logic;
	out192                               :   OUT    std_logic;
	out193                               :   OUT    std_logic;
	out194                               :   OUT    std_logic;
	out195                               :   OUT    std_logic;
	out196                               :   OUT    std_logic;
	out197                               :   OUT    std_logic;
	out198                               :   OUT    std_logic;
	out199                               :   OUT    std_logic;
	out200                               :   OUT    std_logic;
	out201                               :   OUT    std_logic;
	out202                               :   OUT    std_logic;
	out203                               :   OUT    std_logic;
	out204                               :   OUT    std_logic;
	out205                               :   OUT    std_logic;
	out206                               :   OUT    std_logic;
	out207                               :   OUT    std_logic;
	out208                               :   OUT    std_logic;
	out209                               :   OUT    std_logic;
	out210                               :   OUT    std_logic;
	out211                               :   OUT    std_logic;
	out212                               :   OUT    std_logic;
	out213                               :   OUT    std_logic;
	out214                               :   OUT    std_logic;
	out215                               :   OUT    std_logic;
	out216                               :   OUT    std_logic;
	out217                               :   OUT    std_logic;
	out218                               :   OUT    std_logic;
	out219                               :   OUT    std_logic;
	out220                               :   OUT    std_logic;
	out221                               :   OUT    std_logic;
	out222                               :   OUT    std_logic;
	out223                               :   OUT    std_logic;
	out224                               :   OUT    std_logic;
	out225                               :   OUT    std_logic;
	out226                               :   OUT    std_logic;
	out227                               :   OUT    std_logic;
	out228                               :   OUT    std_logic;
	out229                               :   OUT    std_logic;
	out230                               :   OUT    std_logic;
	out231                               :   OUT    std_logic;
	out232                               :   OUT    std_logic;
	out233                               :   OUT    std_logic;
	out234                               :   OUT    std_logic;
	out235                               :   OUT    std_logic;
	out236                               :   OUT    std_logic;
	out237                               :   OUT    std_logic;
	out238                               :   OUT    std_logic;
	out239                               :   OUT    std_logic;
	out240                               :   OUT    std_logic;
	out241                               :   OUT    std_logic;
	out242                               :   OUT    std_logic;
	out243                               :   OUT    std_logic;
	out244                               :   OUT    std_logic;
	out245                               :   OUT    std_logic;
	out246                               :   OUT    std_logic;
	out247                               :   OUT    std_logic;
	out248                               :   OUT    std_logic;
	out249                               :   OUT    std_logic;
	out250                               :   OUT    std_logic;
	out251                               :   OUT    std_logic;
	out252                               :   OUT    std_logic;
	out253                               :   OUT    std_logic;
	out254                               :   OUT    std_logic;
	out255                               :   OUT    std_logic;
	out256                               :   OUT    std_logic;
	out257                               :   OUT    std_logic;
	out258                               :   OUT    std_logic;
	out259                               :   OUT    std_logic;
	out260                               :   OUT    std_logic;
	out261                               :   OUT    std_logic;
	out262                               :   OUT    std_logic;
	out263                               :   OUT    std_logic;
	out264                               :   OUT    std_logic;
	out265                               :   OUT    std_logic;
	out266                               :   OUT    std_logic;
	out267                               :   OUT    std_logic;
	out268                               :   OUT    std_logic;
	out269                               :   OUT    std_logic;
	out270                               :   OUT    std_logic;
	out271                               :   OUT    std_logic;
	out272                               :   OUT    std_logic;
	out273                               :   OUT    std_logic;
	out274                               :   OUT    std_logic;
	out275                               :   OUT    std_logic;
	out276                               :   OUT    std_logic;
	out277                               :   OUT    std_logic;
	out278                               :   OUT    std_logic;
	out279                               :   OUT    std_logic;
	out280                               :   OUT    std_logic;
	out281                               :   OUT    std_logic;
	out282                               :   OUT    std_logic;
	out283                               :   OUT    std_logic;
	out284                               :   OUT    std_logic;
	out285                               :   OUT    std_logic;
	out286                               :   OUT    std_logic;
	out287                               :   OUT    std_logic;
	out288                               :   OUT    std_logic;
	out289                               :   OUT    std_logic;
	out290                               :   OUT    std_logic;
	out291                               :   OUT    std_logic;
	out292                               :   OUT    std_logic;
	out293                               :   OUT    std_logic;
	out294                               :   OUT    std_logic;
	out295                               :   OUT    std_logic;
	out296                               :   OUT    std_logic;
	out297                               :   OUT    std_logic;
	out298                               :   OUT    std_logic;
	out299                               :   OUT    std_logic;
	out300                               :   OUT    std_logic;
	out301                               :   OUT    std_logic;
	out302                               :   OUT    std_logic;
	out303                               :   OUT    std_logic;
	out304                               :   OUT    std_logic;
	out305                               :   OUT    std_logic;
	out306                               :   OUT    std_logic;
	out307                               :   OUT    std_logic;
	out308                               :   OUT    std_logic;
	out309                               :   OUT    std_logic;
	out310                               :   OUT    std_logic;
	out311                               :   OUT    std_logic;
	out312                               :   OUT    std_logic;
	out313                               :   OUT    std_logic;
	out314                               :   OUT    std_logic;
	out315                               :   OUT    std_logic;
	out316                               :   OUT    std_logic;
	out317                               :   OUT    std_logic;
	out318                               :   OUT    std_logic;
	out319                               :   OUT    std_logic;
	out320                               :   OUT    std_logic;
	out321                               :   OUT    std_logic;
	out322                               :   OUT    std_logic;
	out323                               :   OUT    std_logic;
	out324                               :   OUT    std_logic;
	out325                               :   OUT    std_logic;
	out326                               :   OUT    std_logic;
	out327                               :   OUT    std_logic;
	out328                               :   OUT    std_logic;
	out329                               :   OUT    std_logic;
	out330                               :   OUT    std_logic;
	out331                               :   OUT    std_logic;
	out332                               :   OUT    std_logic;
	out333                               :   OUT    std_logic;
	out334                               :   OUT    std_logic;
	out335                               :   OUT    std_logic;
	out336                               :   OUT    std_logic;
	out337                               :   OUT    std_logic;
	out338                               :   OUT    std_logic;
	out339                               :   OUT    std_logic;
	out340                               :   OUT    std_logic;
	out341                               :   OUT    std_logic;
	out342                               :   OUT    std_logic;
	out343                               :   OUT    std_logic;
	out344                               :   OUT    std_logic;
	out345                               :   OUT    std_logic;
	out346                               :   OUT    std_logic;
	out347                               :   OUT    std_logic;
	out348                               :   OUT    std_logic;
	out349                               :   OUT    std_logic;
	out350                               :   OUT    std_logic;
	out351                               :   OUT    std_logic;
	out352                               :   OUT    std_logic;
	out353                               :   OUT    std_logic;
	out354                               :   OUT    std_logic;
	out355                               :   OUT    std_logic;
	out356                               :   OUT    std_logic;
	out357                               :   OUT    std_logic;
	out358                               :   OUT    std_logic;
	out359                               :   OUT    std_logic;
	out360                               :   OUT    std_logic;
	out361                               :   OUT    std_logic;
	out362                               :   OUT    std_logic;
	out363                               :   OUT    std_logic;
	out364                               :   OUT    std_logic;
	out365                               :   OUT    std_logic;
	out366                               :   OUT    std_logic;
	out367                               :   OUT    std_logic;
	out368                               :   OUT    std_logic;
	out369                               :   OUT    std_logic;
	out370                               :   OUT    std_logic;
	out371                               :   OUT    std_logic;
	out372                               :   OUT    std_logic;
	out373                               :   OUT    std_logic;
	out374                               :   OUT    std_logic;
	out375                               :   OUT    std_logic;
	out376                               :   OUT    std_logic;
	out377                               :   OUT    std_logic;
	out378                               :   OUT    std_logic;
	out379                               :   OUT    std_logic;
	out380                               :   OUT    std_logic;
	out381                               :   OUT    std_logic;
	out382                               :   OUT    std_logic;
	out383                               :   OUT    std_logic;
	out384                               :   OUT    std_logic;
	out385                               :   OUT    std_logic;
	out386                               :   OUT    std_logic;
	out387                               :   OUT    std_logic;
	out388                               :   OUT    std_logic;
	out389                               :   OUT    std_logic;
	out390                               :   OUT    std_logic;
	out391                               :   OUT    std_logic;
	out392                               :   OUT    std_logic;
	out393                               :   OUT    std_logic;
	out394                               :   OUT    std_logic;
	out395                               :   OUT    std_logic;
	out396                               :   OUT    std_logic;
	out397                               :   OUT    std_logic;
	out398                               :   OUT    std_logic;
	out399                               :   OUT    std_logic;
	out400                               :   OUT    std_logic;
	out401                               :   OUT    std_logic;
	out402                               :   OUT    std_logic;
	out403                               :   OUT    std_logic;
	out404                               :   OUT    std_logic;
	out405                               :   OUT    std_logic;
	out406                               :   OUT    std_logic;
	out407                               :   OUT    std_logic;
	out408                               :   OUT    std_logic;
	out409                               :   OUT    std_logic;
	out410                               :   OUT    std_logic;
	out411                               :   OUT    std_logic;
	out412                               :   OUT    std_logic;
	out413                               :   OUT    std_logic;
	out414                               :   OUT    std_logic;
	out415                               :   OUT    std_logic;
	out416                               :   OUT    std_logic;
	out417                               :   OUT    std_logic;
	out418                               :   OUT    std_logic;
	out419                               :   OUT    std_logic;
	out420                               :   OUT    std_logic;
	out421                               :   OUT    std_logic;
	out422                               :   OUT    std_logic;
	out423                               :   OUT    std_logic;
	out424                               :   OUT    std_logic;
	out425                               :   OUT    std_logic;
	out426                               :   OUT    std_logic;
	out427                               :   OUT    std_logic;
	out428                               :   OUT    std_logic;
	out429                               :   OUT    std_logic;
	out430                               :   OUT    std_logic;
	out431                               :   OUT    std_logic;
	out432                               :   OUT    std_logic;
	out433                               :   OUT    std_logic;
	out434                               :   OUT    std_logic;
	out435                               :   OUT    std_logic;
	out436                               :   OUT    std_logic;
	out437                               :   OUT    std_logic;
	out438                               :   OUT    std_logic;
	out439                               :   OUT    std_logic;
	out440                               :   OUT    std_logic;
	out441                               :   OUT    std_logic;
	out442                               :   OUT    std_logic;
	out443                               :   OUT    std_logic;
	out444                               :   OUT    std_logic;
	out445                               :   OUT    std_logic;
	out446                               :   OUT    std_logic;
	out447                               :   OUT    std_logic;
	out448                               :   OUT    std_logic;
	out449                               :   OUT    std_logic;
	out450                               :   OUT    std_logic;
	out451                               :   OUT    std_logic;
	out452                               :   OUT    std_logic;
	out453                               :   OUT    std_logic;
	out454                               :   OUT    std_logic;
	out455                               :   OUT    std_logic;
	out456                               :   OUT    std_logic;
	out457                               :   OUT    std_logic;
	out458                               :   OUT    std_logic;
	out459                               :   OUT    std_logic;
	out460                               :   OUT    std_logic;
	out461                               :   OUT    std_logic;
	out462                               :   OUT    std_logic;
	out463                               :   OUT    std_logic;
	out464                               :   OUT    std_logic;
	out465                               :   OUT    std_logic;
	out466                               :   OUT    std_logic;
	out467                               :   OUT    std_logic;
	out468                               :   OUT    std_logic;
	out469                               :   OUT    std_logic;
	out470                               :   OUT    std_logic;
	out471                               :   OUT    std_logic;
	out472                               :   OUT    std_logic;
	out473                               :   OUT    std_logic;
	out474                               :   OUT    std_logic;
	out475                               :   OUT    std_logic;
	out476                               :   OUT    std_logic;
	out477                               :   OUT    std_logic;
	out478                               :   OUT    std_logic;
	out479                               :   OUT    std_logic;
	out480                               :   OUT    std_logic;
	out481                               :   OUT    std_logic;
	out482                               :   OUT    std_logic;
	out483                               :   OUT    std_logic;
	out484                               :   OUT    std_logic;
	out485                               :   OUT    std_logic;
	out486                               :   OUT    std_logic;
	out487                               :   OUT    std_logic;
	out488                               :   OUT    std_logic;
	out489                               :   OUT    std_logic;
	out490                               :   OUT    std_logic;
	out491                               :   OUT    std_logic;
	out492                               :   OUT    std_logic;
	out493                               :   OUT    std_logic;
	out494                               :   OUT    std_logic;
	out495                               :   OUT    std_logic;
	out496                               :   OUT    std_logic;
	out497                               :   OUT    std_logic;
	out498                               :   OUT    std_logic;
	out499                               :   OUT    std_logic;
	out500                               :   OUT    std_logic;
	out501                               :   OUT    std_logic;
	out502                               :   OUT    std_logic;
	out503                               :   OUT    std_logic;
	out504                               :   OUT    std_logic;
	out505                               :   OUT    std_logic;
	out506                               :   OUT    std_logic;
	out507                               :   OUT    std_logic;
	out508                               :   OUT    std_logic;
	out509                               :   OUT    std_logic;
	out510                               :   OUT    std_logic;
	out511                               :   OUT    std_logic;
	out512                               :   OUT    std_logic;
	out513                               :   OUT    std_logic;
	out514                               :   OUT    std_logic;
	out515                               :   OUT    std_logic;
	out516                               :   OUT    std_logic;
	out517                               :   OUT    std_logic;
	out518                               :   OUT    std_logic;
	out519                               :   OUT    std_logic;
	out520                               :   OUT    std_logic;
	out521                               :   OUT    std_logic;
	out522                               :   OUT    std_logic;
	out523                               :   OUT    std_logic;
	out524                               :   OUT    std_logic;
	out525                               :   OUT    std_logic;
	out526                               :   OUT    std_logic;
	out527                               :   OUT    std_logic;
	out528                               :   OUT    std_logic;
	out529                               :   OUT    std_logic;
	out530                               :   OUT    std_logic;
	out531                               :   OUT    std_logic;
	out532                               :   OUT    std_logic;
	out533                               :   OUT    std_logic;
	out534                               :   OUT    std_logic;
	out535                               :   OUT    std_logic;
	out536                               :   OUT    std_logic;
	out537                               :   OUT    std_logic;
	out538                               :   OUT    std_logic;
	out539                               :   OUT    std_logic;
	out540                               :   OUT    std_logic;
	out541                               :   OUT    std_logic;
	out542                               :   OUT    std_logic;
	out543                               :   OUT    std_logic;
	out544                               :   OUT    std_logic;
	out545                               :   OUT    std_logic;
	out546                               :   OUT    std_logic;
	out547                               :   OUT    std_logic;
	out548                               :   OUT    std_logic;
	out549                               :   OUT    std_logic;
	out550                               :   OUT    std_logic;
	out551                               :   OUT    std_logic;
	out552                               :   OUT    std_logic;
	out553                               :   OUT    std_logic;
	out554                               :   OUT    std_logic;
	out555                               :   OUT    std_logic;
	out556                               :   OUT    std_logic;
	out557                               :   OUT    std_logic;
	out558                               :   OUT    std_logic;
	out559                               :   OUT    std_logic;
	out560                               :   OUT    std_logic;
	out561                               :   OUT    std_logic;
	out562                               :   OUT    std_logic;
	out563                               :   OUT    std_logic;
	out564                               :   OUT    std_logic;
	out565                               :   OUT    std_logic;
	out566                               :   OUT    std_logic;
	out567                               :   OUT    std_logic;
	out568                               :   OUT    std_logic;
	out569                               :   OUT    std_logic;
	out570                               :   OUT    std_logic;
	out571                               :   OUT    std_logic;
	out572                               :   OUT    std_logic;
	out573                               :   OUT    std_logic;
	out574                               :   OUT    std_logic;
	out575                               :   OUT    std_logic;
	out576                               :   OUT    std_logic;
	out577                               :   OUT    std_logic;
	out578                               :   OUT    std_logic;
	out579                               :   OUT    std_logic;
	out580                               :   OUT    std_logic;
	out581                               :   OUT    std_logic;
	out582                               :   OUT    std_logic;
	out583                               :   OUT    std_logic;
	out584                               :   OUT    std_logic;
	out585                               :   OUT    std_logic;
	out586                               :   OUT    std_logic;
	out587                               :   OUT    std_logic;
	out588                               :   OUT    std_logic;
	out589                               :   OUT    std_logic;
	out590                               :   OUT    std_logic;
	out591                               :   OUT    std_logic;
	out592                               :   OUT    std_logic;
	out593                               :   OUT    std_logic;
	out594                               :   OUT    std_logic;
	out595                               :   OUT    std_logic;
	out596                               :   OUT    std_logic;
	out597                               :   OUT    std_logic;
	out598                               :   OUT    std_logic;
	out599                               :   OUT    std_logic;
	out600                               :   OUT    std_logic;
	out601                               :   OUT    std_logic;
	out602                               :   OUT    std_logic;
	out603                               :   OUT    std_logic;
	out604                               :   OUT    std_logic;
	out605                               :   OUT    std_logic;
	out606                               :   OUT    std_logic;
	out607                               :   OUT    std_logic;
	out608                               :   OUT    std_logic;
	out609                               :   OUT    std_logic;
	out610                               :   OUT    std_logic;
	out611                               :   OUT    std_logic;
	out612                               :   OUT    std_logic;
	out613                               :   OUT    std_logic;
	out614                               :   OUT    std_logic;
	out615                               :   OUT    std_logic;
	out616                               :   OUT    std_logic;
	out617                               :   OUT    std_logic;
	out618                               :   OUT    std_logic;
	out619                               :   OUT    std_logic;
	out620                               :   OUT    std_logic;
	out621                               :   OUT    std_logic;
	out622                               :   OUT    std_logic;
	out623                               :   OUT    std_logic;
	out624                               :   OUT    std_logic;
	out625                               :   OUT    std_logic;
	out626                               :   OUT    std_logic;
	out627                               :   OUT    std_logic;
	out628                               :   OUT    std_logic;
	out629                               :   OUT    std_logic;
	out630                               :   OUT    std_logic;
	out631                               :   OUT    std_logic;
	out632                               :   OUT    std_logic;
	out633                               :   OUT    std_logic;
	out634                               :   OUT    std_logic;
	out635                               :   OUT    std_logic;
	out636                               :   OUT    std_logic;
	out637                               :   OUT    std_logic;
	out638                               :   OUT    std_logic;
	out639                               :   OUT    std_logic;
	out640                               :   OUT    std_logic;
	out641                               :   OUT    std_logic;
	out642                               :   OUT    std_logic;
	out643                               :   OUT    std_logic;
	out644                               :   OUT    std_logic;
	out645                               :   OUT    std_logic;
	out646                               :   OUT    std_logic;
	out647                               :   OUT    std_logic;
	out648                               :   OUT    std_logic;
	out649                               :   OUT    std_logic;
	out650                               :   OUT    std_logic;
	out651                               :   OUT    std_logic;
	out652                               :   OUT    std_logic;
	out653                               :   OUT    std_logic;
	out654                               :   OUT    std_logic;
	out655                               :   OUT    std_logic;
	out656                               :   OUT    std_logic;
	out657                               :   OUT    std_logic;
	out658                               :   OUT    std_logic;
	out659                               :   OUT    std_logic;
	out660                               :   OUT    std_logic;
	out661                               :   OUT    std_logic;
	out662                               :   OUT    std_logic;
	out663                               :   OUT    std_logic;
	out664                               :   OUT    std_logic;
	out665                               :   OUT    std_logic;
	out666                               :   OUT    std_logic;
	out667                               :   OUT    std_logic;
	out668                               :   OUT    std_logic;
	out669                               :   OUT    std_logic;
	out670                               :   OUT    std_logic;
	out671                               :   OUT    std_logic;
	out672                               :   OUT    std_logic;
	out673                               :   OUT    std_logic;
	out674                               :   OUT    std_logic;
	out675                               :   OUT    std_logic;
	out676                               :   OUT    std_logic;
	out677                               :   OUT    std_logic;
	out678                               :   OUT    std_logic;
	out679                               :   OUT    std_logic;
	out680                               :   OUT    std_logic;
	out681                               :   OUT    std_logic;
	out682                               :   OUT    std_logic;
	out683                               :   OUT    std_logic;
	out684                               :   OUT    std_logic;
	out685                               :   OUT    std_logic;
	out686                               :   OUT    std_logic;
	out687                               :   OUT    std_logic;
	out688                               :   OUT    std_logic;
	out689                               :   OUT    std_logic;
	out690                               :   OUT    std_logic;
	out691                               :   OUT    std_logic;
	out692                               :   OUT    std_logic;
	out693                               :   OUT    std_logic;
	out694                               :   OUT    std_logic;
	out695                               :   OUT    std_logic;
	out696                               :   OUT    std_logic;
	out697                               :   OUT    std_logic;
	out698                               :   OUT    std_logic;
	out699                               :   OUT    std_logic;
	out700                               :   OUT    std_logic;
	out701                               :   OUT    std_logic;
	out702                               :   OUT    std_logic;
	out703                               :   OUT    std_logic;
	out704                               :   OUT    std_logic;
	out705                               :   OUT    std_logic;
	out706                               :   OUT    std_logic;
	out707                               :   OUT    std_logic;
	out708                               :   OUT    std_logic;
	out709                               :   OUT    std_logic;
	out710                               :   OUT    std_logic;
	out711                               :   OUT    std_logic;
	out712                               :   OUT    std_logic;
	out713                               :   OUT    std_logic;
	out714                               :   OUT    std_logic;
	out715                               :   OUT    std_logic;
	out716                               :   OUT    std_logic;
	out717                               :   OUT    std_logic;
	out718                               :   OUT    std_logic;
	out719                               :   OUT    std_logic;
	out720                               :   OUT    std_logic;
	out721                               :   OUT    std_logic;
	out722                               :   OUT    std_logic;
	out723                               :   OUT    std_logic;
	out724                               :   OUT    std_logic;
	out725                               :   OUT    std_logic;
	out726                               :   OUT    std_logic;
	out727                               :   OUT    std_logic;
	out728                               :   OUT    std_logic;
	out729                               :   OUT    std_logic;
	out730                               :   OUT    std_logic;
	out731                               :   OUT    std_logic;
	out732                               :   OUT    std_logic;
	out733                               :   OUT    std_logic;
	out734                               :   OUT    std_logic;
	out735                               :   OUT    std_logic;
	out736                               :   OUT    std_logic;
	out737                               :   OUT    std_logic;
	out738                               :   OUT    std_logic;
	out739                               :   OUT    std_logic;
	out740                               :   OUT    std_logic;
	out741                               :   OUT    std_logic;
	out742                               :   OUT    std_logic;
	out743                               :   OUT    std_logic;
	out744                               :   OUT    std_logic;
	out745                               :   OUT    std_logic;
	out746                               :   OUT    std_logic;
	out747                               :   OUT    std_logic;
	out748                               :   OUT    std_logic;
	out749                               :   OUT    std_logic;
	out750                               :   OUT    std_logic;
	out751                               :   OUT    std_logic;
	out752                               :   OUT    std_logic;
	out753                               :   OUT    std_logic;
	out754                               :   OUT    std_logic;
	out755                               :   OUT    std_logic;
	out756                               :   OUT    std_logic;
	out757                               :   OUT    std_logic;
	out758                               :   OUT    std_logic;
	out759                               :   OUT    std_logic;
	out760                               :   OUT    std_logic;
	out761                               :   OUT    std_logic;
	out762                               :   OUT    std_logic;
	out763                               :   OUT    std_logic;
	out764                               :   OUT    std_logic;
	out765                               :   OUT    std_logic;
	out766                               :   OUT    std_logic;
	out767                               :   OUT    std_logic;
	out768                               :   OUT    std_logic;
	out769                               :   OUT    std_logic;
	out770                               :   OUT    std_logic;
	out771                               :   OUT    std_logic;
	out772                               :   OUT    std_logic;
	out773                               :   OUT    std_logic;
	out774                               :   OUT    std_logic;
	out775                               :   OUT    std_logic;
	out776                               :   OUT    std_logic;
	out777                               :   OUT    std_logic;
	out778                               :   OUT    std_logic;
	out779                               :   OUT    std_logic;
	out780                               :   OUT    std_logic;
	out781                               :   OUT    std_logic;
	out782                               :   OUT    std_logic;
	out783                               :   OUT    std_logic;
	out784                               :   OUT    std_logic;
	out785                               :   OUT    std_logic;
	out786                               :   OUT    std_logic;
	out787                               :   OUT    std_logic;
	out788                               :   OUT    std_logic;
	out789                               :   OUT    std_logic;
	out790                               :   OUT    std_logic;
	out791                               :   OUT    std_logic;
	out792                               :   OUT    std_logic;
	out793                               :   OUT    std_logic;
	out794                               :   OUT    std_logic;
	out795                               :   OUT    std_logic;
	out796                               :   OUT    std_logic;
	out797                               :   OUT    std_logic;
	out798                               :   OUT    std_logic;
	out799                               :   OUT    std_logic;
	out800                               :   OUT    std_logic;
	out801                               :   OUT    std_logic;
	out802                               :   OUT    std_logic;
	out803                               :   OUT    std_logic;
	out804                               :   OUT    std_logic;
	out805                               :   OUT    std_logic;
	out806                               :   OUT    std_logic;
	out807                               :   OUT    std_logic;
	out808                               :   OUT    std_logic;
	out809                               :   OUT    std_logic;
	out810                               :   OUT    std_logic;
	out811                               :   OUT    std_logic;
	out812                               :   OUT    std_logic;
	out813                               :   OUT    std_logic;
	out814                               :   OUT    std_logic;
	out815                               :   OUT    std_logic;
	out816                               :   OUT    std_logic;
	out817                               :   OUT    std_logic;
	out818                               :   OUT    std_logic;
	out819                               :   OUT    std_logic;
	out820                               :   OUT    std_logic;
	out821                               :   OUT    std_logic;
	out822                               :   OUT    std_logic;
	out823                               :   OUT    std_logic;
	out824                               :   OUT    std_logic;
	out825                               :   OUT    std_logic;
	out826                               :   OUT    std_logic;
	out827                               :   OUT    std_logic;
	out828                               :   OUT    std_logic;
	out829                               :   OUT    std_logic;
	out830                               :   OUT    std_logic;
	out831                               :   OUT    std_logic;
	out832                               :   OUT    std_logic;
	out833                               :   OUT    std_logic;
	out834                               :   OUT    std_logic;
	out835                               :   OUT    std_logic;
	out836                               :   OUT    std_logic;
	out837                               :   OUT    std_logic;
	out838                               :   OUT    std_logic;
	out839                               :   OUT    std_logic;
	out840                               :   OUT    std_logic;
	out841                               :   OUT    std_logic;
	out842                               :   OUT    std_logic;
	out843                               :   OUT    std_logic;
	out844                               :   OUT    std_logic;
	out845                               :   OUT    std_logic;
	out846                               :   OUT    std_logic;
	out847                               :   OUT    std_logic;
	out848                               :   OUT    std_logic;
	out849                               :   OUT    std_logic;
	out850                               :   OUT    std_logic;
	out851                               :   OUT    std_logic;
	out852                               :   OUT    std_logic;
	out853                               :   OUT    std_logic;
	out854                               :   OUT    std_logic;
	out855                               :   OUT    std_logic;
	out856                               :   OUT    std_logic;
	out857                               :   OUT    std_logic;
	out858                               :   OUT    std_logic;
	out859                               :   OUT    std_logic;
	out860                               :   OUT    std_logic;
	out861                               :   OUT    std_logic;
	out862                               :   OUT    std_logic;
	out863                               :   OUT    std_logic;
	out864                               :   OUT    std_logic;
	out865                               :   OUT    std_logic;
	out866                               :   OUT    std_logic;
	out867                               :   OUT    std_logic;
	out868                               :   OUT    std_logic;
	out869                               :   OUT    std_logic;
	out870                               :   OUT    std_logic;
	out871                               :   OUT    std_logic;
	out872                               :   OUT    std_logic;
	out873                               :   OUT    std_logic;
	out874                               :   OUT    std_logic;
	out875                               :   OUT    std_logic;
	out876                               :   OUT    std_logic;
	out877                               :   OUT    std_logic;
	out878                               :   OUT    std_logic;
	out879                               :   OUT    std_logic;
	out880                               :   OUT    std_logic;
	out881                               :   OUT    std_logic;
	out882                               :   OUT    std_logic;
	out883                               :   OUT    std_logic;
	out884                               :   OUT    std_logic;
	out885                               :   OUT    std_logic;
	out886                               :   OUT    std_logic;
	out887                               :   OUT    std_logic;
	out888                               :   OUT    std_logic;
	out889                               :   OUT    std_logic;
	out890                               :   OUT    std_logic;
	out891                               :   OUT    std_logic;
	out892                               :   OUT    std_logic;
	out893                               :   OUT    std_logic;
	out894                               :   OUT    std_logic;
	out895                               :   OUT    std_logic;
	out896                               :   OUT    std_logic;
	out897                               :   OUT    std_logic;
	out898                               :   OUT    std_logic;
	out899                               :   OUT    std_logic;
	out900                               :   OUT    std_logic;
	out901                               :   OUT    std_logic;
	out902                               :   OUT    std_logic;
	out903                               :   OUT    std_logic;
	out904                               :   OUT    std_logic;
	out905                               :   OUT    std_logic;
	out906                               :   OUT    std_logic;
	out907                               :   OUT    std_logic;
	out908                               :   OUT    std_logic;
	out909                               :   OUT    std_logic;
	out910                               :   OUT    std_logic;
	out911                               :   OUT    std_logic;
	out912                               :   OUT    std_logic;
	out913                               :   OUT    std_logic;
	out914                               :   OUT    std_logic;
	out915                               :   OUT    std_logic;
	out916                               :   OUT    std_logic;
	out917                               :   OUT    std_logic;
	out918                               :   OUT    std_logic;
	out919                               :   OUT    std_logic;
	out920                               :   OUT    std_logic;
	out921                               :   OUT    std_logic;
	out922                               :   OUT    std_logic;
	out923                               :   OUT    std_logic;
	out924                               :   OUT    std_logic;
	out925                               :   OUT    std_logic;
	out926                               :   OUT    std_logic;
	out927                               :   OUT    std_logic;
	out928                               :   OUT    std_logic;
	out929                               :   OUT    std_logic;
	out930                               :   OUT    std_logic;
	out931                               :   OUT    std_logic;
	out932                               :   OUT    std_logic;
	out933                               :   OUT    std_logic;
	out934                               :   OUT    std_logic;
	out935                               :   OUT    std_logic;
	out936                               :   OUT    std_logic;
	out937                               :   OUT    std_logic;
	out938                               :   OUT    std_logic;
	out939                               :   OUT    std_logic;
	out940                               :   OUT    std_logic;
	out941                               :   OUT    std_logic;
	out942                               :   OUT    std_logic;
	out943                               :   OUT    std_logic;
	out944                               :   OUT    std_logic;
	out945                               :   OUT    std_logic;
	out946                               :   OUT    std_logic;
	out947                               :   OUT    std_logic;
	out948                               :   OUT    std_logic;
	out949                               :   OUT    std_logic;
	out950                               :   OUT    std_logic;
	out951                               :   OUT    std_logic;
	out952                               :   OUT    std_logic;
	out953                               :   OUT    std_logic;
	out954                               :   OUT    std_logic;
	out955                               :   OUT    std_logic;
	out956                               :   OUT    std_logic;
	out957                               :   OUT    std_logic;
	out958                               :   OUT    std_logic;
	out959                               :   OUT    std_logic;
	out960                               :   OUT    std_logic;
	out961                               :   OUT    std_logic;
	out962                               :   OUT    std_logic;
	out963                               :   OUT    std_logic;
	out964                               :   OUT    std_logic;
	out965                               :   OUT    std_logic;
	out966                               :   OUT    std_logic;
	out967                               :   OUT    std_logic;
	out968                               :   OUT    std_logic;
	out969                               :   OUT    std_logic;
	out970                               :   OUT    std_logic;
	out971                               :   OUT    std_logic;
	out972                               :   OUT    std_logic;
	out973                               :   OUT    std_logic;
	out974                               :   OUT    std_logic;
	out975                               :   OUT    std_logic;
	out976                               :   OUT    std_logic;
	out977                               :   OUT    std_logic;
	out978                               :   OUT    std_logic;
	out979                               :   OUT    std_logic;
	out980                               :   OUT    std_logic;
	out981                               :   OUT    std_logic;
	out982                               :   OUT    std_logic;
	out983                               :   OUT    std_logic;
	out984                               :   OUT    std_logic;
	out985                               :   OUT    std_logic;
	out986                               :   OUT    std_logic;
	out987                               :   OUT    std_logic;
	out988                               :   OUT    std_logic;
	out989                               :   OUT    std_logic;
	out990                               :   OUT    std_logic;
	out991                               :   OUT    std_logic;
	out992                               :   OUT    std_logic;
	out993                               :   OUT    std_logic;
	out994                               :   OUT    std_logic;
	out995                               :   OUT    std_logic;
	out996                               :   OUT    std_logic;
	out997                               :   OUT    std_logic;
	out998                               :   OUT    std_logic;
	out999                               :   OUT    std_logic;
	out1000                               :   OUT    std_logic;
	out1001                               :   OUT    std_logic;
	out1002                               :   OUT    std_logic;
	out1003                               :   OUT    std_logic;
	out1004                               :   OUT    std_logic;
	out1005                               :   OUT    std_logic;
	out1006                               :   OUT    std_logic;
	out1007                               :   OUT    std_logic;
	out1008                               :   OUT    std_logic;
	out1009                               :   OUT    std_logic;
	out1010                               :   OUT    std_logic;
	out1011                               :   OUT    std_logic;
	out1012                               :   OUT    std_logic;
	out1013                               :   OUT    std_logic;
	out1014                               :   OUT    std_logic;
	out1015                               :   OUT    std_logic;
	out1016                               :   OUT    std_logic;
	out1017                               :   OUT    std_logic;
	out1018                               :   OUT    std_logic;
	out1019                               :   OUT    std_logic;
	out1020                               :   OUT    std_logic;
	out1021                               :   OUT    std_logic;
	out1022                               :   OUT    std_logic;
	out1023                               :   OUT    std_logic;
	out1024                               :   OUT    std_logic;
	out1025                               :   OUT    std_logic;
	out1026                               :   OUT    std_logic;
	out1027                               :   OUT    std_logic;
	out1028                               :   OUT    std_logic;
	out1029                               :   OUT    std_logic;
	out1030                               :   OUT    std_logic;
	out1031                               :   OUT    std_logic;
	out1032                               :   OUT    std_logic;
	out1033                               :   OUT    std_logic;
	out1034                               :   OUT    std_logic;
	out1035                               :   OUT    std_logic;
	out1036                               :   OUT    std_logic;
	out1037                               :   OUT    std_logic;
	out1038                               :   OUT    std_logic;
	out1039                               :   OUT    std_logic;
	out1040                               :   OUT    std_logic;
	out1041                               :   OUT    std_logic;
	out1042                               :   OUT    std_logic;
	out1043                               :   OUT    std_logic;
	out1044                               :   OUT    std_logic;
	out1045                               :   OUT    std_logic;
	out1046                               :   OUT    std_logic;
	out1047                               :   OUT    std_logic;
	out1048                               :   OUT    std_logic;
	out1049                               :   OUT    std_logic;
	out1050                               :   OUT    std_logic;
	out1051                               :   OUT    std_logic;
	out1052                               :   OUT    std_logic;
	out1053                               :   OUT    std_logic;
	out1054                               :   OUT    std_logic;
	out1055                               :   OUT    std_logic;
	out1056                               :   OUT    std_logic;
	out1057                               :   OUT    std_logic;
	out1058                               :   OUT    std_logic;
	out1059                               :   OUT    std_logic;
	out1060                               :   OUT    std_logic;
	out1061                               :   OUT    std_logic;
	out1062                               :   OUT    std_logic;
	out1063                               :   OUT    std_logic;
	out1064                               :   OUT    std_logic;
	out1065                               :   OUT    std_logic;
	out1066                               :   OUT    std_logic;
	out1067                               :   OUT    std_logic;
	out1068                               :   OUT    std_logic;
	out1069                               :   OUT    std_logic;
	out1070                               :   OUT    std_logic;
	out1071                               :   OUT    std_logic;
	out1072                               :   OUT    std_logic;
	out1073                               :   OUT    std_logic;
	out1074                               :   OUT    std_logic;
	out1075                               :   OUT    std_logic;
	out1076                               :   OUT    std_logic;
	out1077                               :   OUT    std_logic;
	out1078                               :   OUT    std_logic;
	out1079                               :   OUT    std_logic;
	out1080                               :   OUT    std_logic;
	out1081                               :   OUT    std_logic;
	out1082                               :   OUT    std_logic;
	out1083                               :   OUT    std_logic;
	out1084                               :   OUT    std_logic;
	out1085                               :   OUT    std_logic;
	out1086                               :   OUT    std_logic;
	out1087                               :   OUT    std_logic;
	out1088                               :   OUT    std_logic;
	out1089                               :   OUT    std_logic;
	out1090                               :   OUT    std_logic;
	out1091                               :   OUT    std_logic;
	out1092                               :   OUT    std_logic;
	out1093                               :   OUT    std_logic;
	out1094                               :   OUT    std_logic;
	out1095                               :   OUT    std_logic;
	out1096                               :   OUT    std_logic;
	out1097                               :   OUT    std_logic;
	out1098                               :   OUT    std_logic;
	out1099                               :   OUT    std_logic;
	out1100                               :   OUT    std_logic;
	out1101                               :   OUT    std_logic;
	out1102                               :   OUT    std_logic;
	out1103                               :   OUT    std_logic;
	out1104                               :   OUT    std_logic;
	out1105                               :   OUT    std_logic;
	out1106                               :   OUT    std_logic;
	out1107                               :   OUT    std_logic;
	out1108                               :   OUT    std_logic;
	out1109                               :   OUT    std_logic;
	out1110                               :   OUT    std_logic;
	out1111                               :   OUT    std_logic;
	out1112                               :   OUT    std_logic;
	out1113                               :   OUT    std_logic;
	out1114                               :   OUT    std_logic;
	out1115                               :   OUT    std_logic;
	out1116                               :   OUT    std_logic;
	out1117                               :   OUT    std_logic;
	out1118                               :   OUT    std_logic;
	out1119                               :   OUT    std_logic;
	out1120                               :   OUT    std_logic;
	out1121                               :   OUT    std_logic;
	out1122                               :   OUT    std_logic;
	out1123                               :   OUT    std_logic;
	out1124                               :   OUT    std_logic;
	out1125                               :   OUT    std_logic;
	out1126                               :   OUT    std_logic;
	out1127                               :   OUT    std_logic;
	out1128                               :   OUT    std_logic;
	out1129                               :   OUT    std_logic;
	out1130                               :   OUT    std_logic;
	out1131                               :   OUT    std_logic;
	out1132                               :   OUT    std_logic;
	out1133                               :   OUT    std_logic;
	out1134                               :   OUT    std_logic;
	out1135                               :   OUT    std_logic;
	out1136                               :   OUT    std_logic;
	out1137                               :   OUT    std_logic;
	out1138                               :   OUT    std_logic;
	out1139                               :   OUT    std_logic;
	out1140                               :   OUT    std_logic;
	out1141                               :   OUT    std_logic;
	out1142                               :   OUT    std_logic;
	out1143                               :   OUT    std_logic;
	out1144                               :   OUT    std_logic;
	out1145                               :   OUT    std_logic;
	out1146                               :   OUT    std_logic;
	out1147                               :   OUT    std_logic;
	out1148                               :   OUT    std_logic;
	out1149                               :   OUT    std_logic;
	out1150                               :   OUT    std_logic;
	out1151                               :   OUT    std_logic;
	out1152                               :   OUT    std_logic;
	out1153                               :   OUT    std_logic;
	out1154                               :   OUT    std_logic;
	out1155                               :   OUT    std_logic;
	out1156                               :   OUT    std_logic;
	out1157                               :   OUT    std_logic;
	out1158                               :   OUT    std_logic;
	out1159                               :   OUT    std_logic;
	out1160                               :   OUT    std_logic;
	out1161                               :   OUT    std_logic;
	out1162                               :   OUT    std_logic;
	out1163                               :   OUT    std_logic;
	out1164                               :   OUT    std_logic;
	out1165                               :   OUT    std_logic;
	out1166                               :   OUT    std_logic;
	out1167                               :   OUT    std_logic;
	out1168                               :   OUT    std_logic;
	out1169                               :   OUT    std_logic;
	out1170                               :   OUT    std_logic;
	out1171                               :   OUT    std_logic;
	out1172                               :   OUT    std_logic;
	out1173                               :   OUT    std_logic;
	out1174                               :   OUT    std_logic;
	out1175                               :   OUT    std_logic;
	out1176                               :   OUT    std_logic;
	out1177                               :   OUT    std_logic;
	out1178                               :   OUT    std_logic;
	out1179                               :   OUT    std_logic;
	out1180                               :   OUT    std_logic;
	out1181                               :   OUT    std_logic;
	out1182                               :   OUT    std_logic;
	out1183                               :   OUT    std_logic;
	out1184                               :   OUT    std_logic;
	out1185                               :   OUT    std_logic;
	out1186                               :   OUT    std_logic;
	out1187                               :   OUT    std_logic;
	out1188                               :   OUT    std_logic;
	out1189                               :   OUT    std_logic;
	out1190                               :   OUT    std_logic;
	out1191                               :   OUT    std_logic;
	out1192                               :   OUT    std_logic;
	out1193                               :   OUT    std_logic;
	out1194                               :   OUT    std_logic;
	out1195                               :   OUT    std_logic;
	out1196                               :   OUT    std_logic;
	out1197                               :   OUT    std_logic;
	out1198                               :   OUT    std_logic;
	out1199                               :   OUT    std_logic;
	out1200                               :   OUT    std_logic;
	out1201                               :   OUT    std_logic;
	out1202                               :   OUT    std_logic;
	out1203                               :   OUT    std_logic;
	out1204                               :   OUT    std_logic;
	out1205                               :   OUT    std_logic;
	out1206                               :   OUT    std_logic;
	out1207                               :   OUT    std_logic;
	out1208                               :   OUT    std_logic;
	out1209                               :   OUT    std_logic;
	out1210                               :   OUT    std_logic;
	out1211                               :   OUT    std_logic;
	out1212                               :   OUT    std_logic;
	out1213                               :   OUT    std_logic;
	out1214                               :   OUT    std_logic;
	out1215                               :   OUT    std_logic;
	out1216                               :   OUT    std_logic;
	out1217                               :   OUT    std_logic;
	out1218                               :   OUT    std_logic;
	out1219                               :   OUT    std_logic;
	out1220                               :   OUT    std_logic;
	out1221                               :   OUT    std_logic;
	out1222                               :   OUT    std_logic;
	out1223                               :   OUT    std_logic;
	out1224                               :   OUT    std_logic;
	out1225                               :   OUT    std_logic;
	out1226                               :   OUT    std_logic;
	out1227                               :   OUT    std_logic;
	out1228                               :   OUT    std_logic;
	out1229                               :   OUT    std_logic;
	out1230                               :   OUT    std_logic;
	out1231                               :   OUT    std_logic;
	out1232                               :   OUT    std_logic;
	out1233                               :   OUT    std_logic;
	out1234                               :   OUT    std_logic;
	out1235                               :   OUT    std_logic;
	out1236                               :   OUT    std_logic;
	out1237                               :   OUT    std_logic;
	out1238                               :   OUT    std_logic;
	out1239                               :   OUT    std_logic;
	out1240                               :   OUT    std_logic;
	out1241                               :   OUT    std_logic;
	out1242                               :   OUT    std_logic;
	out1243                               :   OUT    std_logic;
	out1244                               :   OUT    std_logic;
	out1245                               :   OUT    std_logic;
	out1246                               :   OUT    std_logic;
	out1247                               :   OUT    std_logic;
	out1248                               :   OUT    std_logic;
	out1249                               :   OUT    std_logic;
	out1250                               :   OUT    std_logic;
	out1251                               :   OUT    std_logic;
	out1252                               :   OUT    std_logic;
	out1253                               :   OUT    std_logic;
	out1254                               :   OUT    std_logic;
	out1255                               :   OUT    std_logic;
	out1256                               :   OUT    std_logic;
	out1257                               :   OUT    std_logic;
	out1258                               :   OUT    std_logic;
	out1259                               :   OUT    std_logic;
	out1260                               :   OUT    std_logic;
	out1261                               :   OUT    std_logic;
	out1262                               :   OUT    std_logic;
	out1263                               :   OUT    std_logic;
	out1264                               :   OUT    std_logic;
	out1265                               :   OUT    std_logic;
	out1266                               :   OUT    std_logic;
	out1267                               :   OUT    std_logic;
	out1268                               :   OUT    std_logic;
	out1269                               :   OUT    std_logic;
	out1270                               :   OUT    std_logic;
	out1271                               :   OUT    std_logic;
	out1272                               :   OUT    std_logic;
	out1273                               :   OUT    std_logic;
	out1274                               :   OUT    std_logic;
	out1275                               :   OUT    std_logic;
	out1276                               :   OUT    std_logic;
	out1277                               :   OUT    std_logic;
	out1278                               :   OUT    std_logic;
	out1279                               :   OUT    std_logic;
	out1280                               :   OUT    std_logic;
	out1281                               :   OUT    std_logic;
	out1282                               :   OUT    std_logic;
	out1283                               :   OUT    std_logic;
	out1284                               :   OUT    std_logic;
	out1285                               :   OUT    std_logic;
	out1286                               :   OUT    std_logic;
	out1287                               :   OUT    std_logic;
	out1288                               :   OUT    std_logic;
	out1289                               :   OUT    std_logic;
	out1290                               :   OUT    std_logic;
	out1291                               :   OUT    std_logic;
	out1292                               :   OUT    std_logic;
	out1293                               :   OUT    std_logic;
	out1294                               :   OUT    std_logic;
	out1295                               :   OUT    std_logic;
	out1296                               :   OUT    std_logic;
	out1297                               :   OUT    std_logic;
	out1298                               :   OUT    std_logic;
	out1299                               :   OUT    std_logic;
	out1300                               :   OUT    std_logic;
	out1301                               :   OUT    std_logic;
	out1302                               :   OUT    std_logic;
	out1303                               :   OUT    std_logic;
	out1304                               :   OUT    std_logic;
	out1305                               :   OUT    std_logic;
	out1306                               :   OUT    std_logic;
	out1307                               :   OUT    std_logic;
	out1308                               :   OUT    std_logic;
	out1309                               :   OUT    std_logic;
	out1310                               :   OUT    std_logic;
	out1311                               :   OUT    std_logic;
	out1312                               :   OUT    std_logic;
	out1313                               :   OUT    std_logic;
	out1314                               :   OUT    std_logic;
	out1315                               :   OUT    std_logic;
	out1316                               :   OUT    std_logic;
	out1317                               :   OUT    std_logic;
	out1318                               :   OUT    std_logic;
	out1319                               :   OUT    std_logic;
	out1320                               :   OUT    std_logic;
	out1321                               :   OUT    std_logic;
	out1322                               :   OUT    std_logic;
	out1323                               :   OUT    std_logic;
	out1324                               :   OUT    std_logic;
	out1325                               :   OUT    std_logic;
	out1326                               :   OUT    std_logic;
	out1327                               :   OUT    std_logic;
	out1328                               :   OUT    std_logic;
	out1329                               :   OUT    std_logic;
	out1330                               :   OUT    std_logic;
	out1331                               :   OUT    std_logic;
	out1332                               :   OUT    std_logic;
	out1333                               :   OUT    std_logic;
	out1334                               :   OUT    std_logic;
	out1335                               :   OUT    std_logic;
	out1336                               :   OUT    std_logic;
	out1337                               :   OUT    std_logic;
	out1338                               :   OUT    std_logic;
	out1339                               :   OUT    std_logic;
	out1340                               :   OUT    std_logic;
	out1341                               :   OUT    std_logic;
	out1342                               :   OUT    std_logic;
	out1343                               :   OUT    std_logic;
	out1344                               :   OUT    std_logic;
	out1345                               :   OUT    std_logic;
	out1346                               :   OUT    std_logic;
	out1347                               :   OUT    std_logic;
	out1348                               :   OUT    std_logic;
	out1349                               :   OUT    std_logic;
	out1350                               :   OUT    std_logic;
	out1351                               :   OUT    std_logic;
	out1352                               :   OUT    std_logic;
	out1353                               :   OUT    std_logic;
	out1354                               :   OUT    std_logic;
	out1355                               :   OUT    std_logic;
	out1356                               :   OUT    std_logic;
	out1357                               :   OUT    std_logic;
	out1358                               :   OUT    std_logic;
	out1359                               :   OUT    std_logic;
	out1360                               :   OUT    std_logic;
	out1361                               :   OUT    std_logic;
	out1362                               :   OUT    std_logic;
	out1363                               :   OUT    std_logic;
	out1364                               :   OUT    std_logic;
	out1365                               :   OUT    std_logic;
	out1366                               :   OUT    std_logic;
	out1367                               :   OUT    std_logic;
	out1368                               :   OUT    std_logic;
	out1369                               :   OUT    std_logic;
	out1370                               :   OUT    std_logic;
	out1371                               :   OUT    std_logic;
	out1372                               :   OUT    std_logic;
	out1373                               :   OUT    std_logic;
	out1374                               :   OUT    std_logic;
	out1375                               :   OUT    std_logic;
	out1376                               :   OUT    std_logic;
	out1377                               :   OUT    std_logic;
	out1378                               :   OUT    std_logic;
	out1379                               :   OUT    std_logic;
	out1380                               :   OUT    std_logic;
	out1381                               :   OUT    std_logic;
	out1382                               :   OUT    std_logic;
	out1383                               :   OUT    std_logic;
	out1384                               :   OUT    std_logic;
	out1385                               :   OUT    std_logic;
	out1386                               :   OUT    std_logic;
	out1387                               :   OUT    std_logic;
	out1388                               :   OUT    std_logic;
	out1389                               :   OUT    std_logic;
	out1390                               :   OUT    std_logic;
	out1391                               :   OUT    std_logic;
	out1392                               :   OUT    std_logic;
	out1393                               :   OUT    std_logic;
	out1394                               :   OUT    std_logic;
	out1395                               :   OUT    std_logic;
	out1396                               :   OUT    std_logic;
	out1397                               :   OUT    std_logic;
	out1398                               :   OUT    std_logic;
	out1399                               :   OUT    std_logic;
	out1400                               :   OUT    std_logic;
	out1401                               :   OUT    std_logic;
	out1402                               :   OUT    std_logic;
	out1403                               :   OUT    std_logic;
	out1404                               :   OUT    std_logic;
	out1405                               :   OUT    std_logic;
	out1406                               :   OUT    std_logic;
	out1407                               :   OUT    std_logic;
	out1408                               :   OUT    std_logic;
	out1409                               :   OUT    std_logic;
	out1410                               :   OUT    std_logic;
	out1411                               :   OUT    std_logic;
	out1412                               :   OUT    std_logic;
	out1413                               :   OUT    std_logic;
	out1414                               :   OUT    std_logic;
	out1415                               :   OUT    std_logic;
	out1416                               :   OUT    std_logic;
	out1417                               :   OUT    std_logic;
	out1418                               :   OUT    std_logic;
	out1419                               :   OUT    std_logic;
	out1420                               :   OUT    std_logic;
	out1421                               :   OUT    std_logic;
	out1422                               :   OUT    std_logic;
	out1423                               :   OUT    std_logic;
	out1424                               :   OUT    std_logic;
	out1425                               :   OUT    std_logic;
	out1426                               :   OUT    std_logic;
	out1427                               :   OUT    std_logic;
	out1428                               :   OUT    std_logic;
	out1429                               :   OUT    std_logic;
	out1430                               :   OUT    std_logic;
	out1431                               :   OUT    std_logic;
	out1432                               :   OUT    std_logic;
	out1433                               :   OUT    std_logic;
	out1434                               :   OUT    std_logic;
	out1435                               :   OUT    std_logic;
	out1436                               :   OUT    std_logic;
	out1437                               :   OUT    std_logic;
	out1438                               :   OUT    std_logic;
	out1439                               :   OUT    std_logic;
	out1440                               :   OUT    std_logic;
	out1441                               :   OUT    std_logic;
	out1442                               :   OUT    std_logic;
	out1443                               :   OUT    std_logic;
	out1444                               :   OUT    std_logic;
	out1445                               :   OUT    std_logic;
	out1446                               :   OUT    std_logic;
	out1447                               :   OUT    std_logic;
	out1448                               :   OUT    std_logic;
	out1449                               :   OUT    std_logic;
	out1450                               :   OUT    std_logic;
	out1451                               :   OUT    std_logic;
	out1452                               :   OUT    std_logic;
	out1453                               :   OUT    std_logic;
	out1454                               :   OUT    std_logic;
	out1455                               :   OUT    std_logic;
	out1456                               :   OUT    std_logic;
	out1457                               :   OUT    std_logic;
	out1458                               :   OUT    std_logic;
	out1459                               :   OUT    std_logic;
	out1460                               :   OUT    std_logic;
	out1461                               :   OUT    std_logic;
	out1462                               :   OUT    std_logic;
	out1463                               :   OUT    std_logic;
	out1464                               :   OUT    std_logic;
	out1465                               :   OUT    std_logic;
	out1466                               :   OUT    std_logic;
	out1467                               :   OUT    std_logic;
	out1468                               :   OUT    std_logic;
	out1469                               :   OUT    std_logic;
	out1470                               :   OUT    std_logic;
	out1471                               :   OUT    std_logic;
	out1472                               :   OUT    std_logic;
	out1473                               :   OUT    std_logic;
	out1474                               :   OUT    std_logic;
	out1475                               :   OUT    std_logic;
	out1476                               :   OUT    std_logic;
	out1477                               :   OUT    std_logic;
	out1478                               :   OUT    std_logic;
	out1479                               :   OUT    std_logic;
	out1480                               :   OUT    std_logic;
	out1481                               :   OUT    std_logic;
	out1482                               :   OUT    std_logic;
	out1483                               :   OUT    std_logic;
	out1484                               :   OUT    std_logic;
	out1485                               :   OUT    std_logic;
	out1486                               :   OUT    std_logic;
	out1487                               :   OUT    std_logic;
	out1488                               :   OUT    std_logic;
	out1489                               :   OUT    std_logic;
	out1490                               :   OUT    std_logic;
	out1491                               :   OUT    std_logic;
	out1492                               :   OUT    std_logic;
	out1493                               :   OUT    std_logic;
	out1494                               :   OUT    std_logic;
	out1495                               :   OUT    std_logic;
	out1496                               :   OUT    std_logic;
	out1497                               :   OUT    std_logic;
	out1498                               :   OUT    std_logic;
	out1499                               :   OUT    std_logic;
	out1500                               :   OUT    std_logic;
	out1501                               :   OUT    std_logic;
	out1502                               :   OUT    std_logic;
	out1503                               :   OUT    std_logic;
	out1504                               :   OUT    std_logic;
	out1505                               :   OUT    std_logic;
	out1506                               :   OUT    std_logic;
	out1507                               :   OUT    std_logic;
	out1508                               :   OUT    std_logic;
	out1509                               :   OUT    std_logic;
	out1510                               :   OUT    std_logic;
	out1511                               :   OUT    std_logic;
	out1512                               :   OUT    std_logic;
	out1513                               :   OUT    std_logic;
	out1514                               :   OUT    std_logic;
	out1515                               :   OUT    std_logic;
	out1516                               :   OUT    std_logic;
	out1517                               :   OUT    std_logic;
	out1518                               :   OUT    std_logic;
	out1519                               :   OUT    std_logic;
	out1520                               :   OUT    std_logic;
	out1521                               :   OUT    std_logic;
	out1522                               :   OUT    std_logic;
	out1523                               :   OUT    std_logic;
	out1524                               :   OUT    std_logic;
	out1525                               :   OUT    std_logic;
	out1526                               :   OUT    std_logic;
	out1527                               :   OUT    std_logic;
	out1528                               :   OUT    std_logic;
	out1529                               :   OUT    std_logic;
	out1530                               :   OUT    std_logic;
	out1531                               :   OUT    std_logic;
	out1532                               :   OUT    std_logic;
	out1533                               :   OUT    std_logic;
	out1534                               :   OUT    std_logic;
	out1535                               :   OUT    std_logic;
	out1536                               :   OUT    std_logic;
	out1537                               :   OUT    std_logic;
	out1538                               :   OUT    std_logic;
	out1539                               :   OUT    std_logic;
	out1540                               :   OUT    std_logic;
	out1541                               :   OUT    std_logic;
	out1542                               :   OUT    std_logic;
	out1543                               :   OUT    std_logic;
	out1544                               :   OUT    std_logic;
	out1545                               :   OUT    std_logic;
	out1546                               :   OUT    std_logic;
	out1547                               :   OUT    std_logic;
	out1548                               :   OUT    std_logic;
	out1549                               :   OUT    std_logic;
	out1550                               :   OUT    std_logic;
	out1551                               :   OUT    std_logic;
	out1552                               :   OUT    std_logic;
	out1553                               :   OUT    std_logic;
	out1554                               :   OUT    std_logic;
	out1555                               :   OUT    std_logic;
	out1556                               :   OUT    std_logic;
	out1557                               :   OUT    std_logic;
	out1558                               :   OUT    std_logic;
	out1559                               :   OUT    std_logic;
	out1560                               :   OUT    std_logic;
	out1561                               :   OUT    std_logic;
	out1562                               :   OUT    std_logic;
	out1563                               :   OUT    std_logic;
	out1564                               :   OUT    std_logic;
	out1565                               :   OUT    std_logic;
	out1566                               :   OUT    std_logic;
	out1567                               :   OUT    std_logic;
	out1568                               :   OUT    std_logic;
	out1569                               :   OUT    std_logic;
	out1570                               :   OUT    std_logic;
	out1571                               :   OUT    std_logic;
	out1572                               :   OUT    std_logic;
	out1573                               :   OUT    std_logic;
	out1574                               :   OUT    std_logic;
	out1575                               :   OUT    std_logic;
	out1576                               :   OUT    std_logic;
	out1577                               :   OUT    std_logic;
	out1578                               :   OUT    std_logic;
	out1579                               :   OUT    std_logic;
	out1580                               :   OUT    std_logic;
	out1581                               :   OUT    std_logic;
	out1582                               :   OUT    std_logic;
	out1583                               :   OUT    std_logic;
	out1584                               :   OUT    std_logic;
	out1585                               :   OUT    std_logic;
	out1586                               :   OUT    std_logic;
	out1587                               :   OUT    std_logic;
	out1588                               :   OUT    std_logic;
	out1589                               :   OUT    std_logic;
	out1590                               :   OUT    std_logic;
	out1591                               :   OUT    std_logic;
	out1592                               :   OUT    std_logic;
	out1593                               :   OUT    std_logic;
	out1594                               :   OUT    std_logic;
	out1595                               :   OUT    std_logic;
	out1596                               :   OUT    std_logic;
	out1597                               :   OUT    std_logic;
	out1598                               :   OUT    std_logic;
	out1599                               :   OUT    std_logic;
	out1600                               :   OUT    std_logic;
	out1601                               :   OUT    std_logic;
	out1602                               :   OUT    std_logic;
	out1603                               :   OUT    std_logic;
	out1604                               :   OUT    std_logic;
	out1605                               :   OUT    std_logic;
	out1606                               :   OUT    std_logic;
	out1607                               :   OUT    std_logic;
	out1608                               :   OUT    std_logic;
	out1609                               :   OUT    std_logic;
	out1610                               :   OUT    std_logic;
	out1611                               :   OUT    std_logic;
	out1612                               :   OUT    std_logic;
	out1613                               :   OUT    std_logic;
	out1614                               :   OUT    std_logic;
	out1615                               :   OUT    std_logic;
	out1616                               :   OUT    std_logic;
	out1617                               :   OUT    std_logic;
	out1618                               :   OUT    std_logic;
	out1619                               :   OUT    std_logic;
	out1620                               :   OUT    std_logic;
	out1621                               :   OUT    std_logic;
	out1622                               :   OUT    std_logic;
	out1623                               :   OUT    std_logic;
	out1624                               :   OUT    std_logic;
	out1625                               :   OUT    std_logic;
	out1626                               :   OUT    std_logic;
	out1627                               :   OUT    std_logic;
	out1628                               :   OUT    std_logic;
	out1629                               :   OUT    std_logic;
	out1630                               :   OUT    std_logic;
	out1631                               :   OUT    std_logic;
	out1632                               :   OUT    std_logic;
	out1633                               :   OUT    std_logic;
	out1634                               :   OUT    std_logic;
	out1635                               :   OUT    std_logic;
	out1636                               :   OUT    std_logic;
	out1637                               :   OUT    std_logic;
	out1638                               :   OUT    std_logic;
	out1639                               :   OUT    std_logic;
	out1640                               :   OUT    std_logic;
	out1641                               :   OUT    std_logic;
	out1642                               :   OUT    std_logic;
	out1643                               :   OUT    std_logic;
	out1644                               :   OUT    std_logic;
	out1645                               :   OUT    std_logic;
	out1646                               :   OUT    std_logic;
	out1647                               :   OUT    std_logic;
	out1648                               :   OUT    std_logic;
	out1649                               :   OUT    std_logic;
	out1650                               :   OUT    std_logic;
	out1651                               :   OUT    std_logic;
	out1652                               :   OUT    std_logic;
	out1653                               :   OUT    std_logic;
	out1654                               :   OUT    std_logic;
	out1655                               :   OUT    std_logic;
	out1656                               :   OUT    std_logic;
	out1657                               :   OUT    std_logic;
	out1658                               :   OUT    std_logic;
	out1659                               :   OUT    std_logic;
	out1660                               :   OUT    std_logic;
	out1661                               :   OUT    std_logic;
	out1662                               :   OUT    std_logic;
	out1663                               :   OUT    std_logic;
	out1664                               :   OUT    std_logic;
	out1665                               :   OUT    std_logic;
	out1666                               :   OUT    std_logic;
	out1667                               :   OUT    std_logic;
	out1668                               :   OUT    std_logic;
	out1669                               :   OUT    std_logic;
	out1670                               :   OUT    std_logic;
	out1671                               :   OUT    std_logic;
	out1672                               :   OUT    std_logic;
	out1673                               :   OUT    std_logic;
	out1674                               :   OUT    std_logic;
	out1675                               :   OUT    std_logic;
	out1676                               :   OUT    std_logic;
	out1677                               :   OUT    std_logic;
	out1678                               :   OUT    std_logic;
	out1679                               :   OUT    std_logic;
	out1680                               :   OUT    std_logic;
	out1681                               :   OUT    std_logic;
	out1682                               :   OUT    std_logic;
	out1683                               :   OUT    std_logic;
	out1684                               :   OUT    std_logic;
	out1685                               :   OUT    std_logic;
	out1686                               :   OUT    std_logic;
	out1687                               :   OUT    std_logic;
	out1688                               :   OUT    std_logic;
	out1689                               :   OUT    std_logic;
	out1690                               :   OUT    std_logic;
	out1691                               :   OUT    std_logic;
	out1692                               :   OUT    std_logic;
	out1693                               :   OUT    std_logic;
	out1694                               :   OUT    std_logic;
	out1695                               :   OUT    std_logic;
	out1696                               :   OUT    std_logic;
	out1697                               :   OUT    std_logic;
	out1698                               :   OUT    std_logic;
	out1699                               :   OUT    std_logic;
	out1700                               :   OUT    std_logic;
	out1701                               :   OUT    std_logic;
	out1702                               :   OUT    std_logic;
	out1703                               :   OUT    std_logic;
	out1704                               :   OUT    std_logic;
	out1705                               :   OUT    std_logic;
	out1706                               :   OUT    std_logic;
	out1707                               :   OUT    std_logic;
	out1708                               :   OUT    std_logic;
	out1709                               :   OUT    std_logic;
	out1710                               :   OUT    std_logic;
	out1711                               :   OUT    std_logic;
	out1712                               :   OUT    std_logic;
	out1713                               :   OUT    std_logic;
	out1714                               :   OUT    std_logic;
	out1715                               :   OUT    std_logic;
	out1716                               :   OUT    std_logic;
	out1717                               :   OUT    std_logic;
	out1718                               :   OUT    std_logic;
	out1719                               :   OUT    std_logic;
	out1720                               :   OUT    std_logic;
	out1721                               :   OUT    std_logic;
	out1722                               :   OUT    std_logic;
	out1723                               :   OUT    std_logic;
	out1724                               :   OUT    std_logic;
	out1725                               :   OUT    std_logic;
	out1726                               :   OUT    std_logic;
	out1727                               :   OUT    std_logic;
	out1728                               :   OUT    std_logic;
	out1729                               :   OUT    std_logic;
	out1730                               :   OUT    std_logic;
	out1731                               :   OUT    std_logic;
	out1732                               :   OUT    std_logic;
	out1733                               :   OUT    std_logic;
	out1734                               :   OUT    std_logic;
	out1735                               :   OUT    std_logic;
	out1736                               :   OUT    std_logic;
	out1737                               :   OUT    std_logic;
	out1738                               :   OUT    std_logic;
	out1739                               :   OUT    std_logic;
	out1740                               :   OUT    std_logic;
	out1741                               :   OUT    std_logic;
	out1742                               :   OUT    std_logic;
	out1743                               :   OUT    std_logic;
	out1744                               :   OUT    std_logic;
	out1745                               :   OUT    std_logic;
	out1746                               :   OUT    std_logic;
	out1747                               :   OUT    std_logic;
	out1748                               :   OUT    std_logic;
	out1749                               :   OUT    std_logic;
	out1750                               :   OUT    std_logic;
	out1751                               :   OUT    std_logic;
	out1752                               :   OUT    std_logic;
	out1753                               :   OUT    std_logic;
	out1754                               :   OUT    std_logic;
	out1755                               :   OUT    std_logic;
	out1756                               :   OUT    std_logic;
	out1757                               :   OUT    std_logic;
	out1758                               :   OUT    std_logic;
	out1759                               :   OUT    std_logic;
	out1760                               :   OUT    std_logic;
	out1761                               :   OUT    std_logic;
	out1762                               :   OUT    std_logic;
	out1763                               :   OUT    std_logic;
	out1764                               :   OUT    std_logic;
	out1765                               :   OUT    std_logic;
	out1766                               :   OUT    std_logic;
	out1767                               :   OUT    std_logic;
	out1768                               :   OUT    std_logic;
	out1769                               :   OUT    std_logic;
	out1770                               :   OUT    std_logic;
	out1771                               :   OUT    std_logic;
	out1772                               :   OUT    std_logic;
	out1773                               :   OUT    std_logic;
	out1774                               :   OUT    std_logic;
	out1775                               :   OUT    std_logic;
	out1776                               :   OUT    std_logic;
	out1777                               :   OUT    std_logic;
	out1778                               :   OUT    std_logic;
	out1779                               :   OUT    std_logic;
	out1780                               :   OUT    std_logic;
	out1781                               :   OUT    std_logic;
	out1782                               :   OUT    std_logic;
	out1783                               :   OUT    std_logic;
	out1784                               :   OUT    std_logic;
	out1785                               :   OUT    std_logic;
	out1786                               :   OUT    std_logic;
	out1787                               :   OUT    std_logic;
	out1788                               :   OUT    std_logic;
	out1789                               :   OUT    std_logic;
	out1790                               :   OUT    std_logic;
	out1791                               :   OUT    std_logic;
	out1792                               :   OUT    std_logic;
	out1793                               :   OUT    std_logic;
	out1794                               :   OUT    std_logic;
	out1795                               :   OUT    std_logic;
	out1796                               :   OUT    std_logic;
	out1797                               :   OUT    std_logic;
	out1798                               :   OUT    std_logic;
	out1799                               :   OUT    std_logic;
	out1800                               :   OUT    std_logic;
	out1801                               :   OUT    std_logic;
	out1802                               :   OUT    std_logic;
	out1803                               :   OUT    std_logic;
	out1804                               :   OUT    std_logic;
	out1805                               :   OUT    std_logic;
	out1806                               :   OUT    std_logic;
	out1807                               :   OUT    std_logic;
	out1808                               :   OUT    std_logic;
	out1809                               :   OUT    std_logic;
	out1810                               :   OUT    std_logic;
	out1811                               :   OUT    std_logic;
	out1812                               :   OUT    std_logic;
	out1813                               :   OUT    std_logic;
	out1814                               :   OUT    std_logic;
	out1815                               :   OUT    std_logic;
	out1816                               :   OUT    std_logic;
	out1817                               :   OUT    std_logic;
	out1818                               :   OUT    std_logic;
	out1819                               :   OUT    std_logic;
	out1820                               :   OUT    std_logic;
	out1821                               :   OUT    std_logic;
	out1822                               :   OUT    std_logic;
	out1823                               :   OUT    std_logic;
	out1824                               :   OUT    std_logic;
	out1825                               :   OUT    std_logic;
	out1826                               :   OUT    std_logic;
	out1827                               :   OUT    std_logic;
	out1828                               :   OUT    std_logic;
	out1829                               :   OUT    std_logic;
	out1830                               :   OUT    std_logic;
	out1831                               :   OUT    std_logic;
	out1832                               :   OUT    std_logic;
	out1833                               :   OUT    std_logic;
	out1834                               :   OUT    std_logic;
	out1835                               :   OUT    std_logic;
	out1836                               :   OUT    std_logic;
	out1837                               :   OUT    std_logic;
	out1838                               :   OUT    std_logic;
	out1839                               :   OUT    std_logic;
	out1840                               :   OUT    std_logic;
	out1841                               :   OUT    std_logic;
	out1842                               :   OUT    std_logic;
	out1843                               :   OUT    std_logic;
	out1844                               :   OUT    std_logic;
	out1845                               :   OUT    std_logic;
	out1846                               :   OUT    std_logic;
	out1847                               :   OUT    std_logic;
	out1848                               :   OUT    std_logic;
	out1849                               :   OUT    std_logic;
	out1850                               :   OUT    std_logic;
	out1851                               :   OUT    std_logic;
	out1852                               :   OUT    std_logic;
	out1853                               :   OUT    std_logic;
	out1854                               :   OUT    std_logic;
	out1855                               :   OUT    std_logic;
	out1856                               :   OUT    std_logic;
	out1857                               :   OUT    std_logic;
	out1858                               :   OUT    std_logic;
	out1859                               :   OUT    std_logic;
	out1860                               :   OUT    std_logic;
	out1861                               :   OUT    std_logic;
	out1862                               :   OUT    std_logic;
	out1863                               :   OUT    std_logic;
	out1864                               :   OUT    std_logic;
	out1865                               :   OUT    std_logic;
	out1866                               :   OUT    std_logic;
	out1867                               :   OUT    std_logic;
	out1868                               :   OUT    std_logic;
	out1869                               :   OUT    std_logic;
	out1870                               :   OUT    std_logic;
	out1871                               :   OUT    std_logic;
	out1872                               :   OUT    std_logic;
	out1873                               :   OUT    std_logic;
	out1874                               :   OUT    std_logic;
	out1875                               :   OUT    std_logic;
	out1876                               :   OUT    std_logic;
	out1877                               :   OUT    std_logic;
	out1878                               :   OUT    std_logic;
	out1879                               :   OUT    std_logic;
	out1880                               :   OUT    std_logic;
	out1881                               :   OUT    std_logic;
	out1882                               :   OUT    std_logic;
	out1883                               :   OUT    std_logic;
	out1884                               :   OUT    std_logic;
	out1885                               :   OUT    std_logic;
	out1886                               :   OUT    std_logic;
	out1887                               :   OUT    std_logic;
	out1888                               :   OUT    std_logic;
	out1889                               :   OUT    std_logic;
	out1890                               :   OUT    std_logic;
	out1891                               :   OUT    std_logic;
	out1892                               :   OUT    std_logic;
	out1893                               :   OUT    std_logic;
	out1894                               :   OUT    std_logic;
	out1895                               :   OUT    std_logic;
	out1896                               :   OUT    std_logic;
	out1897                               :   OUT    std_logic;
	out1898                               :   OUT    std_logic;
	out1899                               :   OUT    std_logic;
	out1900                               :   OUT    std_logic;
	out1901                               :   OUT    std_logic;
	out1902                               :   OUT    std_logic;
	out1903                               :   OUT    std_logic;
	out1904                               :   OUT    std_logic;
	out1905                               :   OUT    std_logic;
	out1906                               :   OUT    std_logic;
	out1907                               :   OUT    std_logic;
	out1908                               :   OUT    std_logic;
	out1909                               :   OUT    std_logic;
	out1910                               :   OUT    std_logic;
	out1911                               :   OUT    std_logic;
	out1912                               :   OUT    std_logic;
	out1913                               :   OUT    std_logic;
	out1914                               :   OUT    std_logic;
	out1915                               :   OUT    std_logic;
	out1916                               :   OUT    std_logic;
	out1917                               :   OUT    std_logic;
	out1918                               :   OUT    std_logic;
	out1919                               :   OUT    std_logic;
	out1920                               :   OUT    std_logic;
	out1921                               :   OUT    std_logic;
	out1922                               :   OUT    std_logic;
	out1923                               :   OUT    std_logic;
	out1924                               :   OUT    std_logic;
	out1925                               :   OUT    std_logic;
	out1926                               :   OUT    std_logic;
	out1927                               :   OUT    std_logic;
	out1928                               :   OUT    std_logic;
	out1929                               :   OUT    std_logic;
	out1930                               :   OUT    std_logic;
	out1931                               :   OUT    std_logic;
	out1932                               :   OUT    std_logic;
	out1933                               :   OUT    std_logic;
	out1934                               :   OUT    std_logic;
	out1935                               :   OUT    std_logic;
	out1936                               :   OUT    std_logic;
	out1937                               :   OUT    std_logic;
	out1938                               :   OUT    std_logic;
	out1939                               :   OUT    std_logic;
	out1940                               :   OUT    std_logic;
	out1941                               :   OUT    std_logic;
	out1942                               :   OUT    std_logic;
	out1943                               :   OUT    std_logic;
	out1944                               :   OUT    std_logic;
	out1945                               :   OUT    std_logic;
	out1946                               :   OUT    std_logic;
	out1947                               :   OUT    std_logic;
	out1948                               :   OUT    std_logic;
	out1949                               :   OUT    std_logic;
	out1950                               :   OUT    std_logic;
	out1951                               :   OUT    std_logic;
	out1952                               :   OUT    std_logic;
	out1953                               :   OUT    std_logic;
	out1954                               :   OUT    std_logic;
	out1955                               :   OUT    std_logic;
	out1956                               :   OUT    std_logic;
	out1957                               :   OUT    std_logic;
	out1958                               :   OUT    std_logic;
	out1959                               :   OUT    std_logic;
	out1960                               :   OUT    std_logic;
	out1961                               :   OUT    std_logic;
	out1962                               :   OUT    std_logic;
	out1963                               :   OUT    std_logic;
	out1964                               :   OUT    std_logic;
	out1965                               :   OUT    std_logic;
	out1966                               :   OUT    std_logic;
	out1967                               :   OUT    std_logic;
	out1968                               :   OUT    std_logic;
	out1969                               :   OUT    std_logic;
	out1970                               :   OUT    std_logic;
	out1971                               :   OUT    std_logic;
	out1972                               :   OUT    std_logic;
	out1973                               :   OUT    std_logic;
	out1974                               :   OUT    std_logic;
	out1975                               :   OUT    std_logic;
	out1976                               :   OUT    std_logic;
	out1977                               :   OUT    std_logic;
	out1978                               :   OUT    std_logic;
	out1979                               :   OUT    std_logic;
	out1980                               :   OUT    std_logic;
	out1981                               :   OUT    std_logic;
	out1982                               :   OUT    std_logic;
	out1983                               :   OUT    std_logic;
	out1984                               :   OUT    std_logic;
	out1985                               :   OUT    std_logic;
	out1986                               :   OUT    std_logic;
	out1987                               :   OUT    std_logic;
	out1988                               :   OUT    std_logic;
	out1989                               :   OUT    std_logic;
	out1990                               :   OUT    std_logic;
	out1991                               :   OUT    std_logic;
	out1992                               :   OUT    std_logic;
	out1993                               :   OUT    std_logic;
	out1994                               :   OUT    std_logic;
	out1995                               :   OUT    std_logic;
	out1996                               :   OUT    std_logic;
	out1997                               :   OUT    std_logic;
	out1998                               :   OUT    std_logic;
	out1999                               :   OUT    std_logic;
	out2000                               :   OUT    std_logic;
	out2001                               :   OUT    std_logic;
	out2002                               :   OUT    std_logic;
	out2003                               :   OUT    std_logic;
	out2004                               :   OUT    std_logic;
	out2005                               :   OUT    std_logic;
	out2006                               :   OUT    std_logic;
	out2007                               :   OUT    std_logic;
	out2008                               :   OUT    std_logic;
	out2009                               :   OUT    std_logic;
	out2010                               :   OUT    std_logic;
	out2011                               :   OUT    std_logic;
	out2012                               :   OUT    std_logic;
	out2013                               :   OUT    std_logic;
	out2014                               :   OUT    std_logic;
	out2015                               :   OUT    std_logic;
	out2016                               :   OUT    std_logic;
	out2017                               :   OUT    std_logic;
	out2018                               :   OUT    std_logic;
	out2019                               :   OUT    std_logic;
	out2020                               :   OUT    std_logic;
	out2021                               :   OUT    std_logic;
	out2022                               :   OUT    std_logic;
	out2023                               :   OUT    std_logic;
	out2024                               :   OUT    std_logic;
	out2025                               :   OUT    std_logic;
	out2026                               :   OUT    std_logic;
	out2027                               :   OUT    std_logic;
	out2028                               :   OUT    std_logic;
	out2029                               :   OUT    std_logic;
	out2030                               :   OUT    std_logic;
	out2031                               :   OUT    std_logic;
	out2032                               :   OUT    std_logic;
	out2033                               :   OUT    std_logic;
	out2034                               :   OUT    std_logic;
	out2035                               :   OUT    std_logic;
	out2036                               :   OUT    std_logic;
	out2037                               :   OUT    std_logic;
	out2038                               :   OUT    std_logic;
	out2039                               :   OUT    std_logic;
	out2040                               :   OUT    std_logic;
	out2041                               :   OUT    std_logic;
	out2042                               :   OUT    std_logic;
	out2043                               :   OUT    std_logic;
	out2044                               :   OUT    std_logic;
	out2045                               :   OUT    std_logic;
	out2046                               :   OUT    std_logic;
	out2047                               :   OUT    std_logic;
	out2048                               :   OUT    std_logic
	);
END encoderN2048;

ARCHITECTURE rtl OF encoderN2048 IS

  SIGNAL Logical_Operator_out1_out1            : std_logic;
  SIGNAL Logical_Operator_out2_out1            : std_logic;
  SIGNAL Logical_Operator_out3_out1            : std_logic;
  SIGNAL Logical_Operator_out4_out1            : std_logic;
  SIGNAL Logical_Operator_out5_out1            : std_logic;
  SIGNAL Logical_Operator_out6_out1            : std_logic;
  SIGNAL Logical_Operator_out7_out1            : std_logic;
  SIGNAL Logical_Operator_out8_out1            : std_logic;
  SIGNAL Logical_Operator_out9_out1            : std_logic;
  SIGNAL Logical_Operator_out10_out1            : std_logic;
  SIGNAL Logical_Operator_out11_out1            : std_logic;
  SIGNAL Logical_Operator_out12_out1            : std_logic;
  SIGNAL Logical_Operator_out13_out1            : std_logic;
  SIGNAL Logical_Operator_out14_out1            : std_logic;
  SIGNAL Logical_Operator_out15_out1            : std_logic;
  SIGNAL Logical_Operator_out16_out1            : std_logic;
  SIGNAL Logical_Operator_out17_out1            : std_logic;
  SIGNAL Logical_Operator_out18_out1            : std_logic;
  SIGNAL Logical_Operator_out19_out1            : std_logic;
  SIGNAL Logical_Operator_out20_out1            : std_logic;
  SIGNAL Logical_Operator_out21_out1            : std_logic;
  SIGNAL Logical_Operator_out22_out1            : std_logic;
  SIGNAL Logical_Operator_out23_out1            : std_logic;
  SIGNAL Logical_Operator_out24_out1            : std_logic;
  SIGNAL Logical_Operator_out25_out1            : std_logic;
  SIGNAL Logical_Operator_out26_out1            : std_logic;
  SIGNAL Logical_Operator_out27_out1            : std_logic;
  SIGNAL Logical_Operator_out28_out1            : std_logic;
  SIGNAL Logical_Operator_out29_out1            : std_logic;
  SIGNAL Logical_Operator_out30_out1            : std_logic;
  SIGNAL Logical_Operator_out31_out1            : std_logic;
  SIGNAL Logical_Operator_out32_out1            : std_logic;
  SIGNAL Logical_Operator_out33_out1            : std_logic;
  SIGNAL Logical_Operator_out34_out1            : std_logic;
  SIGNAL Logical_Operator_out35_out1            : std_logic;
  SIGNAL Logical_Operator_out36_out1            : std_logic;
  SIGNAL Logical_Operator_out37_out1            : std_logic;
  SIGNAL Logical_Operator_out38_out1            : std_logic;
  SIGNAL Logical_Operator_out39_out1            : std_logic;
  SIGNAL Logical_Operator_out40_out1            : std_logic;
  SIGNAL Logical_Operator_out41_out1            : std_logic;
  SIGNAL Logical_Operator_out42_out1            : std_logic;
  SIGNAL Logical_Operator_out43_out1            : std_logic;
  SIGNAL Logical_Operator_out44_out1            : std_logic;
  SIGNAL Logical_Operator_out45_out1            : std_logic;
  SIGNAL Logical_Operator_out46_out1            : std_logic;
  SIGNAL Logical_Operator_out47_out1            : std_logic;
  SIGNAL Logical_Operator_out48_out1            : std_logic;
  SIGNAL Logical_Operator_out49_out1            : std_logic;
  SIGNAL Logical_Operator_out50_out1            : std_logic;
  SIGNAL Logical_Operator_out51_out1            : std_logic;
  SIGNAL Logical_Operator_out52_out1            : std_logic;
  SIGNAL Logical_Operator_out53_out1            : std_logic;
  SIGNAL Logical_Operator_out54_out1            : std_logic;
  SIGNAL Logical_Operator_out55_out1            : std_logic;
  SIGNAL Logical_Operator_out56_out1            : std_logic;
  SIGNAL Logical_Operator_out57_out1            : std_logic;
  SIGNAL Logical_Operator_out58_out1            : std_logic;
  SIGNAL Logical_Operator_out59_out1            : std_logic;
  SIGNAL Logical_Operator_out60_out1            : std_logic;
  SIGNAL Logical_Operator_out61_out1            : std_logic;
  SIGNAL Logical_Operator_out62_out1            : std_logic;
  SIGNAL Logical_Operator_out63_out1            : std_logic;
  SIGNAL Logical_Operator_out64_out1            : std_logic;
  SIGNAL Logical_Operator_out65_out1            : std_logic;
  SIGNAL Logical_Operator_out66_out1            : std_logic;
  SIGNAL Logical_Operator_out67_out1            : std_logic;
  SIGNAL Logical_Operator_out68_out1            : std_logic;
  SIGNAL Logical_Operator_out69_out1            : std_logic;
  SIGNAL Logical_Operator_out70_out1            : std_logic;
  SIGNAL Logical_Operator_out71_out1            : std_logic;
  SIGNAL Logical_Operator_out72_out1            : std_logic;
  SIGNAL Logical_Operator_out73_out1            : std_logic;
  SIGNAL Logical_Operator_out74_out1            : std_logic;
  SIGNAL Logical_Operator_out75_out1            : std_logic;
  SIGNAL Logical_Operator_out76_out1            : std_logic;
  SIGNAL Logical_Operator_out77_out1            : std_logic;
  SIGNAL Logical_Operator_out78_out1            : std_logic;
  SIGNAL Logical_Operator_out79_out1            : std_logic;
  SIGNAL Logical_Operator_out80_out1            : std_logic;
  SIGNAL Logical_Operator_out81_out1            : std_logic;
  SIGNAL Logical_Operator_out82_out1            : std_logic;
  SIGNAL Logical_Operator_out83_out1            : std_logic;
  SIGNAL Logical_Operator_out84_out1            : std_logic;
  SIGNAL Logical_Operator_out85_out1            : std_logic;
  SIGNAL Logical_Operator_out86_out1            : std_logic;
  SIGNAL Logical_Operator_out87_out1            : std_logic;
  SIGNAL Logical_Operator_out88_out1            : std_logic;
  SIGNAL Logical_Operator_out89_out1            : std_logic;
  SIGNAL Logical_Operator_out90_out1            : std_logic;
  SIGNAL Logical_Operator_out91_out1            : std_logic;
  SIGNAL Logical_Operator_out92_out1            : std_logic;
  SIGNAL Logical_Operator_out93_out1            : std_logic;
  SIGNAL Logical_Operator_out94_out1            : std_logic;
  SIGNAL Logical_Operator_out95_out1            : std_logic;
  SIGNAL Logical_Operator_out96_out1            : std_logic;
  SIGNAL Logical_Operator_out97_out1            : std_logic;
  SIGNAL Logical_Operator_out98_out1            : std_logic;
  SIGNAL Logical_Operator_out99_out1            : std_logic;
  SIGNAL Logical_Operator_out100_out1            : std_logic;
  SIGNAL Logical_Operator_out101_out1            : std_logic;
  SIGNAL Logical_Operator_out102_out1            : std_logic;
  SIGNAL Logical_Operator_out103_out1            : std_logic;
  SIGNAL Logical_Operator_out104_out1            : std_logic;
  SIGNAL Logical_Operator_out105_out1            : std_logic;
  SIGNAL Logical_Operator_out106_out1            : std_logic;
  SIGNAL Logical_Operator_out107_out1            : std_logic;
  SIGNAL Logical_Operator_out108_out1            : std_logic;
  SIGNAL Logical_Operator_out109_out1            : std_logic;
  SIGNAL Logical_Operator_out110_out1            : std_logic;
  SIGNAL Logical_Operator_out111_out1            : std_logic;
  SIGNAL Logical_Operator_out112_out1            : std_logic;
  SIGNAL Logical_Operator_out113_out1            : std_logic;
  SIGNAL Logical_Operator_out114_out1            : std_logic;
  SIGNAL Logical_Operator_out115_out1            : std_logic;
  SIGNAL Logical_Operator_out116_out1            : std_logic;
  SIGNAL Logical_Operator_out117_out1            : std_logic;
  SIGNAL Logical_Operator_out118_out1            : std_logic;
  SIGNAL Logical_Operator_out119_out1            : std_logic;
  SIGNAL Logical_Operator_out120_out1            : std_logic;
  SIGNAL Logical_Operator_out121_out1            : std_logic;
  SIGNAL Logical_Operator_out122_out1            : std_logic;
  SIGNAL Logical_Operator_out123_out1            : std_logic;
  SIGNAL Logical_Operator_out124_out1            : std_logic;
  SIGNAL Logical_Operator_out125_out1            : std_logic;
  SIGNAL Logical_Operator_out126_out1            : std_logic;
  SIGNAL Logical_Operator_out127_out1            : std_logic;
  SIGNAL Logical_Operator_out128_out1            : std_logic;
  SIGNAL Logical_Operator_out129_out1            : std_logic;
  SIGNAL Logical_Operator_out130_out1            : std_logic;
  SIGNAL Logical_Operator_out131_out1            : std_logic;
  SIGNAL Logical_Operator_out132_out1            : std_logic;
  SIGNAL Logical_Operator_out133_out1            : std_logic;
  SIGNAL Logical_Operator_out134_out1            : std_logic;
  SIGNAL Logical_Operator_out135_out1            : std_logic;
  SIGNAL Logical_Operator_out136_out1            : std_logic;
  SIGNAL Logical_Operator_out137_out1            : std_logic;
  SIGNAL Logical_Operator_out138_out1            : std_logic;
  SIGNAL Logical_Operator_out139_out1            : std_logic;
  SIGNAL Logical_Operator_out140_out1            : std_logic;
  SIGNAL Logical_Operator_out141_out1            : std_logic;
  SIGNAL Logical_Operator_out142_out1            : std_logic;
  SIGNAL Logical_Operator_out143_out1            : std_logic;
  SIGNAL Logical_Operator_out144_out1            : std_logic;
  SIGNAL Logical_Operator_out145_out1            : std_logic;
  SIGNAL Logical_Operator_out146_out1            : std_logic;
  SIGNAL Logical_Operator_out147_out1            : std_logic;
  SIGNAL Logical_Operator_out148_out1            : std_logic;
  SIGNAL Logical_Operator_out149_out1            : std_logic;
  SIGNAL Logical_Operator_out150_out1            : std_logic;
  SIGNAL Logical_Operator_out151_out1            : std_logic;
  SIGNAL Logical_Operator_out152_out1            : std_logic;
  SIGNAL Logical_Operator_out153_out1            : std_logic;
  SIGNAL Logical_Operator_out154_out1            : std_logic;
  SIGNAL Logical_Operator_out155_out1            : std_logic;
  SIGNAL Logical_Operator_out156_out1            : std_logic;
  SIGNAL Logical_Operator_out157_out1            : std_logic;
  SIGNAL Logical_Operator_out158_out1            : std_logic;
  SIGNAL Logical_Operator_out159_out1            : std_logic;
  SIGNAL Logical_Operator_out160_out1            : std_logic;
  SIGNAL Logical_Operator_out161_out1            : std_logic;
  SIGNAL Logical_Operator_out162_out1            : std_logic;
  SIGNAL Logical_Operator_out163_out1            : std_logic;
  SIGNAL Logical_Operator_out164_out1            : std_logic;
  SIGNAL Logical_Operator_out165_out1            : std_logic;
  SIGNAL Logical_Operator_out166_out1            : std_logic;
  SIGNAL Logical_Operator_out167_out1            : std_logic;
  SIGNAL Logical_Operator_out168_out1            : std_logic;
  SIGNAL Logical_Operator_out169_out1            : std_logic;
  SIGNAL Logical_Operator_out170_out1            : std_logic;
  SIGNAL Logical_Operator_out171_out1            : std_logic;
  SIGNAL Logical_Operator_out172_out1            : std_logic;
  SIGNAL Logical_Operator_out173_out1            : std_logic;
  SIGNAL Logical_Operator_out174_out1            : std_logic;
  SIGNAL Logical_Operator_out175_out1            : std_logic;
  SIGNAL Logical_Operator_out176_out1            : std_logic;
  SIGNAL Logical_Operator_out177_out1            : std_logic;
  SIGNAL Logical_Operator_out178_out1            : std_logic;
  SIGNAL Logical_Operator_out179_out1            : std_logic;
  SIGNAL Logical_Operator_out180_out1            : std_logic;
  SIGNAL Logical_Operator_out181_out1            : std_logic;
  SIGNAL Logical_Operator_out182_out1            : std_logic;
  SIGNAL Logical_Operator_out183_out1            : std_logic;
  SIGNAL Logical_Operator_out184_out1            : std_logic;
  SIGNAL Logical_Operator_out185_out1            : std_logic;
  SIGNAL Logical_Operator_out186_out1            : std_logic;
  SIGNAL Logical_Operator_out187_out1            : std_logic;
  SIGNAL Logical_Operator_out188_out1            : std_logic;
  SIGNAL Logical_Operator_out189_out1            : std_logic;
  SIGNAL Logical_Operator_out190_out1            : std_logic;
  SIGNAL Logical_Operator_out191_out1            : std_logic;
  SIGNAL Logical_Operator_out192_out1            : std_logic;
  SIGNAL Logical_Operator_out193_out1            : std_logic;
  SIGNAL Logical_Operator_out194_out1            : std_logic;
  SIGNAL Logical_Operator_out195_out1            : std_logic;
  SIGNAL Logical_Operator_out196_out1            : std_logic;
  SIGNAL Logical_Operator_out197_out1            : std_logic;
  SIGNAL Logical_Operator_out198_out1            : std_logic;
  SIGNAL Logical_Operator_out199_out1            : std_logic;
  SIGNAL Logical_Operator_out200_out1            : std_logic;
  SIGNAL Logical_Operator_out201_out1            : std_logic;
  SIGNAL Logical_Operator_out202_out1            : std_logic;
  SIGNAL Logical_Operator_out203_out1            : std_logic;
  SIGNAL Logical_Operator_out204_out1            : std_logic;
  SIGNAL Logical_Operator_out205_out1            : std_logic;
  SIGNAL Logical_Operator_out206_out1            : std_logic;
  SIGNAL Logical_Operator_out207_out1            : std_logic;
  SIGNAL Logical_Operator_out208_out1            : std_logic;
  SIGNAL Logical_Operator_out209_out1            : std_logic;
  SIGNAL Logical_Operator_out210_out1            : std_logic;
  SIGNAL Logical_Operator_out211_out1            : std_logic;
  SIGNAL Logical_Operator_out212_out1            : std_logic;
  SIGNAL Logical_Operator_out213_out1            : std_logic;
  SIGNAL Logical_Operator_out214_out1            : std_logic;
  SIGNAL Logical_Operator_out215_out1            : std_logic;
  SIGNAL Logical_Operator_out216_out1            : std_logic;
  SIGNAL Logical_Operator_out217_out1            : std_logic;
  SIGNAL Logical_Operator_out218_out1            : std_logic;
  SIGNAL Logical_Operator_out219_out1            : std_logic;
  SIGNAL Logical_Operator_out220_out1            : std_logic;
  SIGNAL Logical_Operator_out221_out1            : std_logic;
  SIGNAL Logical_Operator_out222_out1            : std_logic;
  SIGNAL Logical_Operator_out223_out1            : std_logic;
  SIGNAL Logical_Operator_out224_out1            : std_logic;
  SIGNAL Logical_Operator_out225_out1            : std_logic;
  SIGNAL Logical_Operator_out226_out1            : std_logic;
  SIGNAL Logical_Operator_out227_out1            : std_logic;
  SIGNAL Logical_Operator_out228_out1            : std_logic;
  SIGNAL Logical_Operator_out229_out1            : std_logic;
  SIGNAL Logical_Operator_out230_out1            : std_logic;
  SIGNAL Logical_Operator_out231_out1            : std_logic;
  SIGNAL Logical_Operator_out232_out1            : std_logic;
  SIGNAL Logical_Operator_out233_out1            : std_logic;
  SIGNAL Logical_Operator_out234_out1            : std_logic;
  SIGNAL Logical_Operator_out235_out1            : std_logic;
  SIGNAL Logical_Operator_out236_out1            : std_logic;
  SIGNAL Logical_Operator_out237_out1            : std_logic;
  SIGNAL Logical_Operator_out238_out1            : std_logic;
  SIGNAL Logical_Operator_out239_out1            : std_logic;
  SIGNAL Logical_Operator_out240_out1            : std_logic;
  SIGNAL Logical_Operator_out241_out1            : std_logic;
  SIGNAL Logical_Operator_out242_out1            : std_logic;
  SIGNAL Logical_Operator_out243_out1            : std_logic;
  SIGNAL Logical_Operator_out244_out1            : std_logic;
  SIGNAL Logical_Operator_out245_out1            : std_logic;
  SIGNAL Logical_Operator_out246_out1            : std_logic;
  SIGNAL Logical_Operator_out247_out1            : std_logic;
  SIGNAL Logical_Operator_out248_out1            : std_logic;
  SIGNAL Logical_Operator_out249_out1            : std_logic;
  SIGNAL Logical_Operator_out250_out1            : std_logic;
  SIGNAL Logical_Operator_out251_out1            : std_logic;
  SIGNAL Logical_Operator_out252_out1            : std_logic;
  SIGNAL Logical_Operator_out253_out1            : std_logic;
  SIGNAL Logical_Operator_out254_out1            : std_logic;
  SIGNAL Logical_Operator_out255_out1            : std_logic;
  SIGNAL Logical_Operator_out256_out1            : std_logic;
  SIGNAL Logical_Operator_out257_out1            : std_logic;
  SIGNAL Logical_Operator_out258_out1            : std_logic;
  SIGNAL Logical_Operator_out259_out1            : std_logic;
  SIGNAL Logical_Operator_out260_out1            : std_logic;
  SIGNAL Logical_Operator_out261_out1            : std_logic;
  SIGNAL Logical_Operator_out262_out1            : std_logic;
  SIGNAL Logical_Operator_out263_out1            : std_logic;
  SIGNAL Logical_Operator_out264_out1            : std_logic;
  SIGNAL Logical_Operator_out265_out1            : std_logic;
  SIGNAL Logical_Operator_out266_out1            : std_logic;
  SIGNAL Logical_Operator_out267_out1            : std_logic;
  SIGNAL Logical_Operator_out268_out1            : std_logic;
  SIGNAL Logical_Operator_out269_out1            : std_logic;
  SIGNAL Logical_Operator_out270_out1            : std_logic;
  SIGNAL Logical_Operator_out271_out1            : std_logic;
  SIGNAL Logical_Operator_out272_out1            : std_logic;
  SIGNAL Logical_Operator_out273_out1            : std_logic;
  SIGNAL Logical_Operator_out274_out1            : std_logic;
  SIGNAL Logical_Operator_out275_out1            : std_logic;
  SIGNAL Logical_Operator_out276_out1            : std_logic;
  SIGNAL Logical_Operator_out277_out1            : std_logic;
  SIGNAL Logical_Operator_out278_out1            : std_logic;
  SIGNAL Logical_Operator_out279_out1            : std_logic;
  SIGNAL Logical_Operator_out280_out1            : std_logic;
  SIGNAL Logical_Operator_out281_out1            : std_logic;
  SIGNAL Logical_Operator_out282_out1            : std_logic;
  SIGNAL Logical_Operator_out283_out1            : std_logic;
  SIGNAL Logical_Operator_out284_out1            : std_logic;
  SIGNAL Logical_Operator_out285_out1            : std_logic;
  SIGNAL Logical_Operator_out286_out1            : std_logic;
  SIGNAL Logical_Operator_out287_out1            : std_logic;
  SIGNAL Logical_Operator_out288_out1            : std_logic;
  SIGNAL Logical_Operator_out289_out1            : std_logic;
  SIGNAL Logical_Operator_out290_out1            : std_logic;
  SIGNAL Logical_Operator_out291_out1            : std_logic;
  SIGNAL Logical_Operator_out292_out1            : std_logic;
  SIGNAL Logical_Operator_out293_out1            : std_logic;
  SIGNAL Logical_Operator_out294_out1            : std_logic;
  SIGNAL Logical_Operator_out295_out1            : std_logic;
  SIGNAL Logical_Operator_out296_out1            : std_logic;
  SIGNAL Logical_Operator_out297_out1            : std_logic;
  SIGNAL Logical_Operator_out298_out1            : std_logic;
  SIGNAL Logical_Operator_out299_out1            : std_logic;
  SIGNAL Logical_Operator_out300_out1            : std_logic;
  SIGNAL Logical_Operator_out301_out1            : std_logic;
  SIGNAL Logical_Operator_out302_out1            : std_logic;
  SIGNAL Logical_Operator_out303_out1            : std_logic;
  SIGNAL Logical_Operator_out304_out1            : std_logic;
  SIGNAL Logical_Operator_out305_out1            : std_logic;
  SIGNAL Logical_Operator_out306_out1            : std_logic;
  SIGNAL Logical_Operator_out307_out1            : std_logic;
  SIGNAL Logical_Operator_out308_out1            : std_logic;
  SIGNAL Logical_Operator_out309_out1            : std_logic;
  SIGNAL Logical_Operator_out310_out1            : std_logic;
  SIGNAL Logical_Operator_out311_out1            : std_logic;
  SIGNAL Logical_Operator_out312_out1            : std_logic;
  SIGNAL Logical_Operator_out313_out1            : std_logic;
  SIGNAL Logical_Operator_out314_out1            : std_logic;
  SIGNAL Logical_Operator_out315_out1            : std_logic;
  SIGNAL Logical_Operator_out316_out1            : std_logic;
  SIGNAL Logical_Operator_out317_out1            : std_logic;
  SIGNAL Logical_Operator_out318_out1            : std_logic;
  SIGNAL Logical_Operator_out319_out1            : std_logic;
  SIGNAL Logical_Operator_out320_out1            : std_logic;
  SIGNAL Logical_Operator_out321_out1            : std_logic;
  SIGNAL Logical_Operator_out322_out1            : std_logic;
  SIGNAL Logical_Operator_out323_out1            : std_logic;
  SIGNAL Logical_Operator_out324_out1            : std_logic;
  SIGNAL Logical_Operator_out325_out1            : std_logic;
  SIGNAL Logical_Operator_out326_out1            : std_logic;
  SIGNAL Logical_Operator_out327_out1            : std_logic;
  SIGNAL Logical_Operator_out328_out1            : std_logic;
  SIGNAL Logical_Operator_out329_out1            : std_logic;
  SIGNAL Logical_Operator_out330_out1            : std_logic;
  SIGNAL Logical_Operator_out331_out1            : std_logic;
  SIGNAL Logical_Operator_out332_out1            : std_logic;
  SIGNAL Logical_Operator_out333_out1            : std_logic;
  SIGNAL Logical_Operator_out334_out1            : std_logic;
  SIGNAL Logical_Operator_out335_out1            : std_logic;
  SIGNAL Logical_Operator_out336_out1            : std_logic;
  SIGNAL Logical_Operator_out337_out1            : std_logic;
  SIGNAL Logical_Operator_out338_out1            : std_logic;
  SIGNAL Logical_Operator_out339_out1            : std_logic;
  SIGNAL Logical_Operator_out340_out1            : std_logic;
  SIGNAL Logical_Operator_out341_out1            : std_logic;
  SIGNAL Logical_Operator_out342_out1            : std_logic;
  SIGNAL Logical_Operator_out343_out1            : std_logic;
  SIGNAL Logical_Operator_out344_out1            : std_logic;
  SIGNAL Logical_Operator_out345_out1            : std_logic;
  SIGNAL Logical_Operator_out346_out1            : std_logic;
  SIGNAL Logical_Operator_out347_out1            : std_logic;
  SIGNAL Logical_Operator_out348_out1            : std_logic;
  SIGNAL Logical_Operator_out349_out1            : std_logic;
  SIGNAL Logical_Operator_out350_out1            : std_logic;
  SIGNAL Logical_Operator_out351_out1            : std_logic;
  SIGNAL Logical_Operator_out352_out1            : std_logic;
  SIGNAL Logical_Operator_out353_out1            : std_logic;
  SIGNAL Logical_Operator_out354_out1            : std_logic;
  SIGNAL Logical_Operator_out355_out1            : std_logic;
  SIGNAL Logical_Operator_out356_out1            : std_logic;
  SIGNAL Logical_Operator_out357_out1            : std_logic;
  SIGNAL Logical_Operator_out358_out1            : std_logic;
  SIGNAL Logical_Operator_out359_out1            : std_logic;
  SIGNAL Logical_Operator_out360_out1            : std_logic;
  SIGNAL Logical_Operator_out361_out1            : std_logic;
  SIGNAL Logical_Operator_out362_out1            : std_logic;
  SIGNAL Logical_Operator_out363_out1            : std_logic;
  SIGNAL Logical_Operator_out364_out1            : std_logic;
  SIGNAL Logical_Operator_out365_out1            : std_logic;
  SIGNAL Logical_Operator_out366_out1            : std_logic;
  SIGNAL Logical_Operator_out367_out1            : std_logic;
  SIGNAL Logical_Operator_out368_out1            : std_logic;
  SIGNAL Logical_Operator_out369_out1            : std_logic;
  SIGNAL Logical_Operator_out370_out1            : std_logic;
  SIGNAL Logical_Operator_out371_out1            : std_logic;
  SIGNAL Logical_Operator_out372_out1            : std_logic;
  SIGNAL Logical_Operator_out373_out1            : std_logic;
  SIGNAL Logical_Operator_out374_out1            : std_logic;
  SIGNAL Logical_Operator_out375_out1            : std_logic;
  SIGNAL Logical_Operator_out376_out1            : std_logic;
  SIGNAL Logical_Operator_out377_out1            : std_logic;
  SIGNAL Logical_Operator_out378_out1            : std_logic;
  SIGNAL Logical_Operator_out379_out1            : std_logic;
  SIGNAL Logical_Operator_out380_out1            : std_logic;
  SIGNAL Logical_Operator_out381_out1            : std_logic;
  SIGNAL Logical_Operator_out382_out1            : std_logic;
  SIGNAL Logical_Operator_out383_out1            : std_logic;
  SIGNAL Logical_Operator_out384_out1            : std_logic;
  SIGNAL Logical_Operator_out385_out1            : std_logic;
  SIGNAL Logical_Operator_out386_out1            : std_logic;
  SIGNAL Logical_Operator_out387_out1            : std_logic;
  SIGNAL Logical_Operator_out388_out1            : std_logic;
  SIGNAL Logical_Operator_out389_out1            : std_logic;
  SIGNAL Logical_Operator_out390_out1            : std_logic;
  SIGNAL Logical_Operator_out391_out1            : std_logic;
  SIGNAL Logical_Operator_out392_out1            : std_logic;
  SIGNAL Logical_Operator_out393_out1            : std_logic;
  SIGNAL Logical_Operator_out394_out1            : std_logic;
  SIGNAL Logical_Operator_out395_out1            : std_logic;
  SIGNAL Logical_Operator_out396_out1            : std_logic;
  SIGNAL Logical_Operator_out397_out1            : std_logic;
  SIGNAL Logical_Operator_out398_out1            : std_logic;
  SIGNAL Logical_Operator_out399_out1            : std_logic;
  SIGNAL Logical_Operator_out400_out1            : std_logic;
  SIGNAL Logical_Operator_out401_out1            : std_logic;
  SIGNAL Logical_Operator_out402_out1            : std_logic;
  SIGNAL Logical_Operator_out403_out1            : std_logic;
  SIGNAL Logical_Operator_out404_out1            : std_logic;
  SIGNAL Logical_Operator_out405_out1            : std_logic;
  SIGNAL Logical_Operator_out406_out1            : std_logic;
  SIGNAL Logical_Operator_out407_out1            : std_logic;
  SIGNAL Logical_Operator_out408_out1            : std_logic;
  SIGNAL Logical_Operator_out409_out1            : std_logic;
  SIGNAL Logical_Operator_out410_out1            : std_logic;
  SIGNAL Logical_Operator_out411_out1            : std_logic;
  SIGNAL Logical_Operator_out412_out1            : std_logic;
  SIGNAL Logical_Operator_out413_out1            : std_logic;
  SIGNAL Logical_Operator_out414_out1            : std_logic;
  SIGNAL Logical_Operator_out415_out1            : std_logic;
  SIGNAL Logical_Operator_out416_out1            : std_logic;
  SIGNAL Logical_Operator_out417_out1            : std_logic;
  SIGNAL Logical_Operator_out418_out1            : std_logic;
  SIGNAL Logical_Operator_out419_out1            : std_logic;
  SIGNAL Logical_Operator_out420_out1            : std_logic;
  SIGNAL Logical_Operator_out421_out1            : std_logic;
  SIGNAL Logical_Operator_out422_out1            : std_logic;
  SIGNAL Logical_Operator_out423_out1            : std_logic;
  SIGNAL Logical_Operator_out424_out1            : std_logic;
  SIGNAL Logical_Operator_out425_out1            : std_logic;
  SIGNAL Logical_Operator_out426_out1            : std_logic;
  SIGNAL Logical_Operator_out427_out1            : std_logic;
  SIGNAL Logical_Operator_out428_out1            : std_logic;
  SIGNAL Logical_Operator_out429_out1            : std_logic;
  SIGNAL Logical_Operator_out430_out1            : std_logic;
  SIGNAL Logical_Operator_out431_out1            : std_logic;
  SIGNAL Logical_Operator_out432_out1            : std_logic;
  SIGNAL Logical_Operator_out433_out1            : std_logic;
  SIGNAL Logical_Operator_out434_out1            : std_logic;
  SIGNAL Logical_Operator_out435_out1            : std_logic;
  SIGNAL Logical_Operator_out436_out1            : std_logic;
  SIGNAL Logical_Operator_out437_out1            : std_logic;
  SIGNAL Logical_Operator_out438_out1            : std_logic;
  SIGNAL Logical_Operator_out439_out1            : std_logic;
  SIGNAL Logical_Operator_out440_out1            : std_logic;
  SIGNAL Logical_Operator_out441_out1            : std_logic;
  SIGNAL Logical_Operator_out442_out1            : std_logic;
  SIGNAL Logical_Operator_out443_out1            : std_logic;
  SIGNAL Logical_Operator_out444_out1            : std_logic;
  SIGNAL Logical_Operator_out445_out1            : std_logic;
  SIGNAL Logical_Operator_out446_out1            : std_logic;
  SIGNAL Logical_Operator_out447_out1            : std_logic;
  SIGNAL Logical_Operator_out448_out1            : std_logic;
  SIGNAL Logical_Operator_out449_out1            : std_logic;
  SIGNAL Logical_Operator_out450_out1            : std_logic;
  SIGNAL Logical_Operator_out451_out1            : std_logic;
  SIGNAL Logical_Operator_out452_out1            : std_logic;
  SIGNAL Logical_Operator_out453_out1            : std_logic;
  SIGNAL Logical_Operator_out454_out1            : std_logic;
  SIGNAL Logical_Operator_out455_out1            : std_logic;
  SIGNAL Logical_Operator_out456_out1            : std_logic;
  SIGNAL Logical_Operator_out457_out1            : std_logic;
  SIGNAL Logical_Operator_out458_out1            : std_logic;
  SIGNAL Logical_Operator_out459_out1            : std_logic;
  SIGNAL Logical_Operator_out460_out1            : std_logic;
  SIGNAL Logical_Operator_out461_out1            : std_logic;
  SIGNAL Logical_Operator_out462_out1            : std_logic;
  SIGNAL Logical_Operator_out463_out1            : std_logic;
  SIGNAL Logical_Operator_out464_out1            : std_logic;
  SIGNAL Logical_Operator_out465_out1            : std_logic;
  SIGNAL Logical_Operator_out466_out1            : std_logic;
  SIGNAL Logical_Operator_out467_out1            : std_logic;
  SIGNAL Logical_Operator_out468_out1            : std_logic;
  SIGNAL Logical_Operator_out469_out1            : std_logic;
  SIGNAL Logical_Operator_out470_out1            : std_logic;
  SIGNAL Logical_Operator_out471_out1            : std_logic;
  SIGNAL Logical_Operator_out472_out1            : std_logic;
  SIGNAL Logical_Operator_out473_out1            : std_logic;
  SIGNAL Logical_Operator_out474_out1            : std_logic;
  SIGNAL Logical_Operator_out475_out1            : std_logic;
  SIGNAL Logical_Operator_out476_out1            : std_logic;
  SIGNAL Logical_Operator_out477_out1            : std_logic;
  SIGNAL Logical_Operator_out478_out1            : std_logic;
  SIGNAL Logical_Operator_out479_out1            : std_logic;
  SIGNAL Logical_Operator_out480_out1            : std_logic;
  SIGNAL Logical_Operator_out481_out1            : std_logic;
  SIGNAL Logical_Operator_out482_out1            : std_logic;
  SIGNAL Logical_Operator_out483_out1            : std_logic;
  SIGNAL Logical_Operator_out484_out1            : std_logic;
  SIGNAL Logical_Operator_out485_out1            : std_logic;
  SIGNAL Logical_Operator_out486_out1            : std_logic;
  SIGNAL Logical_Operator_out487_out1            : std_logic;
  SIGNAL Logical_Operator_out488_out1            : std_logic;
  SIGNAL Logical_Operator_out489_out1            : std_logic;
  SIGNAL Logical_Operator_out490_out1            : std_logic;
  SIGNAL Logical_Operator_out491_out1            : std_logic;
  SIGNAL Logical_Operator_out492_out1            : std_logic;
  SIGNAL Logical_Operator_out493_out1            : std_logic;
  SIGNAL Logical_Operator_out494_out1            : std_logic;
  SIGNAL Logical_Operator_out495_out1            : std_logic;
  SIGNAL Logical_Operator_out496_out1            : std_logic;
  SIGNAL Logical_Operator_out497_out1            : std_logic;
  SIGNAL Logical_Operator_out498_out1            : std_logic;
  SIGNAL Logical_Operator_out499_out1            : std_logic;
  SIGNAL Logical_Operator_out500_out1            : std_logic;
  SIGNAL Logical_Operator_out501_out1            : std_logic;
  SIGNAL Logical_Operator_out502_out1            : std_logic;
  SIGNAL Logical_Operator_out503_out1            : std_logic;
  SIGNAL Logical_Operator_out504_out1            : std_logic;
  SIGNAL Logical_Operator_out505_out1            : std_logic;
  SIGNAL Logical_Operator_out506_out1            : std_logic;
  SIGNAL Logical_Operator_out507_out1            : std_logic;
  SIGNAL Logical_Operator_out508_out1            : std_logic;
  SIGNAL Logical_Operator_out509_out1            : std_logic;
  SIGNAL Logical_Operator_out510_out1            : std_logic;
  SIGNAL Logical_Operator_out511_out1            : std_logic;
  SIGNAL Logical_Operator_out512_out1            : std_logic;
  SIGNAL Logical_Operator_out513_out1            : std_logic;
  SIGNAL Logical_Operator_out514_out1            : std_logic;
  SIGNAL Logical_Operator_out515_out1            : std_logic;
  SIGNAL Logical_Operator_out516_out1            : std_logic;
  SIGNAL Logical_Operator_out517_out1            : std_logic;
  SIGNAL Logical_Operator_out518_out1            : std_logic;
  SIGNAL Logical_Operator_out519_out1            : std_logic;
  SIGNAL Logical_Operator_out520_out1            : std_logic;
  SIGNAL Logical_Operator_out521_out1            : std_logic;
  SIGNAL Logical_Operator_out522_out1            : std_logic;
  SIGNAL Logical_Operator_out523_out1            : std_logic;
  SIGNAL Logical_Operator_out524_out1            : std_logic;
  SIGNAL Logical_Operator_out525_out1            : std_logic;
  SIGNAL Logical_Operator_out526_out1            : std_logic;
  SIGNAL Logical_Operator_out527_out1            : std_logic;
  SIGNAL Logical_Operator_out528_out1            : std_logic;
  SIGNAL Logical_Operator_out529_out1            : std_logic;
  SIGNAL Logical_Operator_out530_out1            : std_logic;
  SIGNAL Logical_Operator_out531_out1            : std_logic;
  SIGNAL Logical_Operator_out532_out1            : std_logic;
  SIGNAL Logical_Operator_out533_out1            : std_logic;
  SIGNAL Logical_Operator_out534_out1            : std_logic;
  SIGNAL Logical_Operator_out535_out1            : std_logic;
  SIGNAL Logical_Operator_out536_out1            : std_logic;
  SIGNAL Logical_Operator_out537_out1            : std_logic;
  SIGNAL Logical_Operator_out538_out1            : std_logic;
  SIGNAL Logical_Operator_out539_out1            : std_logic;
  SIGNAL Logical_Operator_out540_out1            : std_logic;
  SIGNAL Logical_Operator_out541_out1            : std_logic;
  SIGNAL Logical_Operator_out542_out1            : std_logic;
  SIGNAL Logical_Operator_out543_out1            : std_logic;
  SIGNAL Logical_Operator_out544_out1            : std_logic;
  SIGNAL Logical_Operator_out545_out1            : std_logic;
  SIGNAL Logical_Operator_out546_out1            : std_logic;
  SIGNAL Logical_Operator_out547_out1            : std_logic;
  SIGNAL Logical_Operator_out548_out1            : std_logic;
  SIGNAL Logical_Operator_out549_out1            : std_logic;
  SIGNAL Logical_Operator_out550_out1            : std_logic;
  SIGNAL Logical_Operator_out551_out1            : std_logic;
  SIGNAL Logical_Operator_out552_out1            : std_logic;
  SIGNAL Logical_Operator_out553_out1            : std_logic;
  SIGNAL Logical_Operator_out554_out1            : std_logic;
  SIGNAL Logical_Operator_out555_out1            : std_logic;
  SIGNAL Logical_Operator_out556_out1            : std_logic;
  SIGNAL Logical_Operator_out557_out1            : std_logic;
  SIGNAL Logical_Operator_out558_out1            : std_logic;
  SIGNAL Logical_Operator_out559_out1            : std_logic;
  SIGNAL Logical_Operator_out560_out1            : std_logic;
  SIGNAL Logical_Operator_out561_out1            : std_logic;
  SIGNAL Logical_Operator_out562_out1            : std_logic;
  SIGNAL Logical_Operator_out563_out1            : std_logic;
  SIGNAL Logical_Operator_out564_out1            : std_logic;
  SIGNAL Logical_Operator_out565_out1            : std_logic;
  SIGNAL Logical_Operator_out566_out1            : std_logic;
  SIGNAL Logical_Operator_out567_out1            : std_logic;
  SIGNAL Logical_Operator_out568_out1            : std_logic;
  SIGNAL Logical_Operator_out569_out1            : std_logic;
  SIGNAL Logical_Operator_out570_out1            : std_logic;
  SIGNAL Logical_Operator_out571_out1            : std_logic;
  SIGNAL Logical_Operator_out572_out1            : std_logic;
  SIGNAL Logical_Operator_out573_out1            : std_logic;
  SIGNAL Logical_Operator_out574_out1            : std_logic;
  SIGNAL Logical_Operator_out575_out1            : std_logic;
  SIGNAL Logical_Operator_out576_out1            : std_logic;
  SIGNAL Logical_Operator_out577_out1            : std_logic;
  SIGNAL Logical_Operator_out578_out1            : std_logic;
  SIGNAL Logical_Operator_out579_out1            : std_logic;
  SIGNAL Logical_Operator_out580_out1            : std_logic;
  SIGNAL Logical_Operator_out581_out1            : std_logic;
  SIGNAL Logical_Operator_out582_out1            : std_logic;
  SIGNAL Logical_Operator_out583_out1            : std_logic;
  SIGNAL Logical_Operator_out584_out1            : std_logic;
  SIGNAL Logical_Operator_out585_out1            : std_logic;
  SIGNAL Logical_Operator_out586_out1            : std_logic;
  SIGNAL Logical_Operator_out587_out1            : std_logic;
  SIGNAL Logical_Operator_out588_out1            : std_logic;
  SIGNAL Logical_Operator_out589_out1            : std_logic;
  SIGNAL Logical_Operator_out590_out1            : std_logic;
  SIGNAL Logical_Operator_out591_out1            : std_logic;
  SIGNAL Logical_Operator_out592_out1            : std_logic;
  SIGNAL Logical_Operator_out593_out1            : std_logic;
  SIGNAL Logical_Operator_out594_out1            : std_logic;
  SIGNAL Logical_Operator_out595_out1            : std_logic;
  SIGNAL Logical_Operator_out596_out1            : std_logic;
  SIGNAL Logical_Operator_out597_out1            : std_logic;
  SIGNAL Logical_Operator_out598_out1            : std_logic;
  SIGNAL Logical_Operator_out599_out1            : std_logic;
  SIGNAL Logical_Operator_out600_out1            : std_logic;
  SIGNAL Logical_Operator_out601_out1            : std_logic;
  SIGNAL Logical_Operator_out602_out1            : std_logic;
  SIGNAL Logical_Operator_out603_out1            : std_logic;
  SIGNAL Logical_Operator_out604_out1            : std_logic;
  SIGNAL Logical_Operator_out605_out1            : std_logic;
  SIGNAL Logical_Operator_out606_out1            : std_logic;
  SIGNAL Logical_Operator_out607_out1            : std_logic;
  SIGNAL Logical_Operator_out608_out1            : std_logic;
  SIGNAL Logical_Operator_out609_out1            : std_logic;
  SIGNAL Logical_Operator_out610_out1            : std_logic;
  SIGNAL Logical_Operator_out611_out1            : std_logic;
  SIGNAL Logical_Operator_out612_out1            : std_logic;
  SIGNAL Logical_Operator_out613_out1            : std_logic;
  SIGNAL Logical_Operator_out614_out1            : std_logic;
  SIGNAL Logical_Operator_out615_out1            : std_logic;
  SIGNAL Logical_Operator_out616_out1            : std_logic;
  SIGNAL Logical_Operator_out617_out1            : std_logic;
  SIGNAL Logical_Operator_out618_out1            : std_logic;
  SIGNAL Logical_Operator_out619_out1            : std_logic;
  SIGNAL Logical_Operator_out620_out1            : std_logic;
  SIGNAL Logical_Operator_out621_out1            : std_logic;
  SIGNAL Logical_Operator_out622_out1            : std_logic;
  SIGNAL Logical_Operator_out623_out1            : std_logic;
  SIGNAL Logical_Operator_out624_out1            : std_logic;
  SIGNAL Logical_Operator_out625_out1            : std_logic;
  SIGNAL Logical_Operator_out626_out1            : std_logic;
  SIGNAL Logical_Operator_out627_out1            : std_logic;
  SIGNAL Logical_Operator_out628_out1            : std_logic;
  SIGNAL Logical_Operator_out629_out1            : std_logic;
  SIGNAL Logical_Operator_out630_out1            : std_logic;
  SIGNAL Logical_Operator_out631_out1            : std_logic;
  SIGNAL Logical_Operator_out632_out1            : std_logic;
  SIGNAL Logical_Operator_out633_out1            : std_logic;
  SIGNAL Logical_Operator_out634_out1            : std_logic;
  SIGNAL Logical_Operator_out635_out1            : std_logic;
  SIGNAL Logical_Operator_out636_out1            : std_logic;
  SIGNAL Logical_Operator_out637_out1            : std_logic;
  SIGNAL Logical_Operator_out638_out1            : std_logic;
  SIGNAL Logical_Operator_out639_out1            : std_logic;
  SIGNAL Logical_Operator_out640_out1            : std_logic;
  SIGNAL Logical_Operator_out641_out1            : std_logic;
  SIGNAL Logical_Operator_out642_out1            : std_logic;
  SIGNAL Logical_Operator_out643_out1            : std_logic;
  SIGNAL Logical_Operator_out644_out1            : std_logic;
  SIGNAL Logical_Operator_out645_out1            : std_logic;
  SIGNAL Logical_Operator_out646_out1            : std_logic;
  SIGNAL Logical_Operator_out647_out1            : std_logic;
  SIGNAL Logical_Operator_out648_out1            : std_logic;
  SIGNAL Logical_Operator_out649_out1            : std_logic;
  SIGNAL Logical_Operator_out650_out1            : std_logic;
  SIGNAL Logical_Operator_out651_out1            : std_logic;
  SIGNAL Logical_Operator_out652_out1            : std_logic;
  SIGNAL Logical_Operator_out653_out1            : std_logic;
  SIGNAL Logical_Operator_out654_out1            : std_logic;
  SIGNAL Logical_Operator_out655_out1            : std_logic;
  SIGNAL Logical_Operator_out656_out1            : std_logic;
  SIGNAL Logical_Operator_out657_out1            : std_logic;
  SIGNAL Logical_Operator_out658_out1            : std_logic;
  SIGNAL Logical_Operator_out659_out1            : std_logic;
  SIGNAL Logical_Operator_out660_out1            : std_logic;
  SIGNAL Logical_Operator_out661_out1            : std_logic;
  SIGNAL Logical_Operator_out662_out1            : std_logic;
  SIGNAL Logical_Operator_out663_out1            : std_logic;
  SIGNAL Logical_Operator_out664_out1            : std_logic;
  SIGNAL Logical_Operator_out665_out1            : std_logic;
  SIGNAL Logical_Operator_out666_out1            : std_logic;
  SIGNAL Logical_Operator_out667_out1            : std_logic;
  SIGNAL Logical_Operator_out668_out1            : std_logic;
  SIGNAL Logical_Operator_out669_out1            : std_logic;
  SIGNAL Logical_Operator_out670_out1            : std_logic;
  SIGNAL Logical_Operator_out671_out1            : std_logic;
  SIGNAL Logical_Operator_out672_out1            : std_logic;
  SIGNAL Logical_Operator_out673_out1            : std_logic;
  SIGNAL Logical_Operator_out674_out1            : std_logic;
  SIGNAL Logical_Operator_out675_out1            : std_logic;
  SIGNAL Logical_Operator_out676_out1            : std_logic;
  SIGNAL Logical_Operator_out677_out1            : std_logic;
  SIGNAL Logical_Operator_out678_out1            : std_logic;
  SIGNAL Logical_Operator_out679_out1            : std_logic;
  SIGNAL Logical_Operator_out680_out1            : std_logic;
  SIGNAL Logical_Operator_out681_out1            : std_logic;
  SIGNAL Logical_Operator_out682_out1            : std_logic;
  SIGNAL Logical_Operator_out683_out1            : std_logic;
  SIGNAL Logical_Operator_out684_out1            : std_logic;
  SIGNAL Logical_Operator_out685_out1            : std_logic;
  SIGNAL Logical_Operator_out686_out1            : std_logic;
  SIGNAL Logical_Operator_out687_out1            : std_logic;
  SIGNAL Logical_Operator_out688_out1            : std_logic;
  SIGNAL Logical_Operator_out689_out1            : std_logic;
  SIGNAL Logical_Operator_out690_out1            : std_logic;
  SIGNAL Logical_Operator_out691_out1            : std_logic;
  SIGNAL Logical_Operator_out692_out1            : std_logic;
  SIGNAL Logical_Operator_out693_out1            : std_logic;
  SIGNAL Logical_Operator_out694_out1            : std_logic;
  SIGNAL Logical_Operator_out695_out1            : std_logic;
  SIGNAL Logical_Operator_out696_out1            : std_logic;
  SIGNAL Logical_Operator_out697_out1            : std_logic;
  SIGNAL Logical_Operator_out698_out1            : std_logic;
  SIGNAL Logical_Operator_out699_out1            : std_logic;
  SIGNAL Logical_Operator_out700_out1            : std_logic;
  SIGNAL Logical_Operator_out701_out1            : std_logic;
  SIGNAL Logical_Operator_out702_out1            : std_logic;
  SIGNAL Logical_Operator_out703_out1            : std_logic;
  SIGNAL Logical_Operator_out704_out1            : std_logic;
  SIGNAL Logical_Operator_out705_out1            : std_logic;
  SIGNAL Logical_Operator_out706_out1            : std_logic;
  SIGNAL Logical_Operator_out707_out1            : std_logic;
  SIGNAL Logical_Operator_out708_out1            : std_logic;
  SIGNAL Logical_Operator_out709_out1            : std_logic;
  SIGNAL Logical_Operator_out710_out1            : std_logic;
  SIGNAL Logical_Operator_out711_out1            : std_logic;
  SIGNAL Logical_Operator_out712_out1            : std_logic;
  SIGNAL Logical_Operator_out713_out1            : std_logic;
  SIGNAL Logical_Operator_out714_out1            : std_logic;
  SIGNAL Logical_Operator_out715_out1            : std_logic;
  SIGNAL Logical_Operator_out716_out1            : std_logic;
  SIGNAL Logical_Operator_out717_out1            : std_logic;
  SIGNAL Logical_Operator_out718_out1            : std_logic;
  SIGNAL Logical_Operator_out719_out1            : std_logic;
  SIGNAL Logical_Operator_out720_out1            : std_logic;
  SIGNAL Logical_Operator_out721_out1            : std_logic;
  SIGNAL Logical_Operator_out722_out1            : std_logic;
  SIGNAL Logical_Operator_out723_out1            : std_logic;
  SIGNAL Logical_Operator_out724_out1            : std_logic;
  SIGNAL Logical_Operator_out725_out1            : std_logic;
  SIGNAL Logical_Operator_out726_out1            : std_logic;
  SIGNAL Logical_Operator_out727_out1            : std_logic;
  SIGNAL Logical_Operator_out728_out1            : std_logic;
  SIGNAL Logical_Operator_out729_out1            : std_logic;
  SIGNAL Logical_Operator_out730_out1            : std_logic;
  SIGNAL Logical_Operator_out731_out1            : std_logic;
  SIGNAL Logical_Operator_out732_out1            : std_logic;
  SIGNAL Logical_Operator_out733_out1            : std_logic;
  SIGNAL Logical_Operator_out734_out1            : std_logic;
  SIGNAL Logical_Operator_out735_out1            : std_logic;
  SIGNAL Logical_Operator_out736_out1            : std_logic;
  SIGNAL Logical_Operator_out737_out1            : std_logic;
  SIGNAL Logical_Operator_out738_out1            : std_logic;
  SIGNAL Logical_Operator_out739_out1            : std_logic;
  SIGNAL Logical_Operator_out740_out1            : std_logic;
  SIGNAL Logical_Operator_out741_out1            : std_logic;
  SIGNAL Logical_Operator_out742_out1            : std_logic;
  SIGNAL Logical_Operator_out743_out1            : std_logic;
  SIGNAL Logical_Operator_out744_out1            : std_logic;
  SIGNAL Logical_Operator_out745_out1            : std_logic;
  SIGNAL Logical_Operator_out746_out1            : std_logic;
  SIGNAL Logical_Operator_out747_out1            : std_logic;
  SIGNAL Logical_Operator_out748_out1            : std_logic;
  SIGNAL Logical_Operator_out749_out1            : std_logic;
  SIGNAL Logical_Operator_out750_out1            : std_logic;
  SIGNAL Logical_Operator_out751_out1            : std_logic;
  SIGNAL Logical_Operator_out752_out1            : std_logic;
  SIGNAL Logical_Operator_out753_out1            : std_logic;
  SIGNAL Logical_Operator_out754_out1            : std_logic;
  SIGNAL Logical_Operator_out755_out1            : std_logic;
  SIGNAL Logical_Operator_out756_out1            : std_logic;
  SIGNAL Logical_Operator_out757_out1            : std_logic;
  SIGNAL Logical_Operator_out758_out1            : std_logic;
  SIGNAL Logical_Operator_out759_out1            : std_logic;
  SIGNAL Logical_Operator_out760_out1            : std_logic;
  SIGNAL Logical_Operator_out761_out1            : std_logic;
  SIGNAL Logical_Operator_out762_out1            : std_logic;
  SIGNAL Logical_Operator_out763_out1            : std_logic;
  SIGNAL Logical_Operator_out764_out1            : std_logic;
  SIGNAL Logical_Operator_out765_out1            : std_logic;
  SIGNAL Logical_Operator_out766_out1            : std_logic;
  SIGNAL Logical_Operator_out767_out1            : std_logic;
  SIGNAL Logical_Operator_out768_out1            : std_logic;
  SIGNAL Logical_Operator_out769_out1            : std_logic;
  SIGNAL Logical_Operator_out770_out1            : std_logic;
  SIGNAL Logical_Operator_out771_out1            : std_logic;
  SIGNAL Logical_Operator_out772_out1            : std_logic;
  SIGNAL Logical_Operator_out773_out1            : std_logic;
  SIGNAL Logical_Operator_out774_out1            : std_logic;
  SIGNAL Logical_Operator_out775_out1            : std_logic;
  SIGNAL Logical_Operator_out776_out1            : std_logic;
  SIGNAL Logical_Operator_out777_out1            : std_logic;
  SIGNAL Logical_Operator_out778_out1            : std_logic;
  SIGNAL Logical_Operator_out779_out1            : std_logic;
  SIGNAL Logical_Operator_out780_out1            : std_logic;
  SIGNAL Logical_Operator_out781_out1            : std_logic;
  SIGNAL Logical_Operator_out782_out1            : std_logic;
  SIGNAL Logical_Operator_out783_out1            : std_logic;
  SIGNAL Logical_Operator_out784_out1            : std_logic;
  SIGNAL Logical_Operator_out785_out1            : std_logic;
  SIGNAL Logical_Operator_out786_out1            : std_logic;
  SIGNAL Logical_Operator_out787_out1            : std_logic;
  SIGNAL Logical_Operator_out788_out1            : std_logic;
  SIGNAL Logical_Operator_out789_out1            : std_logic;
  SIGNAL Logical_Operator_out790_out1            : std_logic;
  SIGNAL Logical_Operator_out791_out1            : std_logic;
  SIGNAL Logical_Operator_out792_out1            : std_logic;
  SIGNAL Logical_Operator_out793_out1            : std_logic;
  SIGNAL Logical_Operator_out794_out1            : std_logic;
  SIGNAL Logical_Operator_out795_out1            : std_logic;
  SIGNAL Logical_Operator_out796_out1            : std_logic;
  SIGNAL Logical_Operator_out797_out1            : std_logic;
  SIGNAL Logical_Operator_out798_out1            : std_logic;
  SIGNAL Logical_Operator_out799_out1            : std_logic;
  SIGNAL Logical_Operator_out800_out1            : std_logic;
  SIGNAL Logical_Operator_out801_out1            : std_logic;
  SIGNAL Logical_Operator_out802_out1            : std_logic;
  SIGNAL Logical_Operator_out803_out1            : std_logic;
  SIGNAL Logical_Operator_out804_out1            : std_logic;
  SIGNAL Logical_Operator_out805_out1            : std_logic;
  SIGNAL Logical_Operator_out806_out1            : std_logic;
  SIGNAL Logical_Operator_out807_out1            : std_logic;
  SIGNAL Logical_Operator_out808_out1            : std_logic;
  SIGNAL Logical_Operator_out809_out1            : std_logic;
  SIGNAL Logical_Operator_out810_out1            : std_logic;
  SIGNAL Logical_Operator_out811_out1            : std_logic;
  SIGNAL Logical_Operator_out812_out1            : std_logic;
  SIGNAL Logical_Operator_out813_out1            : std_logic;
  SIGNAL Logical_Operator_out814_out1            : std_logic;
  SIGNAL Logical_Operator_out815_out1            : std_logic;
  SIGNAL Logical_Operator_out816_out1            : std_logic;
  SIGNAL Logical_Operator_out817_out1            : std_logic;
  SIGNAL Logical_Operator_out818_out1            : std_logic;
  SIGNAL Logical_Operator_out819_out1            : std_logic;
  SIGNAL Logical_Operator_out820_out1            : std_logic;
  SIGNAL Logical_Operator_out821_out1            : std_logic;
  SIGNAL Logical_Operator_out822_out1            : std_logic;
  SIGNAL Logical_Operator_out823_out1            : std_logic;
  SIGNAL Logical_Operator_out824_out1            : std_logic;
  SIGNAL Logical_Operator_out825_out1            : std_logic;
  SIGNAL Logical_Operator_out826_out1            : std_logic;
  SIGNAL Logical_Operator_out827_out1            : std_logic;
  SIGNAL Logical_Operator_out828_out1            : std_logic;
  SIGNAL Logical_Operator_out829_out1            : std_logic;
  SIGNAL Logical_Operator_out830_out1            : std_logic;
  SIGNAL Logical_Operator_out831_out1            : std_logic;
  SIGNAL Logical_Operator_out832_out1            : std_logic;
  SIGNAL Logical_Operator_out833_out1            : std_logic;
  SIGNAL Logical_Operator_out834_out1            : std_logic;
  SIGNAL Logical_Operator_out835_out1            : std_logic;
  SIGNAL Logical_Operator_out836_out1            : std_logic;
  SIGNAL Logical_Operator_out837_out1            : std_logic;
  SIGNAL Logical_Operator_out838_out1            : std_logic;
  SIGNAL Logical_Operator_out839_out1            : std_logic;
  SIGNAL Logical_Operator_out840_out1            : std_logic;
  SIGNAL Logical_Operator_out841_out1            : std_logic;
  SIGNAL Logical_Operator_out842_out1            : std_logic;
  SIGNAL Logical_Operator_out843_out1            : std_logic;
  SIGNAL Logical_Operator_out844_out1            : std_logic;
  SIGNAL Logical_Operator_out845_out1            : std_logic;
  SIGNAL Logical_Operator_out846_out1            : std_logic;
  SIGNAL Logical_Operator_out847_out1            : std_logic;
  SIGNAL Logical_Operator_out848_out1            : std_logic;
  SIGNAL Logical_Operator_out849_out1            : std_logic;
  SIGNAL Logical_Operator_out850_out1            : std_logic;
  SIGNAL Logical_Operator_out851_out1            : std_logic;
  SIGNAL Logical_Operator_out852_out1            : std_logic;
  SIGNAL Logical_Operator_out853_out1            : std_logic;
  SIGNAL Logical_Operator_out854_out1            : std_logic;
  SIGNAL Logical_Operator_out855_out1            : std_logic;
  SIGNAL Logical_Operator_out856_out1            : std_logic;
  SIGNAL Logical_Operator_out857_out1            : std_logic;
  SIGNAL Logical_Operator_out858_out1            : std_logic;
  SIGNAL Logical_Operator_out859_out1            : std_logic;
  SIGNAL Logical_Operator_out860_out1            : std_logic;
  SIGNAL Logical_Operator_out861_out1            : std_logic;
  SIGNAL Logical_Operator_out862_out1            : std_logic;
  SIGNAL Logical_Operator_out863_out1            : std_logic;
  SIGNAL Logical_Operator_out864_out1            : std_logic;
  SIGNAL Logical_Operator_out865_out1            : std_logic;
  SIGNAL Logical_Operator_out866_out1            : std_logic;
  SIGNAL Logical_Operator_out867_out1            : std_logic;
  SIGNAL Logical_Operator_out868_out1            : std_logic;
  SIGNAL Logical_Operator_out869_out1            : std_logic;
  SIGNAL Logical_Operator_out870_out1            : std_logic;
  SIGNAL Logical_Operator_out871_out1            : std_logic;
  SIGNAL Logical_Operator_out872_out1            : std_logic;
  SIGNAL Logical_Operator_out873_out1            : std_logic;
  SIGNAL Logical_Operator_out874_out1            : std_logic;
  SIGNAL Logical_Operator_out875_out1            : std_logic;
  SIGNAL Logical_Operator_out876_out1            : std_logic;
  SIGNAL Logical_Operator_out877_out1            : std_logic;
  SIGNAL Logical_Operator_out878_out1            : std_logic;
  SIGNAL Logical_Operator_out879_out1            : std_logic;
  SIGNAL Logical_Operator_out880_out1            : std_logic;
  SIGNAL Logical_Operator_out881_out1            : std_logic;
  SIGNAL Logical_Operator_out882_out1            : std_logic;
  SIGNAL Logical_Operator_out883_out1            : std_logic;
  SIGNAL Logical_Operator_out884_out1            : std_logic;
  SIGNAL Logical_Operator_out885_out1            : std_logic;
  SIGNAL Logical_Operator_out886_out1            : std_logic;
  SIGNAL Logical_Operator_out887_out1            : std_logic;
  SIGNAL Logical_Operator_out888_out1            : std_logic;
  SIGNAL Logical_Operator_out889_out1            : std_logic;
  SIGNAL Logical_Operator_out890_out1            : std_logic;
  SIGNAL Logical_Operator_out891_out1            : std_logic;
  SIGNAL Logical_Operator_out892_out1            : std_logic;
  SIGNAL Logical_Operator_out893_out1            : std_logic;
  SIGNAL Logical_Operator_out894_out1            : std_logic;
  SIGNAL Logical_Operator_out895_out1            : std_logic;
  SIGNAL Logical_Operator_out896_out1            : std_logic;
  SIGNAL Logical_Operator_out897_out1            : std_logic;
  SIGNAL Logical_Operator_out898_out1            : std_logic;
  SIGNAL Logical_Operator_out899_out1            : std_logic;
  SIGNAL Logical_Operator_out900_out1            : std_logic;
  SIGNAL Logical_Operator_out901_out1            : std_logic;
  SIGNAL Logical_Operator_out902_out1            : std_logic;
  SIGNAL Logical_Operator_out903_out1            : std_logic;
  SIGNAL Logical_Operator_out904_out1            : std_logic;
  SIGNAL Logical_Operator_out905_out1            : std_logic;
  SIGNAL Logical_Operator_out906_out1            : std_logic;
  SIGNAL Logical_Operator_out907_out1            : std_logic;
  SIGNAL Logical_Operator_out908_out1            : std_logic;
  SIGNAL Logical_Operator_out909_out1            : std_logic;
  SIGNAL Logical_Operator_out910_out1            : std_logic;
  SIGNAL Logical_Operator_out911_out1            : std_logic;
  SIGNAL Logical_Operator_out912_out1            : std_logic;
  SIGNAL Logical_Operator_out913_out1            : std_logic;
  SIGNAL Logical_Operator_out914_out1            : std_logic;
  SIGNAL Logical_Operator_out915_out1            : std_logic;
  SIGNAL Logical_Operator_out916_out1            : std_logic;
  SIGNAL Logical_Operator_out917_out1            : std_logic;
  SIGNAL Logical_Operator_out918_out1            : std_logic;
  SIGNAL Logical_Operator_out919_out1            : std_logic;
  SIGNAL Logical_Operator_out920_out1            : std_logic;
  SIGNAL Logical_Operator_out921_out1            : std_logic;
  SIGNAL Logical_Operator_out922_out1            : std_logic;
  SIGNAL Logical_Operator_out923_out1            : std_logic;
  SIGNAL Logical_Operator_out924_out1            : std_logic;
  SIGNAL Logical_Operator_out925_out1            : std_logic;
  SIGNAL Logical_Operator_out926_out1            : std_logic;
  SIGNAL Logical_Operator_out927_out1            : std_logic;
  SIGNAL Logical_Operator_out928_out1            : std_logic;
  SIGNAL Logical_Operator_out929_out1            : std_logic;
  SIGNAL Logical_Operator_out930_out1            : std_logic;
  SIGNAL Logical_Operator_out931_out1            : std_logic;
  SIGNAL Logical_Operator_out932_out1            : std_logic;
  SIGNAL Logical_Operator_out933_out1            : std_logic;
  SIGNAL Logical_Operator_out934_out1            : std_logic;
  SIGNAL Logical_Operator_out935_out1            : std_logic;
  SIGNAL Logical_Operator_out936_out1            : std_logic;
  SIGNAL Logical_Operator_out937_out1            : std_logic;
  SIGNAL Logical_Operator_out938_out1            : std_logic;
  SIGNAL Logical_Operator_out939_out1            : std_logic;
  SIGNAL Logical_Operator_out940_out1            : std_logic;
  SIGNAL Logical_Operator_out941_out1            : std_logic;
  SIGNAL Logical_Operator_out942_out1            : std_logic;
  SIGNAL Logical_Operator_out943_out1            : std_logic;
  SIGNAL Logical_Operator_out944_out1            : std_logic;
  SIGNAL Logical_Operator_out945_out1            : std_logic;
  SIGNAL Logical_Operator_out946_out1            : std_logic;
  SIGNAL Logical_Operator_out947_out1            : std_logic;
  SIGNAL Logical_Operator_out948_out1            : std_logic;
  SIGNAL Logical_Operator_out949_out1            : std_logic;
  SIGNAL Logical_Operator_out950_out1            : std_logic;
  SIGNAL Logical_Operator_out951_out1            : std_logic;
  SIGNAL Logical_Operator_out952_out1            : std_logic;
  SIGNAL Logical_Operator_out953_out1            : std_logic;
  SIGNAL Logical_Operator_out954_out1            : std_logic;
  SIGNAL Logical_Operator_out955_out1            : std_logic;
  SIGNAL Logical_Operator_out956_out1            : std_logic;
  SIGNAL Logical_Operator_out957_out1            : std_logic;
  SIGNAL Logical_Operator_out958_out1            : std_logic;
  SIGNAL Logical_Operator_out959_out1            : std_logic;
  SIGNAL Logical_Operator_out960_out1            : std_logic;
  SIGNAL Logical_Operator_out961_out1            : std_logic;
  SIGNAL Logical_Operator_out962_out1            : std_logic;
  SIGNAL Logical_Operator_out963_out1            : std_logic;
  SIGNAL Logical_Operator_out964_out1            : std_logic;
  SIGNAL Logical_Operator_out965_out1            : std_logic;
  SIGNAL Logical_Operator_out966_out1            : std_logic;
  SIGNAL Logical_Operator_out967_out1            : std_logic;
  SIGNAL Logical_Operator_out968_out1            : std_logic;
  SIGNAL Logical_Operator_out969_out1            : std_logic;
  SIGNAL Logical_Operator_out970_out1            : std_logic;
  SIGNAL Logical_Operator_out971_out1            : std_logic;
  SIGNAL Logical_Operator_out972_out1            : std_logic;
  SIGNAL Logical_Operator_out973_out1            : std_logic;
  SIGNAL Logical_Operator_out974_out1            : std_logic;
  SIGNAL Logical_Operator_out975_out1            : std_logic;
  SIGNAL Logical_Operator_out976_out1            : std_logic;
  SIGNAL Logical_Operator_out977_out1            : std_logic;
  SIGNAL Logical_Operator_out978_out1            : std_logic;
  SIGNAL Logical_Operator_out979_out1            : std_logic;
  SIGNAL Logical_Operator_out980_out1            : std_logic;
  SIGNAL Logical_Operator_out981_out1            : std_logic;
  SIGNAL Logical_Operator_out982_out1            : std_logic;
  SIGNAL Logical_Operator_out983_out1            : std_logic;
  SIGNAL Logical_Operator_out984_out1            : std_logic;
  SIGNAL Logical_Operator_out985_out1            : std_logic;
  SIGNAL Logical_Operator_out986_out1            : std_logic;
  SIGNAL Logical_Operator_out987_out1            : std_logic;
  SIGNAL Logical_Operator_out988_out1            : std_logic;
  SIGNAL Logical_Operator_out989_out1            : std_logic;
  SIGNAL Logical_Operator_out990_out1            : std_logic;
  SIGNAL Logical_Operator_out991_out1            : std_logic;
  SIGNAL Logical_Operator_out992_out1            : std_logic;
  SIGNAL Logical_Operator_out993_out1            : std_logic;
  SIGNAL Logical_Operator_out994_out1            : std_logic;
  SIGNAL Logical_Operator_out995_out1            : std_logic;
  SIGNAL Logical_Operator_out996_out1            : std_logic;
  SIGNAL Logical_Operator_out997_out1            : std_logic;
  SIGNAL Logical_Operator_out998_out1            : std_logic;
  SIGNAL Logical_Operator_out999_out1            : std_logic;
  SIGNAL Logical_Operator_out1000_out1            : std_logic;
  SIGNAL Logical_Operator_out1001_out1            : std_logic;
  SIGNAL Logical_Operator_out1002_out1            : std_logic;
  SIGNAL Logical_Operator_out1003_out1            : std_logic;
  SIGNAL Logical_Operator_out1004_out1            : std_logic;
  SIGNAL Logical_Operator_out1005_out1            : std_logic;
  SIGNAL Logical_Operator_out1006_out1            : std_logic;
  SIGNAL Logical_Operator_out1007_out1            : std_logic;
  SIGNAL Logical_Operator_out1008_out1            : std_logic;
  SIGNAL Logical_Operator_out1009_out1            : std_logic;
  SIGNAL Logical_Operator_out1010_out1            : std_logic;
  SIGNAL Logical_Operator_out1011_out1            : std_logic;
  SIGNAL Logical_Operator_out1012_out1            : std_logic;
  SIGNAL Logical_Operator_out1013_out1            : std_logic;
  SIGNAL Logical_Operator_out1014_out1            : std_logic;
  SIGNAL Logical_Operator_out1015_out1            : std_logic;
  SIGNAL Logical_Operator_out1016_out1            : std_logic;
  SIGNAL Logical_Operator_out1017_out1            : std_logic;
  SIGNAL Logical_Operator_out1018_out1            : std_logic;
  SIGNAL Logical_Operator_out1019_out1            : std_logic;
  SIGNAL Logical_Operator_out1020_out1            : std_logic;
  SIGNAL Logical_Operator_out1021_out1            : std_logic;
  SIGNAL Logical_Operator_out1022_out1            : std_logic;
  SIGNAL Logical_Operator_out1023_out1            : std_logic;
  SIGNAL Logical_Operator_out1024_out1            : std_logic;
  SIGNAL Logical_Operator_out1025_out1            : std_logic;
  SIGNAL Logical_Operator_out1026_out1            : std_logic;
  SIGNAL Logical_Operator_out1027_out1            : std_logic;
  SIGNAL Logical_Operator_out1028_out1            : std_logic;
  SIGNAL Logical_Operator_out1029_out1            : std_logic;
  SIGNAL Logical_Operator_out1030_out1            : std_logic;
  SIGNAL Logical_Operator_out1031_out1            : std_logic;
  SIGNAL Logical_Operator_out1032_out1            : std_logic;
  SIGNAL Logical_Operator_out1033_out1            : std_logic;
  SIGNAL Logical_Operator_out1034_out1            : std_logic;
  SIGNAL Logical_Operator_out1035_out1            : std_logic;
  SIGNAL Logical_Operator_out1036_out1            : std_logic;
  SIGNAL Logical_Operator_out1037_out1            : std_logic;
  SIGNAL Logical_Operator_out1038_out1            : std_logic;
  SIGNAL Logical_Operator_out1039_out1            : std_logic;
  SIGNAL Logical_Operator_out1040_out1            : std_logic;
  SIGNAL Logical_Operator_out1041_out1            : std_logic;
  SIGNAL Logical_Operator_out1042_out1            : std_logic;
  SIGNAL Logical_Operator_out1043_out1            : std_logic;
  SIGNAL Logical_Operator_out1044_out1            : std_logic;
  SIGNAL Logical_Operator_out1045_out1            : std_logic;
  SIGNAL Logical_Operator_out1046_out1            : std_logic;
  SIGNAL Logical_Operator_out1047_out1            : std_logic;
  SIGNAL Logical_Operator_out1048_out1            : std_logic;
  SIGNAL Logical_Operator_out1049_out1            : std_logic;
  SIGNAL Logical_Operator_out1050_out1            : std_logic;
  SIGNAL Logical_Operator_out1051_out1            : std_logic;
  SIGNAL Logical_Operator_out1052_out1            : std_logic;
  SIGNAL Logical_Operator_out1053_out1            : std_logic;
  SIGNAL Logical_Operator_out1054_out1            : std_logic;
  SIGNAL Logical_Operator_out1055_out1            : std_logic;
  SIGNAL Logical_Operator_out1056_out1            : std_logic;
  SIGNAL Logical_Operator_out1057_out1            : std_logic;
  SIGNAL Logical_Operator_out1058_out1            : std_logic;
  SIGNAL Logical_Operator_out1059_out1            : std_logic;
  SIGNAL Logical_Operator_out1060_out1            : std_logic;
  SIGNAL Logical_Operator_out1061_out1            : std_logic;
  SIGNAL Logical_Operator_out1062_out1            : std_logic;
  SIGNAL Logical_Operator_out1063_out1            : std_logic;
  SIGNAL Logical_Operator_out1064_out1            : std_logic;
  SIGNAL Logical_Operator_out1065_out1            : std_logic;
  SIGNAL Logical_Operator_out1066_out1            : std_logic;
  SIGNAL Logical_Operator_out1067_out1            : std_logic;
  SIGNAL Logical_Operator_out1068_out1            : std_logic;
  SIGNAL Logical_Operator_out1069_out1            : std_logic;
  SIGNAL Logical_Operator_out1070_out1            : std_logic;
  SIGNAL Logical_Operator_out1071_out1            : std_logic;
  SIGNAL Logical_Operator_out1072_out1            : std_logic;
  SIGNAL Logical_Operator_out1073_out1            : std_logic;
  SIGNAL Logical_Operator_out1074_out1            : std_logic;
  SIGNAL Logical_Operator_out1075_out1            : std_logic;
  SIGNAL Logical_Operator_out1076_out1            : std_logic;
  SIGNAL Logical_Operator_out1077_out1            : std_logic;
  SIGNAL Logical_Operator_out1078_out1            : std_logic;
  SIGNAL Logical_Operator_out1079_out1            : std_logic;
  SIGNAL Logical_Operator_out1080_out1            : std_logic;
  SIGNAL Logical_Operator_out1081_out1            : std_logic;
  SIGNAL Logical_Operator_out1082_out1            : std_logic;
  SIGNAL Logical_Operator_out1083_out1            : std_logic;
  SIGNAL Logical_Operator_out1084_out1            : std_logic;
  SIGNAL Logical_Operator_out1085_out1            : std_logic;
  SIGNAL Logical_Operator_out1086_out1            : std_logic;
  SIGNAL Logical_Operator_out1087_out1            : std_logic;
  SIGNAL Logical_Operator_out1088_out1            : std_logic;
  SIGNAL Logical_Operator_out1089_out1            : std_logic;
  SIGNAL Logical_Operator_out1090_out1            : std_logic;
  SIGNAL Logical_Operator_out1091_out1            : std_logic;
  SIGNAL Logical_Operator_out1092_out1            : std_logic;
  SIGNAL Logical_Operator_out1093_out1            : std_logic;
  SIGNAL Logical_Operator_out1094_out1            : std_logic;
  SIGNAL Logical_Operator_out1095_out1            : std_logic;
  SIGNAL Logical_Operator_out1096_out1            : std_logic;
  SIGNAL Logical_Operator_out1097_out1            : std_logic;
  SIGNAL Logical_Operator_out1098_out1            : std_logic;
  SIGNAL Logical_Operator_out1099_out1            : std_logic;
  SIGNAL Logical_Operator_out1100_out1            : std_logic;
  SIGNAL Logical_Operator_out1101_out1            : std_logic;
  SIGNAL Logical_Operator_out1102_out1            : std_logic;
  SIGNAL Logical_Operator_out1103_out1            : std_logic;
  SIGNAL Logical_Operator_out1104_out1            : std_logic;
  SIGNAL Logical_Operator_out1105_out1            : std_logic;
  SIGNAL Logical_Operator_out1106_out1            : std_logic;
  SIGNAL Logical_Operator_out1107_out1            : std_logic;
  SIGNAL Logical_Operator_out1108_out1            : std_logic;
  SIGNAL Logical_Operator_out1109_out1            : std_logic;
  SIGNAL Logical_Operator_out1110_out1            : std_logic;
  SIGNAL Logical_Operator_out1111_out1            : std_logic;
  SIGNAL Logical_Operator_out1112_out1            : std_logic;
  SIGNAL Logical_Operator_out1113_out1            : std_logic;
  SIGNAL Logical_Operator_out1114_out1            : std_logic;
  SIGNAL Logical_Operator_out1115_out1            : std_logic;
  SIGNAL Logical_Operator_out1116_out1            : std_logic;
  SIGNAL Logical_Operator_out1117_out1            : std_logic;
  SIGNAL Logical_Operator_out1118_out1            : std_logic;
  SIGNAL Logical_Operator_out1119_out1            : std_logic;
  SIGNAL Logical_Operator_out1120_out1            : std_logic;
  SIGNAL Logical_Operator_out1121_out1            : std_logic;
  SIGNAL Logical_Operator_out1122_out1            : std_logic;
  SIGNAL Logical_Operator_out1123_out1            : std_logic;
  SIGNAL Logical_Operator_out1124_out1            : std_logic;
  SIGNAL Logical_Operator_out1125_out1            : std_logic;
  SIGNAL Logical_Operator_out1126_out1            : std_logic;
  SIGNAL Logical_Operator_out1127_out1            : std_logic;
  SIGNAL Logical_Operator_out1128_out1            : std_logic;
  SIGNAL Logical_Operator_out1129_out1            : std_logic;
  SIGNAL Logical_Operator_out1130_out1            : std_logic;
  SIGNAL Logical_Operator_out1131_out1            : std_logic;
  SIGNAL Logical_Operator_out1132_out1            : std_logic;
  SIGNAL Logical_Operator_out1133_out1            : std_logic;
  SIGNAL Logical_Operator_out1134_out1            : std_logic;
  SIGNAL Logical_Operator_out1135_out1            : std_logic;
  SIGNAL Logical_Operator_out1136_out1            : std_logic;
  SIGNAL Logical_Operator_out1137_out1            : std_logic;
  SIGNAL Logical_Operator_out1138_out1            : std_logic;
  SIGNAL Logical_Operator_out1139_out1            : std_logic;
  SIGNAL Logical_Operator_out1140_out1            : std_logic;
  SIGNAL Logical_Operator_out1141_out1            : std_logic;
  SIGNAL Logical_Operator_out1142_out1            : std_logic;
  SIGNAL Logical_Operator_out1143_out1            : std_logic;
  SIGNAL Logical_Operator_out1144_out1            : std_logic;
  SIGNAL Logical_Operator_out1145_out1            : std_logic;
  SIGNAL Logical_Operator_out1146_out1            : std_logic;
  SIGNAL Logical_Operator_out1147_out1            : std_logic;
  SIGNAL Logical_Operator_out1148_out1            : std_logic;
  SIGNAL Logical_Operator_out1149_out1            : std_logic;
  SIGNAL Logical_Operator_out1150_out1            : std_logic;
  SIGNAL Logical_Operator_out1151_out1            : std_logic;
  SIGNAL Logical_Operator_out1152_out1            : std_logic;
  SIGNAL Logical_Operator_out1153_out1            : std_logic;
  SIGNAL Logical_Operator_out1154_out1            : std_logic;
  SIGNAL Logical_Operator_out1155_out1            : std_logic;
  SIGNAL Logical_Operator_out1156_out1            : std_logic;
  SIGNAL Logical_Operator_out1157_out1            : std_logic;
  SIGNAL Logical_Operator_out1158_out1            : std_logic;
  SIGNAL Logical_Operator_out1159_out1            : std_logic;
  SIGNAL Logical_Operator_out1160_out1            : std_logic;
  SIGNAL Logical_Operator_out1161_out1            : std_logic;
  SIGNAL Logical_Operator_out1162_out1            : std_logic;
  SIGNAL Logical_Operator_out1163_out1            : std_logic;
  SIGNAL Logical_Operator_out1164_out1            : std_logic;
  SIGNAL Logical_Operator_out1165_out1            : std_logic;
  SIGNAL Logical_Operator_out1166_out1            : std_logic;
  SIGNAL Logical_Operator_out1167_out1            : std_logic;
  SIGNAL Logical_Operator_out1168_out1            : std_logic;
  SIGNAL Logical_Operator_out1169_out1            : std_logic;
  SIGNAL Logical_Operator_out1170_out1            : std_logic;
  SIGNAL Logical_Operator_out1171_out1            : std_logic;
  SIGNAL Logical_Operator_out1172_out1            : std_logic;
  SIGNAL Logical_Operator_out1173_out1            : std_logic;
  SIGNAL Logical_Operator_out1174_out1            : std_logic;
  SIGNAL Logical_Operator_out1175_out1            : std_logic;
  SIGNAL Logical_Operator_out1176_out1            : std_logic;
  SIGNAL Logical_Operator_out1177_out1            : std_logic;
  SIGNAL Logical_Operator_out1178_out1            : std_logic;
  SIGNAL Logical_Operator_out1179_out1            : std_logic;
  SIGNAL Logical_Operator_out1180_out1            : std_logic;
  SIGNAL Logical_Operator_out1181_out1            : std_logic;
  SIGNAL Logical_Operator_out1182_out1            : std_logic;
  SIGNAL Logical_Operator_out1183_out1            : std_logic;
  SIGNAL Logical_Operator_out1184_out1            : std_logic;
  SIGNAL Logical_Operator_out1185_out1            : std_logic;
  SIGNAL Logical_Operator_out1186_out1            : std_logic;
  SIGNAL Logical_Operator_out1187_out1            : std_logic;
  SIGNAL Logical_Operator_out1188_out1            : std_logic;
  SIGNAL Logical_Operator_out1189_out1            : std_logic;
  SIGNAL Logical_Operator_out1190_out1            : std_logic;
  SIGNAL Logical_Operator_out1191_out1            : std_logic;
  SIGNAL Logical_Operator_out1192_out1            : std_logic;
  SIGNAL Logical_Operator_out1193_out1            : std_logic;
  SIGNAL Logical_Operator_out1194_out1            : std_logic;
  SIGNAL Logical_Operator_out1195_out1            : std_logic;
  SIGNAL Logical_Operator_out1196_out1            : std_logic;
  SIGNAL Logical_Operator_out1197_out1            : std_logic;
  SIGNAL Logical_Operator_out1198_out1            : std_logic;
  SIGNAL Logical_Operator_out1199_out1            : std_logic;
  SIGNAL Logical_Operator_out1200_out1            : std_logic;
  SIGNAL Logical_Operator_out1201_out1            : std_logic;
  SIGNAL Logical_Operator_out1202_out1            : std_logic;
  SIGNAL Logical_Operator_out1203_out1            : std_logic;
  SIGNAL Logical_Operator_out1204_out1            : std_logic;
  SIGNAL Logical_Operator_out1205_out1            : std_logic;
  SIGNAL Logical_Operator_out1206_out1            : std_logic;
  SIGNAL Logical_Operator_out1207_out1            : std_logic;
  SIGNAL Logical_Operator_out1208_out1            : std_logic;
  SIGNAL Logical_Operator_out1209_out1            : std_logic;
  SIGNAL Logical_Operator_out1210_out1            : std_logic;
  SIGNAL Logical_Operator_out1211_out1            : std_logic;
  SIGNAL Logical_Operator_out1212_out1            : std_logic;
  SIGNAL Logical_Operator_out1213_out1            : std_logic;
  SIGNAL Logical_Operator_out1214_out1            : std_logic;
  SIGNAL Logical_Operator_out1215_out1            : std_logic;
  SIGNAL Logical_Operator_out1216_out1            : std_logic;
  SIGNAL Logical_Operator_out1217_out1            : std_logic;
  SIGNAL Logical_Operator_out1218_out1            : std_logic;
  SIGNAL Logical_Operator_out1219_out1            : std_logic;
  SIGNAL Logical_Operator_out1220_out1            : std_logic;
  SIGNAL Logical_Operator_out1221_out1            : std_logic;
  SIGNAL Logical_Operator_out1222_out1            : std_logic;
  SIGNAL Logical_Operator_out1223_out1            : std_logic;
  SIGNAL Logical_Operator_out1224_out1            : std_logic;
  SIGNAL Logical_Operator_out1225_out1            : std_logic;
  SIGNAL Logical_Operator_out1226_out1            : std_logic;
  SIGNAL Logical_Operator_out1227_out1            : std_logic;
  SIGNAL Logical_Operator_out1228_out1            : std_logic;
  SIGNAL Logical_Operator_out1229_out1            : std_logic;
  SIGNAL Logical_Operator_out1230_out1            : std_logic;
  SIGNAL Logical_Operator_out1231_out1            : std_logic;
  SIGNAL Logical_Operator_out1232_out1            : std_logic;
  SIGNAL Logical_Operator_out1233_out1            : std_logic;
  SIGNAL Logical_Operator_out1234_out1            : std_logic;
  SIGNAL Logical_Operator_out1235_out1            : std_logic;
  SIGNAL Logical_Operator_out1236_out1            : std_logic;
  SIGNAL Logical_Operator_out1237_out1            : std_logic;
  SIGNAL Logical_Operator_out1238_out1            : std_logic;
  SIGNAL Logical_Operator_out1239_out1            : std_logic;
  SIGNAL Logical_Operator_out1240_out1            : std_logic;
  SIGNAL Logical_Operator_out1241_out1            : std_logic;
  SIGNAL Logical_Operator_out1242_out1            : std_logic;
  SIGNAL Logical_Operator_out1243_out1            : std_logic;
  SIGNAL Logical_Operator_out1244_out1            : std_logic;
  SIGNAL Logical_Operator_out1245_out1            : std_logic;
  SIGNAL Logical_Operator_out1246_out1            : std_logic;
  SIGNAL Logical_Operator_out1247_out1            : std_logic;
  SIGNAL Logical_Operator_out1248_out1            : std_logic;
  SIGNAL Logical_Operator_out1249_out1            : std_logic;
  SIGNAL Logical_Operator_out1250_out1            : std_logic;
  SIGNAL Logical_Operator_out1251_out1            : std_logic;
  SIGNAL Logical_Operator_out1252_out1            : std_logic;
  SIGNAL Logical_Operator_out1253_out1            : std_logic;
  SIGNAL Logical_Operator_out1254_out1            : std_logic;
  SIGNAL Logical_Operator_out1255_out1            : std_logic;
  SIGNAL Logical_Operator_out1256_out1            : std_logic;
  SIGNAL Logical_Operator_out1257_out1            : std_logic;
  SIGNAL Logical_Operator_out1258_out1            : std_logic;
  SIGNAL Logical_Operator_out1259_out1            : std_logic;
  SIGNAL Logical_Operator_out1260_out1            : std_logic;
  SIGNAL Logical_Operator_out1261_out1            : std_logic;
  SIGNAL Logical_Operator_out1262_out1            : std_logic;
  SIGNAL Logical_Operator_out1263_out1            : std_logic;
  SIGNAL Logical_Operator_out1264_out1            : std_logic;
  SIGNAL Logical_Operator_out1265_out1            : std_logic;
  SIGNAL Logical_Operator_out1266_out1            : std_logic;
  SIGNAL Logical_Operator_out1267_out1            : std_logic;
  SIGNAL Logical_Operator_out1268_out1            : std_logic;
  SIGNAL Logical_Operator_out1269_out1            : std_logic;
  SIGNAL Logical_Operator_out1270_out1            : std_logic;
  SIGNAL Logical_Operator_out1271_out1            : std_logic;
  SIGNAL Logical_Operator_out1272_out1            : std_logic;
  SIGNAL Logical_Operator_out1273_out1            : std_logic;
  SIGNAL Logical_Operator_out1274_out1            : std_logic;
  SIGNAL Logical_Operator_out1275_out1            : std_logic;
  SIGNAL Logical_Operator_out1276_out1            : std_logic;
  SIGNAL Logical_Operator_out1277_out1            : std_logic;
  SIGNAL Logical_Operator_out1278_out1            : std_logic;
  SIGNAL Logical_Operator_out1279_out1            : std_logic;
  SIGNAL Logical_Operator_out1280_out1            : std_logic;
  SIGNAL Logical_Operator_out1281_out1            : std_logic;
  SIGNAL Logical_Operator_out1282_out1            : std_logic;
  SIGNAL Logical_Operator_out1283_out1            : std_logic;
  SIGNAL Logical_Operator_out1284_out1            : std_logic;
  SIGNAL Logical_Operator_out1285_out1            : std_logic;
  SIGNAL Logical_Operator_out1286_out1            : std_logic;
  SIGNAL Logical_Operator_out1287_out1            : std_logic;
  SIGNAL Logical_Operator_out1288_out1            : std_logic;
  SIGNAL Logical_Operator_out1289_out1            : std_logic;
  SIGNAL Logical_Operator_out1290_out1            : std_logic;
  SIGNAL Logical_Operator_out1291_out1            : std_logic;
  SIGNAL Logical_Operator_out1292_out1            : std_logic;
  SIGNAL Logical_Operator_out1293_out1            : std_logic;
  SIGNAL Logical_Operator_out1294_out1            : std_logic;
  SIGNAL Logical_Operator_out1295_out1            : std_logic;
  SIGNAL Logical_Operator_out1296_out1            : std_logic;
  SIGNAL Logical_Operator_out1297_out1            : std_logic;
  SIGNAL Logical_Operator_out1298_out1            : std_logic;
  SIGNAL Logical_Operator_out1299_out1            : std_logic;
  SIGNAL Logical_Operator_out1300_out1            : std_logic;
  SIGNAL Logical_Operator_out1301_out1            : std_logic;
  SIGNAL Logical_Operator_out1302_out1            : std_logic;
  SIGNAL Logical_Operator_out1303_out1            : std_logic;
  SIGNAL Logical_Operator_out1304_out1            : std_logic;
  SIGNAL Logical_Operator_out1305_out1            : std_logic;
  SIGNAL Logical_Operator_out1306_out1            : std_logic;
  SIGNAL Logical_Operator_out1307_out1            : std_logic;
  SIGNAL Logical_Operator_out1308_out1            : std_logic;
  SIGNAL Logical_Operator_out1309_out1            : std_logic;
  SIGNAL Logical_Operator_out1310_out1            : std_logic;
  SIGNAL Logical_Operator_out1311_out1            : std_logic;
  SIGNAL Logical_Operator_out1312_out1            : std_logic;
  SIGNAL Logical_Operator_out1313_out1            : std_logic;
  SIGNAL Logical_Operator_out1314_out1            : std_logic;
  SIGNAL Logical_Operator_out1315_out1            : std_logic;
  SIGNAL Logical_Operator_out1316_out1            : std_logic;
  SIGNAL Logical_Operator_out1317_out1            : std_logic;
  SIGNAL Logical_Operator_out1318_out1            : std_logic;
  SIGNAL Logical_Operator_out1319_out1            : std_logic;
  SIGNAL Logical_Operator_out1320_out1            : std_logic;
  SIGNAL Logical_Operator_out1321_out1            : std_logic;
  SIGNAL Logical_Operator_out1322_out1            : std_logic;
  SIGNAL Logical_Operator_out1323_out1            : std_logic;
  SIGNAL Logical_Operator_out1324_out1            : std_logic;
  SIGNAL Logical_Operator_out1325_out1            : std_logic;
  SIGNAL Logical_Operator_out1326_out1            : std_logic;
  SIGNAL Logical_Operator_out1327_out1            : std_logic;
  SIGNAL Logical_Operator_out1328_out1            : std_logic;
  SIGNAL Logical_Operator_out1329_out1            : std_logic;
  SIGNAL Logical_Operator_out1330_out1            : std_logic;
  SIGNAL Logical_Operator_out1331_out1            : std_logic;
  SIGNAL Logical_Operator_out1332_out1            : std_logic;
  SIGNAL Logical_Operator_out1333_out1            : std_logic;
  SIGNAL Logical_Operator_out1334_out1            : std_logic;
  SIGNAL Logical_Operator_out1335_out1            : std_logic;
  SIGNAL Logical_Operator_out1336_out1            : std_logic;
  SIGNAL Logical_Operator_out1337_out1            : std_logic;
  SIGNAL Logical_Operator_out1338_out1            : std_logic;
  SIGNAL Logical_Operator_out1339_out1            : std_logic;
  SIGNAL Logical_Operator_out1340_out1            : std_logic;
  SIGNAL Logical_Operator_out1341_out1            : std_logic;
  SIGNAL Logical_Operator_out1342_out1            : std_logic;
  SIGNAL Logical_Operator_out1343_out1            : std_logic;
  SIGNAL Logical_Operator_out1344_out1            : std_logic;
  SIGNAL Logical_Operator_out1345_out1            : std_logic;
  SIGNAL Logical_Operator_out1346_out1            : std_logic;
  SIGNAL Logical_Operator_out1347_out1            : std_logic;
  SIGNAL Logical_Operator_out1348_out1            : std_logic;
  SIGNAL Logical_Operator_out1349_out1            : std_logic;
  SIGNAL Logical_Operator_out1350_out1            : std_logic;
  SIGNAL Logical_Operator_out1351_out1            : std_logic;
  SIGNAL Logical_Operator_out1352_out1            : std_logic;
  SIGNAL Logical_Operator_out1353_out1            : std_logic;
  SIGNAL Logical_Operator_out1354_out1            : std_logic;
  SIGNAL Logical_Operator_out1355_out1            : std_logic;
  SIGNAL Logical_Operator_out1356_out1            : std_logic;
  SIGNAL Logical_Operator_out1357_out1            : std_logic;
  SIGNAL Logical_Operator_out1358_out1            : std_logic;
  SIGNAL Logical_Operator_out1359_out1            : std_logic;
  SIGNAL Logical_Operator_out1360_out1            : std_logic;
  SIGNAL Logical_Operator_out1361_out1            : std_logic;
  SIGNAL Logical_Operator_out1362_out1            : std_logic;
  SIGNAL Logical_Operator_out1363_out1            : std_logic;
  SIGNAL Logical_Operator_out1364_out1            : std_logic;
  SIGNAL Logical_Operator_out1365_out1            : std_logic;
  SIGNAL Logical_Operator_out1366_out1            : std_logic;
  SIGNAL Logical_Operator_out1367_out1            : std_logic;
  SIGNAL Logical_Operator_out1368_out1            : std_logic;
  SIGNAL Logical_Operator_out1369_out1            : std_logic;
  SIGNAL Logical_Operator_out1370_out1            : std_logic;
  SIGNAL Logical_Operator_out1371_out1            : std_logic;
  SIGNAL Logical_Operator_out1372_out1            : std_logic;
  SIGNAL Logical_Operator_out1373_out1            : std_logic;
  SIGNAL Logical_Operator_out1374_out1            : std_logic;
  SIGNAL Logical_Operator_out1375_out1            : std_logic;
  SIGNAL Logical_Operator_out1376_out1            : std_logic;
  SIGNAL Logical_Operator_out1377_out1            : std_logic;
  SIGNAL Logical_Operator_out1378_out1            : std_logic;
  SIGNAL Logical_Operator_out1379_out1            : std_logic;
  SIGNAL Logical_Operator_out1380_out1            : std_logic;
  SIGNAL Logical_Operator_out1381_out1            : std_logic;
  SIGNAL Logical_Operator_out1382_out1            : std_logic;
  SIGNAL Logical_Operator_out1383_out1            : std_logic;
  SIGNAL Logical_Operator_out1384_out1            : std_logic;
  SIGNAL Logical_Operator_out1385_out1            : std_logic;
  SIGNAL Logical_Operator_out1386_out1            : std_logic;
  SIGNAL Logical_Operator_out1387_out1            : std_logic;
  SIGNAL Logical_Operator_out1388_out1            : std_logic;
  SIGNAL Logical_Operator_out1389_out1            : std_logic;
  SIGNAL Logical_Operator_out1390_out1            : std_logic;
  SIGNAL Logical_Operator_out1391_out1            : std_logic;
  SIGNAL Logical_Operator_out1392_out1            : std_logic;
  SIGNAL Logical_Operator_out1393_out1            : std_logic;
  SIGNAL Logical_Operator_out1394_out1            : std_logic;
  SIGNAL Logical_Operator_out1395_out1            : std_logic;
  SIGNAL Logical_Operator_out1396_out1            : std_logic;
  SIGNAL Logical_Operator_out1397_out1            : std_logic;
  SIGNAL Logical_Operator_out1398_out1            : std_logic;
  SIGNAL Logical_Operator_out1399_out1            : std_logic;
  SIGNAL Logical_Operator_out1400_out1            : std_logic;
  SIGNAL Logical_Operator_out1401_out1            : std_logic;
  SIGNAL Logical_Operator_out1402_out1            : std_logic;
  SIGNAL Logical_Operator_out1403_out1            : std_logic;
  SIGNAL Logical_Operator_out1404_out1            : std_logic;
  SIGNAL Logical_Operator_out1405_out1            : std_logic;
  SIGNAL Logical_Operator_out1406_out1            : std_logic;
  SIGNAL Logical_Operator_out1407_out1            : std_logic;
  SIGNAL Logical_Operator_out1408_out1            : std_logic;
  SIGNAL Logical_Operator_out1409_out1            : std_logic;
  SIGNAL Logical_Operator_out1410_out1            : std_logic;
  SIGNAL Logical_Operator_out1411_out1            : std_logic;
  SIGNAL Logical_Operator_out1412_out1            : std_logic;
  SIGNAL Logical_Operator_out1413_out1            : std_logic;
  SIGNAL Logical_Operator_out1414_out1            : std_logic;
  SIGNAL Logical_Operator_out1415_out1            : std_logic;
  SIGNAL Logical_Operator_out1416_out1            : std_logic;
  SIGNAL Logical_Operator_out1417_out1            : std_logic;
  SIGNAL Logical_Operator_out1418_out1            : std_logic;
  SIGNAL Logical_Operator_out1419_out1            : std_logic;
  SIGNAL Logical_Operator_out1420_out1            : std_logic;
  SIGNAL Logical_Operator_out1421_out1            : std_logic;
  SIGNAL Logical_Operator_out1422_out1            : std_logic;
  SIGNAL Logical_Operator_out1423_out1            : std_logic;
  SIGNAL Logical_Operator_out1424_out1            : std_logic;
  SIGNAL Logical_Operator_out1425_out1            : std_logic;
  SIGNAL Logical_Operator_out1426_out1            : std_logic;
  SIGNAL Logical_Operator_out1427_out1            : std_logic;
  SIGNAL Logical_Operator_out1428_out1            : std_logic;
  SIGNAL Logical_Operator_out1429_out1            : std_logic;
  SIGNAL Logical_Operator_out1430_out1            : std_logic;
  SIGNAL Logical_Operator_out1431_out1            : std_logic;
  SIGNAL Logical_Operator_out1432_out1            : std_logic;
  SIGNAL Logical_Operator_out1433_out1            : std_logic;
  SIGNAL Logical_Operator_out1434_out1            : std_logic;
  SIGNAL Logical_Operator_out1435_out1            : std_logic;
  SIGNAL Logical_Operator_out1436_out1            : std_logic;
  SIGNAL Logical_Operator_out1437_out1            : std_logic;
  SIGNAL Logical_Operator_out1438_out1            : std_logic;
  SIGNAL Logical_Operator_out1439_out1            : std_logic;
  SIGNAL Logical_Operator_out1440_out1            : std_logic;
  SIGNAL Logical_Operator_out1441_out1            : std_logic;
  SIGNAL Logical_Operator_out1442_out1            : std_logic;
  SIGNAL Logical_Operator_out1443_out1            : std_logic;
  SIGNAL Logical_Operator_out1444_out1            : std_logic;
  SIGNAL Logical_Operator_out1445_out1            : std_logic;
  SIGNAL Logical_Operator_out1446_out1            : std_logic;
  SIGNAL Logical_Operator_out1447_out1            : std_logic;
  SIGNAL Logical_Operator_out1448_out1            : std_logic;
  SIGNAL Logical_Operator_out1449_out1            : std_logic;
  SIGNAL Logical_Operator_out1450_out1            : std_logic;
  SIGNAL Logical_Operator_out1451_out1            : std_logic;
  SIGNAL Logical_Operator_out1452_out1            : std_logic;
  SIGNAL Logical_Operator_out1453_out1            : std_logic;
  SIGNAL Logical_Operator_out1454_out1            : std_logic;
  SIGNAL Logical_Operator_out1455_out1            : std_logic;
  SIGNAL Logical_Operator_out1456_out1            : std_logic;
  SIGNAL Logical_Operator_out1457_out1            : std_logic;
  SIGNAL Logical_Operator_out1458_out1            : std_logic;
  SIGNAL Logical_Operator_out1459_out1            : std_logic;
  SIGNAL Logical_Operator_out1460_out1            : std_logic;
  SIGNAL Logical_Operator_out1461_out1            : std_logic;
  SIGNAL Logical_Operator_out1462_out1            : std_logic;
  SIGNAL Logical_Operator_out1463_out1            : std_logic;
  SIGNAL Logical_Operator_out1464_out1            : std_logic;
  SIGNAL Logical_Operator_out1465_out1            : std_logic;
  SIGNAL Logical_Operator_out1466_out1            : std_logic;
  SIGNAL Logical_Operator_out1467_out1            : std_logic;
  SIGNAL Logical_Operator_out1468_out1            : std_logic;
  SIGNAL Logical_Operator_out1469_out1            : std_logic;
  SIGNAL Logical_Operator_out1470_out1            : std_logic;
  SIGNAL Logical_Operator_out1471_out1            : std_logic;
  SIGNAL Logical_Operator_out1472_out1            : std_logic;
  SIGNAL Logical_Operator_out1473_out1            : std_logic;
  SIGNAL Logical_Operator_out1474_out1            : std_logic;
  SIGNAL Logical_Operator_out1475_out1            : std_logic;
  SIGNAL Logical_Operator_out1476_out1            : std_logic;
  SIGNAL Logical_Operator_out1477_out1            : std_logic;
  SIGNAL Logical_Operator_out1478_out1            : std_logic;
  SIGNAL Logical_Operator_out1479_out1            : std_logic;
  SIGNAL Logical_Operator_out1480_out1            : std_logic;
  SIGNAL Logical_Operator_out1481_out1            : std_logic;
  SIGNAL Logical_Operator_out1482_out1            : std_logic;
  SIGNAL Logical_Operator_out1483_out1            : std_logic;
  SIGNAL Logical_Operator_out1484_out1            : std_logic;
  SIGNAL Logical_Operator_out1485_out1            : std_logic;
  SIGNAL Logical_Operator_out1486_out1            : std_logic;
  SIGNAL Logical_Operator_out1487_out1            : std_logic;
  SIGNAL Logical_Operator_out1488_out1            : std_logic;
  SIGNAL Logical_Operator_out1489_out1            : std_logic;
  SIGNAL Logical_Operator_out1490_out1            : std_logic;
  SIGNAL Logical_Operator_out1491_out1            : std_logic;
  SIGNAL Logical_Operator_out1492_out1            : std_logic;
  SIGNAL Logical_Operator_out1493_out1            : std_logic;
  SIGNAL Logical_Operator_out1494_out1            : std_logic;
  SIGNAL Logical_Operator_out1495_out1            : std_logic;
  SIGNAL Logical_Operator_out1496_out1            : std_logic;
  SIGNAL Logical_Operator_out1497_out1            : std_logic;
  SIGNAL Logical_Operator_out1498_out1            : std_logic;
  SIGNAL Logical_Operator_out1499_out1            : std_logic;
  SIGNAL Logical_Operator_out1500_out1            : std_logic;
  SIGNAL Logical_Operator_out1501_out1            : std_logic;
  SIGNAL Logical_Operator_out1502_out1            : std_logic;
  SIGNAL Logical_Operator_out1503_out1            : std_logic;
  SIGNAL Logical_Operator_out1504_out1            : std_logic;
  SIGNAL Logical_Operator_out1505_out1            : std_logic;
  SIGNAL Logical_Operator_out1506_out1            : std_logic;
  SIGNAL Logical_Operator_out1507_out1            : std_logic;
  SIGNAL Logical_Operator_out1508_out1            : std_logic;
  SIGNAL Logical_Operator_out1509_out1            : std_logic;
  SIGNAL Logical_Operator_out1510_out1            : std_logic;
  SIGNAL Logical_Operator_out1511_out1            : std_logic;
  SIGNAL Logical_Operator_out1512_out1            : std_logic;
  SIGNAL Logical_Operator_out1513_out1            : std_logic;
  SIGNAL Logical_Operator_out1514_out1            : std_logic;
  SIGNAL Logical_Operator_out1515_out1            : std_logic;
  SIGNAL Logical_Operator_out1516_out1            : std_logic;
  SIGNAL Logical_Operator_out1517_out1            : std_logic;
  SIGNAL Logical_Operator_out1518_out1            : std_logic;
  SIGNAL Logical_Operator_out1519_out1            : std_logic;
  SIGNAL Logical_Operator_out1520_out1            : std_logic;
  SIGNAL Logical_Operator_out1521_out1            : std_logic;
  SIGNAL Logical_Operator_out1522_out1            : std_logic;
  SIGNAL Logical_Operator_out1523_out1            : std_logic;
  SIGNAL Logical_Operator_out1524_out1            : std_logic;
  SIGNAL Logical_Operator_out1525_out1            : std_logic;
  SIGNAL Logical_Operator_out1526_out1            : std_logic;
  SIGNAL Logical_Operator_out1527_out1            : std_logic;
  SIGNAL Logical_Operator_out1528_out1            : std_logic;
  SIGNAL Logical_Operator_out1529_out1            : std_logic;
  SIGNAL Logical_Operator_out1530_out1            : std_logic;
  SIGNAL Logical_Operator_out1531_out1            : std_logic;
  SIGNAL Logical_Operator_out1532_out1            : std_logic;
  SIGNAL Logical_Operator_out1533_out1            : std_logic;
  SIGNAL Logical_Operator_out1534_out1            : std_logic;
  SIGNAL Logical_Operator_out1535_out1            : std_logic;
  SIGNAL Logical_Operator_out1536_out1            : std_logic;
  SIGNAL Logical_Operator_out1537_out1            : std_logic;
  SIGNAL Logical_Operator_out1538_out1            : std_logic;
  SIGNAL Logical_Operator_out1539_out1            : std_logic;
  SIGNAL Logical_Operator_out1540_out1            : std_logic;
  SIGNAL Logical_Operator_out1541_out1            : std_logic;
  SIGNAL Logical_Operator_out1542_out1            : std_logic;
  SIGNAL Logical_Operator_out1543_out1            : std_logic;
  SIGNAL Logical_Operator_out1544_out1            : std_logic;
  SIGNAL Logical_Operator_out1545_out1            : std_logic;
  SIGNAL Logical_Operator_out1546_out1            : std_logic;
  SIGNAL Logical_Operator_out1547_out1            : std_logic;
  SIGNAL Logical_Operator_out1548_out1            : std_logic;
  SIGNAL Logical_Operator_out1549_out1            : std_logic;
  SIGNAL Logical_Operator_out1550_out1            : std_logic;
  SIGNAL Logical_Operator_out1551_out1            : std_logic;
  SIGNAL Logical_Operator_out1552_out1            : std_logic;
  SIGNAL Logical_Operator_out1553_out1            : std_logic;
  SIGNAL Logical_Operator_out1554_out1            : std_logic;
  SIGNAL Logical_Operator_out1555_out1            : std_logic;
  SIGNAL Logical_Operator_out1556_out1            : std_logic;
  SIGNAL Logical_Operator_out1557_out1            : std_logic;
  SIGNAL Logical_Operator_out1558_out1            : std_logic;
  SIGNAL Logical_Operator_out1559_out1            : std_logic;
  SIGNAL Logical_Operator_out1560_out1            : std_logic;
  SIGNAL Logical_Operator_out1561_out1            : std_logic;
  SIGNAL Logical_Operator_out1562_out1            : std_logic;
  SIGNAL Logical_Operator_out1563_out1            : std_logic;
  SIGNAL Logical_Operator_out1564_out1            : std_logic;
  SIGNAL Logical_Operator_out1565_out1            : std_logic;
  SIGNAL Logical_Operator_out1566_out1            : std_logic;
  SIGNAL Logical_Operator_out1567_out1            : std_logic;
  SIGNAL Logical_Operator_out1568_out1            : std_logic;
  SIGNAL Logical_Operator_out1569_out1            : std_logic;
  SIGNAL Logical_Operator_out1570_out1            : std_logic;
  SIGNAL Logical_Operator_out1571_out1            : std_logic;
  SIGNAL Logical_Operator_out1572_out1            : std_logic;
  SIGNAL Logical_Operator_out1573_out1            : std_logic;
  SIGNAL Logical_Operator_out1574_out1            : std_logic;
  SIGNAL Logical_Operator_out1575_out1            : std_logic;
  SIGNAL Logical_Operator_out1576_out1            : std_logic;
  SIGNAL Logical_Operator_out1577_out1            : std_logic;
  SIGNAL Logical_Operator_out1578_out1            : std_logic;
  SIGNAL Logical_Operator_out1579_out1            : std_logic;
  SIGNAL Logical_Operator_out1580_out1            : std_logic;
  SIGNAL Logical_Operator_out1581_out1            : std_logic;
  SIGNAL Logical_Operator_out1582_out1            : std_logic;
  SIGNAL Logical_Operator_out1583_out1            : std_logic;
  SIGNAL Logical_Operator_out1584_out1            : std_logic;
  SIGNAL Logical_Operator_out1585_out1            : std_logic;
  SIGNAL Logical_Operator_out1586_out1            : std_logic;
  SIGNAL Logical_Operator_out1587_out1            : std_logic;
  SIGNAL Logical_Operator_out1588_out1            : std_logic;
  SIGNAL Logical_Operator_out1589_out1            : std_logic;
  SIGNAL Logical_Operator_out1590_out1            : std_logic;
  SIGNAL Logical_Operator_out1591_out1            : std_logic;
  SIGNAL Logical_Operator_out1592_out1            : std_logic;
  SIGNAL Logical_Operator_out1593_out1            : std_logic;
  SIGNAL Logical_Operator_out1594_out1            : std_logic;
  SIGNAL Logical_Operator_out1595_out1            : std_logic;
  SIGNAL Logical_Operator_out1596_out1            : std_logic;
  SIGNAL Logical_Operator_out1597_out1            : std_logic;
  SIGNAL Logical_Operator_out1598_out1            : std_logic;
  SIGNAL Logical_Operator_out1599_out1            : std_logic;
  SIGNAL Logical_Operator_out1600_out1            : std_logic;
  SIGNAL Logical_Operator_out1601_out1            : std_logic;
  SIGNAL Logical_Operator_out1602_out1            : std_logic;
  SIGNAL Logical_Operator_out1603_out1            : std_logic;
  SIGNAL Logical_Operator_out1604_out1            : std_logic;
  SIGNAL Logical_Operator_out1605_out1            : std_logic;
  SIGNAL Logical_Operator_out1606_out1            : std_logic;
  SIGNAL Logical_Operator_out1607_out1            : std_logic;
  SIGNAL Logical_Operator_out1608_out1            : std_logic;
  SIGNAL Logical_Operator_out1609_out1            : std_logic;
  SIGNAL Logical_Operator_out1610_out1            : std_logic;
  SIGNAL Logical_Operator_out1611_out1            : std_logic;
  SIGNAL Logical_Operator_out1612_out1            : std_logic;
  SIGNAL Logical_Operator_out1613_out1            : std_logic;
  SIGNAL Logical_Operator_out1614_out1            : std_logic;
  SIGNAL Logical_Operator_out1615_out1            : std_logic;
  SIGNAL Logical_Operator_out1616_out1            : std_logic;
  SIGNAL Logical_Operator_out1617_out1            : std_logic;
  SIGNAL Logical_Operator_out1618_out1            : std_logic;
  SIGNAL Logical_Operator_out1619_out1            : std_logic;
  SIGNAL Logical_Operator_out1620_out1            : std_logic;
  SIGNAL Logical_Operator_out1621_out1            : std_logic;
  SIGNAL Logical_Operator_out1622_out1            : std_logic;
  SIGNAL Logical_Operator_out1623_out1            : std_logic;
  SIGNAL Logical_Operator_out1624_out1            : std_logic;
  SIGNAL Logical_Operator_out1625_out1            : std_logic;
  SIGNAL Logical_Operator_out1626_out1            : std_logic;
  SIGNAL Logical_Operator_out1627_out1            : std_logic;
  SIGNAL Logical_Operator_out1628_out1            : std_logic;
  SIGNAL Logical_Operator_out1629_out1            : std_logic;
  SIGNAL Logical_Operator_out1630_out1            : std_logic;
  SIGNAL Logical_Operator_out1631_out1            : std_logic;
  SIGNAL Logical_Operator_out1632_out1            : std_logic;
  SIGNAL Logical_Operator_out1633_out1            : std_logic;
  SIGNAL Logical_Operator_out1634_out1            : std_logic;
  SIGNAL Logical_Operator_out1635_out1            : std_logic;
  SIGNAL Logical_Operator_out1636_out1            : std_logic;
  SIGNAL Logical_Operator_out1637_out1            : std_logic;
  SIGNAL Logical_Operator_out1638_out1            : std_logic;
  SIGNAL Logical_Operator_out1639_out1            : std_logic;
  SIGNAL Logical_Operator_out1640_out1            : std_logic;
  SIGNAL Logical_Operator_out1641_out1            : std_logic;
  SIGNAL Logical_Operator_out1642_out1            : std_logic;
  SIGNAL Logical_Operator_out1643_out1            : std_logic;
  SIGNAL Logical_Operator_out1644_out1            : std_logic;
  SIGNAL Logical_Operator_out1645_out1            : std_logic;
  SIGNAL Logical_Operator_out1646_out1            : std_logic;
  SIGNAL Logical_Operator_out1647_out1            : std_logic;
  SIGNAL Logical_Operator_out1648_out1            : std_logic;
  SIGNAL Logical_Operator_out1649_out1            : std_logic;
  SIGNAL Logical_Operator_out1650_out1            : std_logic;
  SIGNAL Logical_Operator_out1651_out1            : std_logic;
  SIGNAL Logical_Operator_out1652_out1            : std_logic;
  SIGNAL Logical_Operator_out1653_out1            : std_logic;
  SIGNAL Logical_Operator_out1654_out1            : std_logic;
  SIGNAL Logical_Operator_out1655_out1            : std_logic;
  SIGNAL Logical_Operator_out1656_out1            : std_logic;
  SIGNAL Logical_Operator_out1657_out1            : std_logic;
  SIGNAL Logical_Operator_out1658_out1            : std_logic;
  SIGNAL Logical_Operator_out1659_out1            : std_logic;
  SIGNAL Logical_Operator_out1660_out1            : std_logic;
  SIGNAL Logical_Operator_out1661_out1            : std_logic;
  SIGNAL Logical_Operator_out1662_out1            : std_logic;
  SIGNAL Logical_Operator_out1663_out1            : std_logic;
  SIGNAL Logical_Operator_out1664_out1            : std_logic;
  SIGNAL Logical_Operator_out1665_out1            : std_logic;
  SIGNAL Logical_Operator_out1666_out1            : std_logic;
  SIGNAL Logical_Operator_out1667_out1            : std_logic;
  SIGNAL Logical_Operator_out1668_out1            : std_logic;
  SIGNAL Logical_Operator_out1669_out1            : std_logic;
  SIGNAL Logical_Operator_out1670_out1            : std_logic;
  SIGNAL Logical_Operator_out1671_out1            : std_logic;
  SIGNAL Logical_Operator_out1672_out1            : std_logic;
  SIGNAL Logical_Operator_out1673_out1            : std_logic;
  SIGNAL Logical_Operator_out1674_out1            : std_logic;
  SIGNAL Logical_Operator_out1675_out1            : std_logic;
  SIGNAL Logical_Operator_out1676_out1            : std_logic;
  SIGNAL Logical_Operator_out1677_out1            : std_logic;
  SIGNAL Logical_Operator_out1678_out1            : std_logic;
  SIGNAL Logical_Operator_out1679_out1            : std_logic;
  SIGNAL Logical_Operator_out1680_out1            : std_logic;
  SIGNAL Logical_Operator_out1681_out1            : std_logic;
  SIGNAL Logical_Operator_out1682_out1            : std_logic;
  SIGNAL Logical_Operator_out1683_out1            : std_logic;
  SIGNAL Logical_Operator_out1684_out1            : std_logic;
  SIGNAL Logical_Operator_out1685_out1            : std_logic;
  SIGNAL Logical_Operator_out1686_out1            : std_logic;
  SIGNAL Logical_Operator_out1687_out1            : std_logic;
  SIGNAL Logical_Operator_out1688_out1            : std_logic;
  SIGNAL Logical_Operator_out1689_out1            : std_logic;
  SIGNAL Logical_Operator_out1690_out1            : std_logic;
  SIGNAL Logical_Operator_out1691_out1            : std_logic;
  SIGNAL Logical_Operator_out1692_out1            : std_logic;
  SIGNAL Logical_Operator_out1693_out1            : std_logic;
  SIGNAL Logical_Operator_out1694_out1            : std_logic;
  SIGNAL Logical_Operator_out1695_out1            : std_logic;
  SIGNAL Logical_Operator_out1696_out1            : std_logic;
  SIGNAL Logical_Operator_out1697_out1            : std_logic;
  SIGNAL Logical_Operator_out1698_out1            : std_logic;
  SIGNAL Logical_Operator_out1699_out1            : std_logic;
  SIGNAL Logical_Operator_out1700_out1            : std_logic;
  SIGNAL Logical_Operator_out1701_out1            : std_logic;
  SIGNAL Logical_Operator_out1702_out1            : std_logic;
  SIGNAL Logical_Operator_out1703_out1            : std_logic;
  SIGNAL Logical_Operator_out1704_out1            : std_logic;
  SIGNAL Logical_Operator_out1705_out1            : std_logic;
  SIGNAL Logical_Operator_out1706_out1            : std_logic;
  SIGNAL Logical_Operator_out1707_out1            : std_logic;
  SIGNAL Logical_Operator_out1708_out1            : std_logic;
  SIGNAL Logical_Operator_out1709_out1            : std_logic;
  SIGNAL Logical_Operator_out1710_out1            : std_logic;
  SIGNAL Logical_Operator_out1711_out1            : std_logic;
  SIGNAL Logical_Operator_out1712_out1            : std_logic;
  SIGNAL Logical_Operator_out1713_out1            : std_logic;
  SIGNAL Logical_Operator_out1714_out1            : std_logic;
  SIGNAL Logical_Operator_out1715_out1            : std_logic;
  SIGNAL Logical_Operator_out1716_out1            : std_logic;
  SIGNAL Logical_Operator_out1717_out1            : std_logic;
  SIGNAL Logical_Operator_out1718_out1            : std_logic;
  SIGNAL Logical_Operator_out1719_out1            : std_logic;
  SIGNAL Logical_Operator_out1720_out1            : std_logic;
  SIGNAL Logical_Operator_out1721_out1            : std_logic;
  SIGNAL Logical_Operator_out1722_out1            : std_logic;
  SIGNAL Logical_Operator_out1723_out1            : std_logic;
  SIGNAL Logical_Operator_out1724_out1            : std_logic;
  SIGNAL Logical_Operator_out1725_out1            : std_logic;
  SIGNAL Logical_Operator_out1726_out1            : std_logic;
  SIGNAL Logical_Operator_out1727_out1            : std_logic;
  SIGNAL Logical_Operator_out1728_out1            : std_logic;
  SIGNAL Logical_Operator_out1729_out1            : std_logic;
  SIGNAL Logical_Operator_out1730_out1            : std_logic;
  SIGNAL Logical_Operator_out1731_out1            : std_logic;
  SIGNAL Logical_Operator_out1732_out1            : std_logic;
  SIGNAL Logical_Operator_out1733_out1            : std_logic;
  SIGNAL Logical_Operator_out1734_out1            : std_logic;
  SIGNAL Logical_Operator_out1735_out1            : std_logic;
  SIGNAL Logical_Operator_out1736_out1            : std_logic;
  SIGNAL Logical_Operator_out1737_out1            : std_logic;
  SIGNAL Logical_Operator_out1738_out1            : std_logic;
  SIGNAL Logical_Operator_out1739_out1            : std_logic;
  SIGNAL Logical_Operator_out1740_out1            : std_logic;
  SIGNAL Logical_Operator_out1741_out1            : std_logic;
  SIGNAL Logical_Operator_out1742_out1            : std_logic;
  SIGNAL Logical_Operator_out1743_out1            : std_logic;
  SIGNAL Logical_Operator_out1744_out1            : std_logic;
  SIGNAL Logical_Operator_out1745_out1            : std_logic;
  SIGNAL Logical_Operator_out1746_out1            : std_logic;
  SIGNAL Logical_Operator_out1747_out1            : std_logic;
  SIGNAL Logical_Operator_out1748_out1            : std_logic;
  SIGNAL Logical_Operator_out1749_out1            : std_logic;
  SIGNAL Logical_Operator_out1750_out1            : std_logic;
  SIGNAL Logical_Operator_out1751_out1            : std_logic;
  SIGNAL Logical_Operator_out1752_out1            : std_logic;
  SIGNAL Logical_Operator_out1753_out1            : std_logic;
  SIGNAL Logical_Operator_out1754_out1            : std_logic;
  SIGNAL Logical_Operator_out1755_out1            : std_logic;
  SIGNAL Logical_Operator_out1756_out1            : std_logic;
  SIGNAL Logical_Operator_out1757_out1            : std_logic;
  SIGNAL Logical_Operator_out1758_out1            : std_logic;
  SIGNAL Logical_Operator_out1759_out1            : std_logic;
  SIGNAL Logical_Operator_out1760_out1            : std_logic;
  SIGNAL Logical_Operator_out1761_out1            : std_logic;
  SIGNAL Logical_Operator_out1762_out1            : std_logic;
  SIGNAL Logical_Operator_out1763_out1            : std_logic;
  SIGNAL Logical_Operator_out1764_out1            : std_logic;
  SIGNAL Logical_Operator_out1765_out1            : std_logic;
  SIGNAL Logical_Operator_out1766_out1            : std_logic;
  SIGNAL Logical_Operator_out1767_out1            : std_logic;
  SIGNAL Logical_Operator_out1768_out1            : std_logic;
  SIGNAL Logical_Operator_out1769_out1            : std_logic;
  SIGNAL Logical_Operator_out1770_out1            : std_logic;
  SIGNAL Logical_Operator_out1771_out1            : std_logic;
  SIGNAL Logical_Operator_out1772_out1            : std_logic;
  SIGNAL Logical_Operator_out1773_out1            : std_logic;
  SIGNAL Logical_Operator_out1774_out1            : std_logic;
  SIGNAL Logical_Operator_out1775_out1            : std_logic;
  SIGNAL Logical_Operator_out1776_out1            : std_logic;
  SIGNAL Logical_Operator_out1777_out1            : std_logic;
  SIGNAL Logical_Operator_out1778_out1            : std_logic;
  SIGNAL Logical_Operator_out1779_out1            : std_logic;
  SIGNAL Logical_Operator_out1780_out1            : std_logic;
  SIGNAL Logical_Operator_out1781_out1            : std_logic;
  SIGNAL Logical_Operator_out1782_out1            : std_logic;
  SIGNAL Logical_Operator_out1783_out1            : std_logic;
  SIGNAL Logical_Operator_out1784_out1            : std_logic;
  SIGNAL Logical_Operator_out1785_out1            : std_logic;
  SIGNAL Logical_Operator_out1786_out1            : std_logic;
  SIGNAL Logical_Operator_out1787_out1            : std_logic;
  SIGNAL Logical_Operator_out1788_out1            : std_logic;
  SIGNAL Logical_Operator_out1789_out1            : std_logic;
  SIGNAL Logical_Operator_out1790_out1            : std_logic;
  SIGNAL Logical_Operator_out1791_out1            : std_logic;
  SIGNAL Logical_Operator_out1792_out1            : std_logic;
  SIGNAL Logical_Operator_out1793_out1            : std_logic;
  SIGNAL Logical_Operator_out1794_out1            : std_logic;
  SIGNAL Logical_Operator_out1795_out1            : std_logic;
  SIGNAL Logical_Operator_out1796_out1            : std_logic;
  SIGNAL Logical_Operator_out1797_out1            : std_logic;
  SIGNAL Logical_Operator_out1798_out1            : std_logic;
  SIGNAL Logical_Operator_out1799_out1            : std_logic;
  SIGNAL Logical_Operator_out1800_out1            : std_logic;
  SIGNAL Logical_Operator_out1801_out1            : std_logic;
  SIGNAL Logical_Operator_out1802_out1            : std_logic;
  SIGNAL Logical_Operator_out1803_out1            : std_logic;
  SIGNAL Logical_Operator_out1804_out1            : std_logic;
  SIGNAL Logical_Operator_out1805_out1            : std_logic;
  SIGNAL Logical_Operator_out1806_out1            : std_logic;
  SIGNAL Logical_Operator_out1807_out1            : std_logic;
  SIGNAL Logical_Operator_out1808_out1            : std_logic;
  SIGNAL Logical_Operator_out1809_out1            : std_logic;
  SIGNAL Logical_Operator_out1810_out1            : std_logic;
  SIGNAL Logical_Operator_out1811_out1            : std_logic;
  SIGNAL Logical_Operator_out1812_out1            : std_logic;
  SIGNAL Logical_Operator_out1813_out1            : std_logic;
  SIGNAL Logical_Operator_out1814_out1            : std_logic;
  SIGNAL Logical_Operator_out1815_out1            : std_logic;
  SIGNAL Logical_Operator_out1816_out1            : std_logic;
  SIGNAL Logical_Operator_out1817_out1            : std_logic;
  SIGNAL Logical_Operator_out1818_out1            : std_logic;
  SIGNAL Logical_Operator_out1819_out1            : std_logic;
  SIGNAL Logical_Operator_out1820_out1            : std_logic;
  SIGNAL Logical_Operator_out1821_out1            : std_logic;
  SIGNAL Logical_Operator_out1822_out1            : std_logic;
  SIGNAL Logical_Operator_out1823_out1            : std_logic;
  SIGNAL Logical_Operator_out1824_out1            : std_logic;
  SIGNAL Logical_Operator_out1825_out1            : std_logic;
  SIGNAL Logical_Operator_out1826_out1            : std_logic;
  SIGNAL Logical_Operator_out1827_out1            : std_logic;
  SIGNAL Logical_Operator_out1828_out1            : std_logic;
  SIGNAL Logical_Operator_out1829_out1            : std_logic;
  SIGNAL Logical_Operator_out1830_out1            : std_logic;
  SIGNAL Logical_Operator_out1831_out1            : std_logic;
  SIGNAL Logical_Operator_out1832_out1            : std_logic;
  SIGNAL Logical_Operator_out1833_out1            : std_logic;
  SIGNAL Logical_Operator_out1834_out1            : std_logic;
  SIGNAL Logical_Operator_out1835_out1            : std_logic;
  SIGNAL Logical_Operator_out1836_out1            : std_logic;
  SIGNAL Logical_Operator_out1837_out1            : std_logic;
  SIGNAL Logical_Operator_out1838_out1            : std_logic;
  SIGNAL Logical_Operator_out1839_out1            : std_logic;
  SIGNAL Logical_Operator_out1840_out1            : std_logic;
  SIGNAL Logical_Operator_out1841_out1            : std_logic;
  SIGNAL Logical_Operator_out1842_out1            : std_logic;
  SIGNAL Logical_Operator_out1843_out1            : std_logic;
  SIGNAL Logical_Operator_out1844_out1            : std_logic;
  SIGNAL Logical_Operator_out1845_out1            : std_logic;
  SIGNAL Logical_Operator_out1846_out1            : std_logic;
  SIGNAL Logical_Operator_out1847_out1            : std_logic;
  SIGNAL Logical_Operator_out1848_out1            : std_logic;
  SIGNAL Logical_Operator_out1849_out1            : std_logic;
  SIGNAL Logical_Operator_out1850_out1            : std_logic;
  SIGNAL Logical_Operator_out1851_out1            : std_logic;
  SIGNAL Logical_Operator_out1852_out1            : std_logic;
  SIGNAL Logical_Operator_out1853_out1            : std_logic;
  SIGNAL Logical_Operator_out1854_out1            : std_logic;
  SIGNAL Logical_Operator_out1855_out1            : std_logic;
  SIGNAL Logical_Operator_out1856_out1            : std_logic;
  SIGNAL Logical_Operator_out1857_out1            : std_logic;
  SIGNAL Logical_Operator_out1858_out1            : std_logic;
  SIGNAL Logical_Operator_out1859_out1            : std_logic;
  SIGNAL Logical_Operator_out1860_out1            : std_logic;
  SIGNAL Logical_Operator_out1861_out1            : std_logic;
  SIGNAL Logical_Operator_out1862_out1            : std_logic;
  SIGNAL Logical_Operator_out1863_out1            : std_logic;
  SIGNAL Logical_Operator_out1864_out1            : std_logic;
  SIGNAL Logical_Operator_out1865_out1            : std_logic;
  SIGNAL Logical_Operator_out1866_out1            : std_logic;
  SIGNAL Logical_Operator_out1867_out1            : std_logic;
  SIGNAL Logical_Operator_out1868_out1            : std_logic;
  SIGNAL Logical_Operator_out1869_out1            : std_logic;
  SIGNAL Logical_Operator_out1870_out1            : std_logic;
  SIGNAL Logical_Operator_out1871_out1            : std_logic;
  SIGNAL Logical_Operator_out1872_out1            : std_logic;
  SIGNAL Logical_Operator_out1873_out1            : std_logic;
  SIGNAL Logical_Operator_out1874_out1            : std_logic;
  SIGNAL Logical_Operator_out1875_out1            : std_logic;
  SIGNAL Logical_Operator_out1876_out1            : std_logic;
  SIGNAL Logical_Operator_out1877_out1            : std_logic;
  SIGNAL Logical_Operator_out1878_out1            : std_logic;
  SIGNAL Logical_Operator_out1879_out1            : std_logic;
  SIGNAL Logical_Operator_out1880_out1            : std_logic;
  SIGNAL Logical_Operator_out1881_out1            : std_logic;
  SIGNAL Logical_Operator_out1882_out1            : std_logic;
  SIGNAL Logical_Operator_out1883_out1            : std_logic;
  SIGNAL Logical_Operator_out1884_out1            : std_logic;
  SIGNAL Logical_Operator_out1885_out1            : std_logic;
  SIGNAL Logical_Operator_out1886_out1            : std_logic;
  SIGNAL Logical_Operator_out1887_out1            : std_logic;
  SIGNAL Logical_Operator_out1888_out1            : std_logic;
  SIGNAL Logical_Operator_out1889_out1            : std_logic;
  SIGNAL Logical_Operator_out1890_out1            : std_logic;
  SIGNAL Logical_Operator_out1891_out1            : std_logic;
  SIGNAL Logical_Operator_out1892_out1            : std_logic;
  SIGNAL Logical_Operator_out1893_out1            : std_logic;
  SIGNAL Logical_Operator_out1894_out1            : std_logic;
  SIGNAL Logical_Operator_out1895_out1            : std_logic;
  SIGNAL Logical_Operator_out1896_out1            : std_logic;
  SIGNAL Logical_Operator_out1897_out1            : std_logic;
  SIGNAL Logical_Operator_out1898_out1            : std_logic;
  SIGNAL Logical_Operator_out1899_out1            : std_logic;
  SIGNAL Logical_Operator_out1900_out1            : std_logic;
  SIGNAL Logical_Operator_out1901_out1            : std_logic;
  SIGNAL Logical_Operator_out1902_out1            : std_logic;
  SIGNAL Logical_Operator_out1903_out1            : std_logic;
  SIGNAL Logical_Operator_out1904_out1            : std_logic;
  SIGNAL Logical_Operator_out1905_out1            : std_logic;
  SIGNAL Logical_Operator_out1906_out1            : std_logic;
  SIGNAL Logical_Operator_out1907_out1            : std_logic;
  SIGNAL Logical_Operator_out1908_out1            : std_logic;
  SIGNAL Logical_Operator_out1909_out1            : std_logic;
  SIGNAL Logical_Operator_out1910_out1            : std_logic;
  SIGNAL Logical_Operator_out1911_out1            : std_logic;
  SIGNAL Logical_Operator_out1912_out1            : std_logic;
  SIGNAL Logical_Operator_out1913_out1            : std_logic;
  SIGNAL Logical_Operator_out1914_out1            : std_logic;
  SIGNAL Logical_Operator_out1915_out1            : std_logic;
  SIGNAL Logical_Operator_out1916_out1            : std_logic;
  SIGNAL Logical_Operator_out1917_out1            : std_logic;
  SIGNAL Logical_Operator_out1918_out1            : std_logic;
  SIGNAL Logical_Operator_out1919_out1            : std_logic;
  SIGNAL Logical_Operator_out1920_out1            : std_logic;
  SIGNAL Logical_Operator_out1921_out1            : std_logic;
  SIGNAL Logical_Operator_out1922_out1            : std_logic;
  SIGNAL Logical_Operator_out1923_out1            : std_logic;
  SIGNAL Logical_Operator_out1924_out1            : std_logic;
  SIGNAL Logical_Operator_out1925_out1            : std_logic;
  SIGNAL Logical_Operator_out1926_out1            : std_logic;
  SIGNAL Logical_Operator_out1927_out1            : std_logic;
  SIGNAL Logical_Operator_out1928_out1            : std_logic;
  SIGNAL Logical_Operator_out1929_out1            : std_logic;
  SIGNAL Logical_Operator_out1930_out1            : std_logic;
  SIGNAL Logical_Operator_out1931_out1            : std_logic;
  SIGNAL Logical_Operator_out1932_out1            : std_logic;
  SIGNAL Logical_Operator_out1933_out1            : std_logic;
  SIGNAL Logical_Operator_out1934_out1            : std_logic;
  SIGNAL Logical_Operator_out1935_out1            : std_logic;
  SIGNAL Logical_Operator_out1936_out1            : std_logic;
  SIGNAL Logical_Operator_out1937_out1            : std_logic;
  SIGNAL Logical_Operator_out1938_out1            : std_logic;
  SIGNAL Logical_Operator_out1939_out1            : std_logic;
  SIGNAL Logical_Operator_out1940_out1            : std_logic;
  SIGNAL Logical_Operator_out1941_out1            : std_logic;
  SIGNAL Logical_Operator_out1942_out1            : std_logic;
  SIGNAL Logical_Operator_out1943_out1            : std_logic;
  SIGNAL Logical_Operator_out1944_out1            : std_logic;
  SIGNAL Logical_Operator_out1945_out1            : std_logic;
  SIGNAL Logical_Operator_out1946_out1            : std_logic;
  SIGNAL Logical_Operator_out1947_out1            : std_logic;
  SIGNAL Logical_Operator_out1948_out1            : std_logic;
  SIGNAL Logical_Operator_out1949_out1            : std_logic;
  SIGNAL Logical_Operator_out1950_out1            : std_logic;
  SIGNAL Logical_Operator_out1951_out1            : std_logic;
  SIGNAL Logical_Operator_out1952_out1            : std_logic;
  SIGNAL Logical_Operator_out1953_out1            : std_logic;
  SIGNAL Logical_Operator_out1954_out1            : std_logic;
  SIGNAL Logical_Operator_out1955_out1            : std_logic;
  SIGNAL Logical_Operator_out1956_out1            : std_logic;
  SIGNAL Logical_Operator_out1957_out1            : std_logic;
  SIGNAL Logical_Operator_out1958_out1            : std_logic;
  SIGNAL Logical_Operator_out1959_out1            : std_logic;
  SIGNAL Logical_Operator_out1960_out1            : std_logic;
  SIGNAL Logical_Operator_out1961_out1            : std_logic;
  SIGNAL Logical_Operator_out1962_out1            : std_logic;
  SIGNAL Logical_Operator_out1963_out1            : std_logic;
  SIGNAL Logical_Operator_out1964_out1            : std_logic;
  SIGNAL Logical_Operator_out1965_out1            : std_logic;
  SIGNAL Logical_Operator_out1966_out1            : std_logic;
  SIGNAL Logical_Operator_out1967_out1            : std_logic;
  SIGNAL Logical_Operator_out1968_out1            : std_logic;
  SIGNAL Logical_Operator_out1969_out1            : std_logic;
  SIGNAL Logical_Operator_out1970_out1            : std_logic;
  SIGNAL Logical_Operator_out1971_out1            : std_logic;
  SIGNAL Logical_Operator_out1972_out1            : std_logic;
  SIGNAL Logical_Operator_out1973_out1            : std_logic;
  SIGNAL Logical_Operator_out1974_out1            : std_logic;
  SIGNAL Logical_Operator_out1975_out1            : std_logic;
  SIGNAL Logical_Operator_out1976_out1            : std_logic;
  SIGNAL Logical_Operator_out1977_out1            : std_logic;
  SIGNAL Logical_Operator_out1978_out1            : std_logic;
  SIGNAL Logical_Operator_out1979_out1            : std_logic;
  SIGNAL Logical_Operator_out1980_out1            : std_logic;
  SIGNAL Logical_Operator_out1981_out1            : std_logic;
  SIGNAL Logical_Operator_out1982_out1            : std_logic;
  SIGNAL Logical_Operator_out1983_out1            : std_logic;
  SIGNAL Logical_Operator_out1984_out1            : std_logic;
  SIGNAL Logical_Operator_out1985_out1            : std_logic;
  SIGNAL Logical_Operator_out1986_out1            : std_logic;
  SIGNAL Logical_Operator_out1987_out1            : std_logic;
  SIGNAL Logical_Operator_out1988_out1            : std_logic;
  SIGNAL Logical_Operator_out1989_out1            : std_logic;
  SIGNAL Logical_Operator_out1990_out1            : std_logic;
  SIGNAL Logical_Operator_out1991_out1            : std_logic;
  SIGNAL Logical_Operator_out1992_out1            : std_logic;
  SIGNAL Logical_Operator_out1993_out1            : std_logic;
  SIGNAL Logical_Operator_out1994_out1            : std_logic;
  SIGNAL Logical_Operator_out1995_out1            : std_logic;
  SIGNAL Logical_Operator_out1996_out1            : std_logic;
  SIGNAL Logical_Operator_out1997_out1            : std_logic;
  SIGNAL Logical_Operator_out1998_out1            : std_logic;
  SIGNAL Logical_Operator_out1999_out1            : std_logic;
  SIGNAL Logical_Operator_out2000_out1            : std_logic;
  SIGNAL Logical_Operator_out2001_out1            : std_logic;
  SIGNAL Logical_Operator_out2002_out1            : std_logic;
  SIGNAL Logical_Operator_out2003_out1            : std_logic;
  SIGNAL Logical_Operator_out2004_out1            : std_logic;
  SIGNAL Logical_Operator_out2005_out1            : std_logic;
  SIGNAL Logical_Operator_out2006_out1            : std_logic;
  SIGNAL Logical_Operator_out2007_out1            : std_logic;
  SIGNAL Logical_Operator_out2008_out1            : std_logic;
  SIGNAL Logical_Operator_out2009_out1            : std_logic;
  SIGNAL Logical_Operator_out2010_out1            : std_logic;
  SIGNAL Logical_Operator_out2011_out1            : std_logic;
  SIGNAL Logical_Operator_out2012_out1            : std_logic;
  SIGNAL Logical_Operator_out2013_out1            : std_logic;
  SIGNAL Logical_Operator_out2014_out1            : std_logic;
  SIGNAL Logical_Operator_out2015_out1            : std_logic;
  SIGNAL Logical_Operator_out2016_out1            : std_logic;
  SIGNAL Logical_Operator_out2017_out1            : std_logic;
  SIGNAL Logical_Operator_out2018_out1            : std_logic;
  SIGNAL Logical_Operator_out2019_out1            : std_logic;
  SIGNAL Logical_Operator_out2020_out1            : std_logic;
  SIGNAL Logical_Operator_out2021_out1            : std_logic;
  SIGNAL Logical_Operator_out2022_out1            : std_logic;
  SIGNAL Logical_Operator_out2023_out1            : std_logic;
  SIGNAL Logical_Operator_out2024_out1            : std_logic;
  SIGNAL Logical_Operator_out2025_out1            : std_logic;
  SIGNAL Logical_Operator_out2026_out1            : std_logic;
  SIGNAL Logical_Operator_out2027_out1            : std_logic;
  SIGNAL Logical_Operator_out2028_out1            : std_logic;
  SIGNAL Logical_Operator_out2029_out1            : std_logic;
  SIGNAL Logical_Operator_out2030_out1            : std_logic;
  SIGNAL Logical_Operator_out2031_out1            : std_logic;
  SIGNAL Logical_Operator_out2032_out1            : std_logic;
  SIGNAL Logical_Operator_out2033_out1            : std_logic;
  SIGNAL Logical_Operator_out2034_out1            : std_logic;
  SIGNAL Logical_Operator_out2035_out1            : std_logic;
  SIGNAL Logical_Operator_out2036_out1            : std_logic;
  SIGNAL Logical_Operator_out2037_out1            : std_logic;
  SIGNAL Logical_Operator_out2038_out1            : std_logic;
  SIGNAL Logical_Operator_out2039_out1            : std_logic;
  SIGNAL Logical_Operator_out2040_out1            : std_logic;
  SIGNAL Logical_Operator_out2041_out1            : std_logic;
  SIGNAL Logical_Operator_out2042_out1            : std_logic;
  SIGNAL Logical_Operator_out2043_out1            : std_logic;
  SIGNAL Logical_Operator_out2044_out1            : std_logic;
  SIGNAL Logical_Operator_out2045_out1            : std_logic;
  SIGNAL Logical_Operator_out2046_out1            : std_logic;
  SIGNAL Logical_Operator_out2047_out1            : std_logic;
  SIGNAL Logical_Operator_out2048_out1            : std_logic;
  SIGNAL Logical_Operator_out2049_out1            : std_logic;
  SIGNAL Logical_Operator_out2050_out1            : std_logic;
  SIGNAL Logical_Operator_out2051_out1            : std_logic;
  SIGNAL Logical_Operator_out2052_out1            : std_logic;
  SIGNAL Logical_Operator_out2053_out1            : std_logic;
  SIGNAL Logical_Operator_out2054_out1            : std_logic;
  SIGNAL Logical_Operator_out2055_out1            : std_logic;
  SIGNAL Logical_Operator_out2056_out1            : std_logic;
  SIGNAL Logical_Operator_out2057_out1            : std_logic;
  SIGNAL Logical_Operator_out2058_out1            : std_logic;
  SIGNAL Logical_Operator_out2059_out1            : std_logic;
  SIGNAL Logical_Operator_out2060_out1            : std_logic;
  SIGNAL Logical_Operator_out2061_out1            : std_logic;
  SIGNAL Logical_Operator_out2062_out1            : std_logic;
  SIGNAL Logical_Operator_out2063_out1            : std_logic;
  SIGNAL Logical_Operator_out2064_out1            : std_logic;
  SIGNAL Logical_Operator_out2065_out1            : std_logic;
  SIGNAL Logical_Operator_out2066_out1            : std_logic;
  SIGNAL Logical_Operator_out2067_out1            : std_logic;
  SIGNAL Logical_Operator_out2068_out1            : std_logic;
  SIGNAL Logical_Operator_out2069_out1            : std_logic;
  SIGNAL Logical_Operator_out2070_out1            : std_logic;
  SIGNAL Logical_Operator_out2071_out1            : std_logic;
  SIGNAL Logical_Operator_out2072_out1            : std_logic;
  SIGNAL Logical_Operator_out2073_out1            : std_logic;
  SIGNAL Logical_Operator_out2074_out1            : std_logic;
  SIGNAL Logical_Operator_out2075_out1            : std_logic;
  SIGNAL Logical_Operator_out2076_out1            : std_logic;
  SIGNAL Logical_Operator_out2077_out1            : std_logic;
  SIGNAL Logical_Operator_out2078_out1            : std_logic;
  SIGNAL Logical_Operator_out2079_out1            : std_logic;
  SIGNAL Logical_Operator_out2080_out1            : std_logic;
  SIGNAL Logical_Operator_out2081_out1            : std_logic;
  SIGNAL Logical_Operator_out2082_out1            : std_logic;
  SIGNAL Logical_Operator_out2083_out1            : std_logic;
  SIGNAL Logical_Operator_out2084_out1            : std_logic;
  SIGNAL Logical_Operator_out2085_out1            : std_logic;
  SIGNAL Logical_Operator_out2086_out1            : std_logic;
  SIGNAL Logical_Operator_out2087_out1            : std_logic;
  SIGNAL Logical_Operator_out2088_out1            : std_logic;
  SIGNAL Logical_Operator_out2089_out1            : std_logic;
  SIGNAL Logical_Operator_out2090_out1            : std_logic;
  SIGNAL Logical_Operator_out2091_out1            : std_logic;
  SIGNAL Logical_Operator_out2092_out1            : std_logic;
  SIGNAL Logical_Operator_out2093_out1            : std_logic;
  SIGNAL Logical_Operator_out2094_out1            : std_logic;
  SIGNAL Logical_Operator_out2095_out1            : std_logic;
  SIGNAL Logical_Operator_out2096_out1            : std_logic;
  SIGNAL Logical_Operator_out2097_out1            : std_logic;
  SIGNAL Logical_Operator_out2098_out1            : std_logic;
  SIGNAL Logical_Operator_out2099_out1            : std_logic;
  SIGNAL Logical_Operator_out2100_out1            : std_logic;
  SIGNAL Logical_Operator_out2101_out1            : std_logic;
  SIGNAL Logical_Operator_out2102_out1            : std_logic;
  SIGNAL Logical_Operator_out2103_out1            : std_logic;
  SIGNAL Logical_Operator_out2104_out1            : std_logic;
  SIGNAL Logical_Operator_out2105_out1            : std_logic;
  SIGNAL Logical_Operator_out2106_out1            : std_logic;
  SIGNAL Logical_Operator_out2107_out1            : std_logic;
  SIGNAL Logical_Operator_out2108_out1            : std_logic;
  SIGNAL Logical_Operator_out2109_out1            : std_logic;
  SIGNAL Logical_Operator_out2110_out1            : std_logic;
  SIGNAL Logical_Operator_out2111_out1            : std_logic;
  SIGNAL Logical_Operator_out2112_out1            : std_logic;
  SIGNAL Logical_Operator_out2113_out1            : std_logic;
  SIGNAL Logical_Operator_out2114_out1            : std_logic;
  SIGNAL Logical_Operator_out2115_out1            : std_logic;
  SIGNAL Logical_Operator_out2116_out1            : std_logic;
  SIGNAL Logical_Operator_out2117_out1            : std_logic;
  SIGNAL Logical_Operator_out2118_out1            : std_logic;
  SIGNAL Logical_Operator_out2119_out1            : std_logic;
  SIGNAL Logical_Operator_out2120_out1            : std_logic;
  SIGNAL Logical_Operator_out2121_out1            : std_logic;
  SIGNAL Logical_Operator_out2122_out1            : std_logic;
  SIGNAL Logical_Operator_out2123_out1            : std_logic;
  SIGNAL Logical_Operator_out2124_out1            : std_logic;
  SIGNAL Logical_Operator_out2125_out1            : std_logic;
  SIGNAL Logical_Operator_out2126_out1            : std_logic;
  SIGNAL Logical_Operator_out2127_out1            : std_logic;
  SIGNAL Logical_Operator_out2128_out1            : std_logic;
  SIGNAL Logical_Operator_out2129_out1            : std_logic;
  SIGNAL Logical_Operator_out2130_out1            : std_logic;
  SIGNAL Logical_Operator_out2131_out1            : std_logic;
  SIGNAL Logical_Operator_out2132_out1            : std_logic;
  SIGNAL Logical_Operator_out2133_out1            : std_logic;
  SIGNAL Logical_Operator_out2134_out1            : std_logic;
  SIGNAL Logical_Operator_out2135_out1            : std_logic;
  SIGNAL Logical_Operator_out2136_out1            : std_logic;
  SIGNAL Logical_Operator_out2137_out1            : std_logic;
  SIGNAL Logical_Operator_out2138_out1            : std_logic;
  SIGNAL Logical_Operator_out2139_out1            : std_logic;
  SIGNAL Logical_Operator_out2140_out1            : std_logic;
  SIGNAL Logical_Operator_out2141_out1            : std_logic;
  SIGNAL Logical_Operator_out2142_out1            : std_logic;
  SIGNAL Logical_Operator_out2143_out1            : std_logic;
  SIGNAL Logical_Operator_out2144_out1            : std_logic;
  SIGNAL Logical_Operator_out2145_out1            : std_logic;
  SIGNAL Logical_Operator_out2146_out1            : std_logic;
  SIGNAL Logical_Operator_out2147_out1            : std_logic;
  SIGNAL Logical_Operator_out2148_out1            : std_logic;
  SIGNAL Logical_Operator_out2149_out1            : std_logic;
  SIGNAL Logical_Operator_out2150_out1            : std_logic;
  SIGNAL Logical_Operator_out2151_out1            : std_logic;
  SIGNAL Logical_Operator_out2152_out1            : std_logic;
  SIGNAL Logical_Operator_out2153_out1            : std_logic;
  SIGNAL Logical_Operator_out2154_out1            : std_logic;
  SIGNAL Logical_Operator_out2155_out1            : std_logic;
  SIGNAL Logical_Operator_out2156_out1            : std_logic;
  SIGNAL Logical_Operator_out2157_out1            : std_logic;
  SIGNAL Logical_Operator_out2158_out1            : std_logic;
  SIGNAL Logical_Operator_out2159_out1            : std_logic;
  SIGNAL Logical_Operator_out2160_out1            : std_logic;
  SIGNAL Logical_Operator_out2161_out1            : std_logic;
  SIGNAL Logical_Operator_out2162_out1            : std_logic;
  SIGNAL Logical_Operator_out2163_out1            : std_logic;
  SIGNAL Logical_Operator_out2164_out1            : std_logic;
  SIGNAL Logical_Operator_out2165_out1            : std_logic;
  SIGNAL Logical_Operator_out2166_out1            : std_logic;
  SIGNAL Logical_Operator_out2167_out1            : std_logic;
  SIGNAL Logical_Operator_out2168_out1            : std_logic;
  SIGNAL Logical_Operator_out2169_out1            : std_logic;
  SIGNAL Logical_Operator_out2170_out1            : std_logic;
  SIGNAL Logical_Operator_out2171_out1            : std_logic;
  SIGNAL Logical_Operator_out2172_out1            : std_logic;
  SIGNAL Logical_Operator_out2173_out1            : std_logic;
  SIGNAL Logical_Operator_out2174_out1            : std_logic;
  SIGNAL Logical_Operator_out2175_out1            : std_logic;
  SIGNAL Logical_Operator_out2176_out1            : std_logic;
  SIGNAL Logical_Operator_out2177_out1            : std_logic;
  SIGNAL Logical_Operator_out2178_out1            : std_logic;
  SIGNAL Logical_Operator_out2179_out1            : std_logic;
  SIGNAL Logical_Operator_out2180_out1            : std_logic;
  SIGNAL Logical_Operator_out2181_out1            : std_logic;
  SIGNAL Logical_Operator_out2182_out1            : std_logic;
  SIGNAL Logical_Operator_out2183_out1            : std_logic;
  SIGNAL Logical_Operator_out2184_out1            : std_logic;
  SIGNAL Logical_Operator_out2185_out1            : std_logic;
  SIGNAL Logical_Operator_out2186_out1            : std_logic;
  SIGNAL Logical_Operator_out2187_out1            : std_logic;
  SIGNAL Logical_Operator_out2188_out1            : std_logic;
  SIGNAL Logical_Operator_out2189_out1            : std_logic;
  SIGNAL Logical_Operator_out2190_out1            : std_logic;
  SIGNAL Logical_Operator_out2191_out1            : std_logic;
  SIGNAL Logical_Operator_out2192_out1            : std_logic;
  SIGNAL Logical_Operator_out2193_out1            : std_logic;
  SIGNAL Logical_Operator_out2194_out1            : std_logic;
  SIGNAL Logical_Operator_out2195_out1            : std_logic;
  SIGNAL Logical_Operator_out2196_out1            : std_logic;
  SIGNAL Logical_Operator_out2197_out1            : std_logic;
  SIGNAL Logical_Operator_out2198_out1            : std_logic;
  SIGNAL Logical_Operator_out2199_out1            : std_logic;
  SIGNAL Logical_Operator_out2200_out1            : std_logic;
  SIGNAL Logical_Operator_out2201_out1            : std_logic;
  SIGNAL Logical_Operator_out2202_out1            : std_logic;
  SIGNAL Logical_Operator_out2203_out1            : std_logic;
  SIGNAL Logical_Operator_out2204_out1            : std_logic;
  SIGNAL Logical_Operator_out2205_out1            : std_logic;
  SIGNAL Logical_Operator_out2206_out1            : std_logic;
  SIGNAL Logical_Operator_out2207_out1            : std_logic;
  SIGNAL Logical_Operator_out2208_out1            : std_logic;
  SIGNAL Logical_Operator_out2209_out1            : std_logic;
  SIGNAL Logical_Operator_out2210_out1            : std_logic;
  SIGNAL Logical_Operator_out2211_out1            : std_logic;
  SIGNAL Logical_Operator_out2212_out1            : std_logic;
  SIGNAL Logical_Operator_out2213_out1            : std_logic;
  SIGNAL Logical_Operator_out2214_out1            : std_logic;
  SIGNAL Logical_Operator_out2215_out1            : std_logic;
  SIGNAL Logical_Operator_out2216_out1            : std_logic;
  SIGNAL Logical_Operator_out2217_out1            : std_logic;
  SIGNAL Logical_Operator_out2218_out1            : std_logic;
  SIGNAL Logical_Operator_out2219_out1            : std_logic;
  SIGNAL Logical_Operator_out2220_out1            : std_logic;
  SIGNAL Logical_Operator_out2221_out1            : std_logic;
  SIGNAL Logical_Operator_out2222_out1            : std_logic;
  SIGNAL Logical_Operator_out2223_out1            : std_logic;
  SIGNAL Logical_Operator_out2224_out1            : std_logic;
  SIGNAL Logical_Operator_out2225_out1            : std_logic;
  SIGNAL Logical_Operator_out2226_out1            : std_logic;
  SIGNAL Logical_Operator_out2227_out1            : std_logic;
  SIGNAL Logical_Operator_out2228_out1            : std_logic;
  SIGNAL Logical_Operator_out2229_out1            : std_logic;
  SIGNAL Logical_Operator_out2230_out1            : std_logic;
  SIGNAL Logical_Operator_out2231_out1            : std_logic;
  SIGNAL Logical_Operator_out2232_out1            : std_logic;
  SIGNAL Logical_Operator_out2233_out1            : std_logic;
  SIGNAL Logical_Operator_out2234_out1            : std_logic;
  SIGNAL Logical_Operator_out2235_out1            : std_logic;
  SIGNAL Logical_Operator_out2236_out1            : std_logic;
  SIGNAL Logical_Operator_out2237_out1            : std_logic;
  SIGNAL Logical_Operator_out2238_out1            : std_logic;
  SIGNAL Logical_Operator_out2239_out1            : std_logic;
  SIGNAL Logical_Operator_out2240_out1            : std_logic;
  SIGNAL Logical_Operator_out2241_out1            : std_logic;
  SIGNAL Logical_Operator_out2242_out1            : std_logic;
  SIGNAL Logical_Operator_out2243_out1            : std_logic;
  SIGNAL Logical_Operator_out2244_out1            : std_logic;
  SIGNAL Logical_Operator_out2245_out1            : std_logic;
  SIGNAL Logical_Operator_out2246_out1            : std_logic;
  SIGNAL Logical_Operator_out2247_out1            : std_logic;
  SIGNAL Logical_Operator_out2248_out1            : std_logic;
  SIGNAL Logical_Operator_out2249_out1            : std_logic;
  SIGNAL Logical_Operator_out2250_out1            : std_logic;
  SIGNAL Logical_Operator_out2251_out1            : std_logic;
  SIGNAL Logical_Operator_out2252_out1            : std_logic;
  SIGNAL Logical_Operator_out2253_out1            : std_logic;
  SIGNAL Logical_Operator_out2254_out1            : std_logic;
  SIGNAL Logical_Operator_out2255_out1            : std_logic;
  SIGNAL Logical_Operator_out2256_out1            : std_logic;
  SIGNAL Logical_Operator_out2257_out1            : std_logic;
  SIGNAL Logical_Operator_out2258_out1            : std_logic;
  SIGNAL Logical_Operator_out2259_out1            : std_logic;
  SIGNAL Logical_Operator_out2260_out1            : std_logic;
  SIGNAL Logical_Operator_out2261_out1            : std_logic;
  SIGNAL Logical_Operator_out2262_out1            : std_logic;
  SIGNAL Logical_Operator_out2263_out1            : std_logic;
  SIGNAL Logical_Operator_out2264_out1            : std_logic;
  SIGNAL Logical_Operator_out2265_out1            : std_logic;
  SIGNAL Logical_Operator_out2266_out1            : std_logic;
  SIGNAL Logical_Operator_out2267_out1            : std_logic;
  SIGNAL Logical_Operator_out2268_out1            : std_logic;
  SIGNAL Logical_Operator_out2269_out1            : std_logic;
  SIGNAL Logical_Operator_out2270_out1            : std_logic;
  SIGNAL Logical_Operator_out2271_out1            : std_logic;
  SIGNAL Logical_Operator_out2272_out1            : std_logic;
  SIGNAL Logical_Operator_out2273_out1            : std_logic;
  SIGNAL Logical_Operator_out2274_out1            : std_logic;
  SIGNAL Logical_Operator_out2275_out1            : std_logic;
  SIGNAL Logical_Operator_out2276_out1            : std_logic;
  SIGNAL Logical_Operator_out2277_out1            : std_logic;
  SIGNAL Logical_Operator_out2278_out1            : std_logic;
  SIGNAL Logical_Operator_out2279_out1            : std_logic;
  SIGNAL Logical_Operator_out2280_out1            : std_logic;
  SIGNAL Logical_Operator_out2281_out1            : std_logic;
  SIGNAL Logical_Operator_out2282_out1            : std_logic;
  SIGNAL Logical_Operator_out2283_out1            : std_logic;
  SIGNAL Logical_Operator_out2284_out1            : std_logic;
  SIGNAL Logical_Operator_out2285_out1            : std_logic;
  SIGNAL Logical_Operator_out2286_out1            : std_logic;
  SIGNAL Logical_Operator_out2287_out1            : std_logic;
  SIGNAL Logical_Operator_out2288_out1            : std_logic;
  SIGNAL Logical_Operator_out2289_out1            : std_logic;
  SIGNAL Logical_Operator_out2290_out1            : std_logic;
  SIGNAL Logical_Operator_out2291_out1            : std_logic;
  SIGNAL Logical_Operator_out2292_out1            : std_logic;
  SIGNAL Logical_Operator_out2293_out1            : std_logic;
  SIGNAL Logical_Operator_out2294_out1            : std_logic;
  SIGNAL Logical_Operator_out2295_out1            : std_logic;
  SIGNAL Logical_Operator_out2296_out1            : std_logic;
  SIGNAL Logical_Operator_out2297_out1            : std_logic;
  SIGNAL Logical_Operator_out2298_out1            : std_logic;
  SIGNAL Logical_Operator_out2299_out1            : std_logic;
  SIGNAL Logical_Operator_out2300_out1            : std_logic;
  SIGNAL Logical_Operator_out2301_out1            : std_logic;
  SIGNAL Logical_Operator_out2302_out1            : std_logic;
  SIGNAL Logical_Operator_out2303_out1            : std_logic;
  SIGNAL Logical_Operator_out2304_out1            : std_logic;
  SIGNAL Logical_Operator_out2305_out1            : std_logic;
  SIGNAL Logical_Operator_out2306_out1            : std_logic;
  SIGNAL Logical_Operator_out2307_out1            : std_logic;
  SIGNAL Logical_Operator_out2308_out1            : std_logic;
  SIGNAL Logical_Operator_out2309_out1            : std_logic;
  SIGNAL Logical_Operator_out2310_out1            : std_logic;
  SIGNAL Logical_Operator_out2311_out1            : std_logic;
  SIGNAL Logical_Operator_out2312_out1            : std_logic;
  SIGNAL Logical_Operator_out2313_out1            : std_logic;
  SIGNAL Logical_Operator_out2314_out1            : std_logic;
  SIGNAL Logical_Operator_out2315_out1            : std_logic;
  SIGNAL Logical_Operator_out2316_out1            : std_logic;
  SIGNAL Logical_Operator_out2317_out1            : std_logic;
  SIGNAL Logical_Operator_out2318_out1            : std_logic;
  SIGNAL Logical_Operator_out2319_out1            : std_logic;
  SIGNAL Logical_Operator_out2320_out1            : std_logic;
  SIGNAL Logical_Operator_out2321_out1            : std_logic;
  SIGNAL Logical_Operator_out2322_out1            : std_logic;
  SIGNAL Logical_Operator_out2323_out1            : std_logic;
  SIGNAL Logical_Operator_out2324_out1            : std_logic;
  SIGNAL Logical_Operator_out2325_out1            : std_logic;
  SIGNAL Logical_Operator_out2326_out1            : std_logic;
  SIGNAL Logical_Operator_out2327_out1            : std_logic;
  SIGNAL Logical_Operator_out2328_out1            : std_logic;
  SIGNAL Logical_Operator_out2329_out1            : std_logic;
  SIGNAL Logical_Operator_out2330_out1            : std_logic;
  SIGNAL Logical_Operator_out2331_out1            : std_logic;
  SIGNAL Logical_Operator_out2332_out1            : std_logic;
  SIGNAL Logical_Operator_out2333_out1            : std_logic;
  SIGNAL Logical_Operator_out2334_out1            : std_logic;
  SIGNAL Logical_Operator_out2335_out1            : std_logic;
  SIGNAL Logical_Operator_out2336_out1            : std_logic;
  SIGNAL Logical_Operator_out2337_out1            : std_logic;
  SIGNAL Logical_Operator_out2338_out1            : std_logic;
  SIGNAL Logical_Operator_out2339_out1            : std_logic;
  SIGNAL Logical_Operator_out2340_out1            : std_logic;
  SIGNAL Logical_Operator_out2341_out1            : std_logic;
  SIGNAL Logical_Operator_out2342_out1            : std_logic;
  SIGNAL Logical_Operator_out2343_out1            : std_logic;
  SIGNAL Logical_Operator_out2344_out1            : std_logic;
  SIGNAL Logical_Operator_out2345_out1            : std_logic;
  SIGNAL Logical_Operator_out2346_out1            : std_logic;
  SIGNAL Logical_Operator_out2347_out1            : std_logic;
  SIGNAL Logical_Operator_out2348_out1            : std_logic;
  SIGNAL Logical_Operator_out2349_out1            : std_logic;
  SIGNAL Logical_Operator_out2350_out1            : std_logic;
  SIGNAL Logical_Operator_out2351_out1            : std_logic;
  SIGNAL Logical_Operator_out2352_out1            : std_logic;
  SIGNAL Logical_Operator_out2353_out1            : std_logic;
  SIGNAL Logical_Operator_out2354_out1            : std_logic;
  SIGNAL Logical_Operator_out2355_out1            : std_logic;
  SIGNAL Logical_Operator_out2356_out1            : std_logic;
  SIGNAL Logical_Operator_out2357_out1            : std_logic;
  SIGNAL Logical_Operator_out2358_out1            : std_logic;
  SIGNAL Logical_Operator_out2359_out1            : std_logic;
  SIGNAL Logical_Operator_out2360_out1            : std_logic;
  SIGNAL Logical_Operator_out2361_out1            : std_logic;
  SIGNAL Logical_Operator_out2362_out1            : std_logic;
  SIGNAL Logical_Operator_out2363_out1            : std_logic;
  SIGNAL Logical_Operator_out2364_out1            : std_logic;
  SIGNAL Logical_Operator_out2365_out1            : std_logic;
  SIGNAL Logical_Operator_out2366_out1            : std_logic;
  SIGNAL Logical_Operator_out2367_out1            : std_logic;
  SIGNAL Logical_Operator_out2368_out1            : std_logic;
  SIGNAL Logical_Operator_out2369_out1            : std_logic;
  SIGNAL Logical_Operator_out2370_out1            : std_logic;
  SIGNAL Logical_Operator_out2371_out1            : std_logic;
  SIGNAL Logical_Operator_out2372_out1            : std_logic;
  SIGNAL Logical_Operator_out2373_out1            : std_logic;
  SIGNAL Logical_Operator_out2374_out1            : std_logic;
  SIGNAL Logical_Operator_out2375_out1            : std_logic;
  SIGNAL Logical_Operator_out2376_out1            : std_logic;
  SIGNAL Logical_Operator_out2377_out1            : std_logic;
  SIGNAL Logical_Operator_out2378_out1            : std_logic;
  SIGNAL Logical_Operator_out2379_out1            : std_logic;
  SIGNAL Logical_Operator_out2380_out1            : std_logic;
  SIGNAL Logical_Operator_out2381_out1            : std_logic;
  SIGNAL Logical_Operator_out2382_out1            : std_logic;
  SIGNAL Logical_Operator_out2383_out1            : std_logic;
  SIGNAL Logical_Operator_out2384_out1            : std_logic;
  SIGNAL Logical_Operator_out2385_out1            : std_logic;
  SIGNAL Logical_Operator_out2386_out1            : std_logic;
  SIGNAL Logical_Operator_out2387_out1            : std_logic;
  SIGNAL Logical_Operator_out2388_out1            : std_logic;
  SIGNAL Logical_Operator_out2389_out1            : std_logic;
  SIGNAL Logical_Operator_out2390_out1            : std_logic;
  SIGNAL Logical_Operator_out2391_out1            : std_logic;
  SIGNAL Logical_Operator_out2392_out1            : std_logic;
  SIGNAL Logical_Operator_out2393_out1            : std_logic;
  SIGNAL Logical_Operator_out2394_out1            : std_logic;
  SIGNAL Logical_Operator_out2395_out1            : std_logic;
  SIGNAL Logical_Operator_out2396_out1            : std_logic;
  SIGNAL Logical_Operator_out2397_out1            : std_logic;
  SIGNAL Logical_Operator_out2398_out1            : std_logic;
  SIGNAL Logical_Operator_out2399_out1            : std_logic;
  SIGNAL Logical_Operator_out2400_out1            : std_logic;
  SIGNAL Logical_Operator_out2401_out1            : std_logic;
  SIGNAL Logical_Operator_out2402_out1            : std_logic;
  SIGNAL Logical_Operator_out2403_out1            : std_logic;
  SIGNAL Logical_Operator_out2404_out1            : std_logic;
  SIGNAL Logical_Operator_out2405_out1            : std_logic;
  SIGNAL Logical_Operator_out2406_out1            : std_logic;
  SIGNAL Logical_Operator_out2407_out1            : std_logic;
  SIGNAL Logical_Operator_out2408_out1            : std_logic;
  SIGNAL Logical_Operator_out2409_out1            : std_logic;
  SIGNAL Logical_Operator_out2410_out1            : std_logic;
  SIGNAL Logical_Operator_out2411_out1            : std_logic;
  SIGNAL Logical_Operator_out2412_out1            : std_logic;
  SIGNAL Logical_Operator_out2413_out1            : std_logic;
  SIGNAL Logical_Operator_out2414_out1            : std_logic;
  SIGNAL Logical_Operator_out2415_out1            : std_logic;
  SIGNAL Logical_Operator_out2416_out1            : std_logic;
  SIGNAL Logical_Operator_out2417_out1            : std_logic;
  SIGNAL Logical_Operator_out2418_out1            : std_logic;
  SIGNAL Logical_Operator_out2419_out1            : std_logic;
  SIGNAL Logical_Operator_out2420_out1            : std_logic;
  SIGNAL Logical_Operator_out2421_out1            : std_logic;
  SIGNAL Logical_Operator_out2422_out1            : std_logic;
  SIGNAL Logical_Operator_out2423_out1            : std_logic;
  SIGNAL Logical_Operator_out2424_out1            : std_logic;
  SIGNAL Logical_Operator_out2425_out1            : std_logic;
  SIGNAL Logical_Operator_out2426_out1            : std_logic;
  SIGNAL Logical_Operator_out2427_out1            : std_logic;
  SIGNAL Logical_Operator_out2428_out1            : std_logic;
  SIGNAL Logical_Operator_out2429_out1            : std_logic;
  SIGNAL Logical_Operator_out2430_out1            : std_logic;
  SIGNAL Logical_Operator_out2431_out1            : std_logic;
  SIGNAL Logical_Operator_out2432_out1            : std_logic;
  SIGNAL Logical_Operator_out2433_out1            : std_logic;
  SIGNAL Logical_Operator_out2434_out1            : std_logic;
  SIGNAL Logical_Operator_out2435_out1            : std_logic;
  SIGNAL Logical_Operator_out2436_out1            : std_logic;
  SIGNAL Logical_Operator_out2437_out1            : std_logic;
  SIGNAL Logical_Operator_out2438_out1            : std_logic;
  SIGNAL Logical_Operator_out2439_out1            : std_logic;
  SIGNAL Logical_Operator_out2440_out1            : std_logic;
  SIGNAL Logical_Operator_out2441_out1            : std_logic;
  SIGNAL Logical_Operator_out2442_out1            : std_logic;
  SIGNAL Logical_Operator_out2443_out1            : std_logic;
  SIGNAL Logical_Operator_out2444_out1            : std_logic;
  SIGNAL Logical_Operator_out2445_out1            : std_logic;
  SIGNAL Logical_Operator_out2446_out1            : std_logic;
  SIGNAL Logical_Operator_out2447_out1            : std_logic;
  SIGNAL Logical_Operator_out2448_out1            : std_logic;
  SIGNAL Logical_Operator_out2449_out1            : std_logic;
  SIGNAL Logical_Operator_out2450_out1            : std_logic;
  SIGNAL Logical_Operator_out2451_out1            : std_logic;
  SIGNAL Logical_Operator_out2452_out1            : std_logic;
  SIGNAL Logical_Operator_out2453_out1            : std_logic;
  SIGNAL Logical_Operator_out2454_out1            : std_logic;
  SIGNAL Logical_Operator_out2455_out1            : std_logic;
  SIGNAL Logical_Operator_out2456_out1            : std_logic;
  SIGNAL Logical_Operator_out2457_out1            : std_logic;
  SIGNAL Logical_Operator_out2458_out1            : std_logic;
  SIGNAL Logical_Operator_out2459_out1            : std_logic;
  SIGNAL Logical_Operator_out2460_out1            : std_logic;
  SIGNAL Logical_Operator_out2461_out1            : std_logic;
  SIGNAL Logical_Operator_out2462_out1            : std_logic;
  SIGNAL Logical_Operator_out2463_out1            : std_logic;
  SIGNAL Logical_Operator_out2464_out1            : std_logic;
  SIGNAL Logical_Operator_out2465_out1            : std_logic;
  SIGNAL Logical_Operator_out2466_out1            : std_logic;
  SIGNAL Logical_Operator_out2467_out1            : std_logic;
  SIGNAL Logical_Operator_out2468_out1            : std_logic;
  SIGNAL Logical_Operator_out2469_out1            : std_logic;
  SIGNAL Logical_Operator_out2470_out1            : std_logic;
  SIGNAL Logical_Operator_out2471_out1            : std_logic;
  SIGNAL Logical_Operator_out2472_out1            : std_logic;
  SIGNAL Logical_Operator_out2473_out1            : std_logic;
  SIGNAL Logical_Operator_out2474_out1            : std_logic;
  SIGNAL Logical_Operator_out2475_out1            : std_logic;
  SIGNAL Logical_Operator_out2476_out1            : std_logic;
  SIGNAL Logical_Operator_out2477_out1            : std_logic;
  SIGNAL Logical_Operator_out2478_out1            : std_logic;
  SIGNAL Logical_Operator_out2479_out1            : std_logic;
  SIGNAL Logical_Operator_out2480_out1            : std_logic;
  SIGNAL Logical_Operator_out2481_out1            : std_logic;
  SIGNAL Logical_Operator_out2482_out1            : std_logic;
  SIGNAL Logical_Operator_out2483_out1            : std_logic;
  SIGNAL Logical_Operator_out2484_out1            : std_logic;
  SIGNAL Logical_Operator_out2485_out1            : std_logic;
  SIGNAL Logical_Operator_out2486_out1            : std_logic;
  SIGNAL Logical_Operator_out2487_out1            : std_logic;
  SIGNAL Logical_Operator_out2488_out1            : std_logic;
  SIGNAL Logical_Operator_out2489_out1            : std_logic;
  SIGNAL Logical_Operator_out2490_out1            : std_logic;
  SIGNAL Logical_Operator_out2491_out1            : std_logic;
  SIGNAL Logical_Operator_out2492_out1            : std_logic;
  SIGNAL Logical_Operator_out2493_out1            : std_logic;
  SIGNAL Logical_Operator_out2494_out1            : std_logic;
  SIGNAL Logical_Operator_out2495_out1            : std_logic;
  SIGNAL Logical_Operator_out2496_out1            : std_logic;
  SIGNAL Logical_Operator_out2497_out1            : std_logic;
  SIGNAL Logical_Operator_out2498_out1            : std_logic;
  SIGNAL Logical_Operator_out2499_out1            : std_logic;
  SIGNAL Logical_Operator_out2500_out1            : std_logic;
  SIGNAL Logical_Operator_out2501_out1            : std_logic;
  SIGNAL Logical_Operator_out2502_out1            : std_logic;
  SIGNAL Logical_Operator_out2503_out1            : std_logic;
  SIGNAL Logical_Operator_out2504_out1            : std_logic;
  SIGNAL Logical_Operator_out2505_out1            : std_logic;
  SIGNAL Logical_Operator_out2506_out1            : std_logic;
  SIGNAL Logical_Operator_out2507_out1            : std_logic;
  SIGNAL Logical_Operator_out2508_out1            : std_logic;
  SIGNAL Logical_Operator_out2509_out1            : std_logic;
  SIGNAL Logical_Operator_out2510_out1            : std_logic;
  SIGNAL Logical_Operator_out2511_out1            : std_logic;
  SIGNAL Logical_Operator_out2512_out1            : std_logic;
  SIGNAL Logical_Operator_out2513_out1            : std_logic;
  SIGNAL Logical_Operator_out2514_out1            : std_logic;
  SIGNAL Logical_Operator_out2515_out1            : std_logic;
  SIGNAL Logical_Operator_out2516_out1            : std_logic;
  SIGNAL Logical_Operator_out2517_out1            : std_logic;
  SIGNAL Logical_Operator_out2518_out1            : std_logic;
  SIGNAL Logical_Operator_out2519_out1            : std_logic;
  SIGNAL Logical_Operator_out2520_out1            : std_logic;
  SIGNAL Logical_Operator_out2521_out1            : std_logic;
  SIGNAL Logical_Operator_out2522_out1            : std_logic;
  SIGNAL Logical_Operator_out2523_out1            : std_logic;
  SIGNAL Logical_Operator_out2524_out1            : std_logic;
  SIGNAL Logical_Operator_out2525_out1            : std_logic;
  SIGNAL Logical_Operator_out2526_out1            : std_logic;
  SIGNAL Logical_Operator_out2527_out1            : std_logic;
  SIGNAL Logical_Operator_out2528_out1            : std_logic;
  SIGNAL Logical_Operator_out2529_out1            : std_logic;
  SIGNAL Logical_Operator_out2530_out1            : std_logic;
  SIGNAL Logical_Operator_out2531_out1            : std_logic;
  SIGNAL Logical_Operator_out2532_out1            : std_logic;
  SIGNAL Logical_Operator_out2533_out1            : std_logic;
  SIGNAL Logical_Operator_out2534_out1            : std_logic;
  SIGNAL Logical_Operator_out2535_out1            : std_logic;
  SIGNAL Logical_Operator_out2536_out1            : std_logic;
  SIGNAL Logical_Operator_out2537_out1            : std_logic;
  SIGNAL Logical_Operator_out2538_out1            : std_logic;
  SIGNAL Logical_Operator_out2539_out1            : std_logic;
  SIGNAL Logical_Operator_out2540_out1            : std_logic;
  SIGNAL Logical_Operator_out2541_out1            : std_logic;
  SIGNAL Logical_Operator_out2542_out1            : std_logic;
  SIGNAL Logical_Operator_out2543_out1            : std_logic;
  SIGNAL Logical_Operator_out2544_out1            : std_logic;
  SIGNAL Logical_Operator_out2545_out1            : std_logic;
  SIGNAL Logical_Operator_out2546_out1            : std_logic;
  SIGNAL Logical_Operator_out2547_out1            : std_logic;
  SIGNAL Logical_Operator_out2548_out1            : std_logic;
  SIGNAL Logical_Operator_out2549_out1            : std_logic;
  SIGNAL Logical_Operator_out2550_out1            : std_logic;
  SIGNAL Logical_Operator_out2551_out1            : std_logic;
  SIGNAL Logical_Operator_out2552_out1            : std_logic;
  SIGNAL Logical_Operator_out2553_out1            : std_logic;
  SIGNAL Logical_Operator_out2554_out1            : std_logic;
  SIGNAL Logical_Operator_out2555_out1            : std_logic;
  SIGNAL Logical_Operator_out2556_out1            : std_logic;
  SIGNAL Logical_Operator_out2557_out1            : std_logic;
  SIGNAL Logical_Operator_out2558_out1            : std_logic;
  SIGNAL Logical_Operator_out2559_out1            : std_logic;
  SIGNAL Logical_Operator_out2560_out1            : std_logic;
  SIGNAL Logical_Operator_out2561_out1            : std_logic;
  SIGNAL Logical_Operator_out2562_out1            : std_logic;
  SIGNAL Logical_Operator_out2563_out1            : std_logic;
  SIGNAL Logical_Operator_out2564_out1            : std_logic;
  SIGNAL Logical_Operator_out2565_out1            : std_logic;
  SIGNAL Logical_Operator_out2566_out1            : std_logic;
  SIGNAL Logical_Operator_out2567_out1            : std_logic;
  SIGNAL Logical_Operator_out2568_out1            : std_logic;
  SIGNAL Logical_Operator_out2569_out1            : std_logic;
  SIGNAL Logical_Operator_out2570_out1            : std_logic;
  SIGNAL Logical_Operator_out2571_out1            : std_logic;
  SIGNAL Logical_Operator_out2572_out1            : std_logic;
  SIGNAL Logical_Operator_out2573_out1            : std_logic;
  SIGNAL Logical_Operator_out2574_out1            : std_logic;
  SIGNAL Logical_Operator_out2575_out1            : std_logic;
  SIGNAL Logical_Operator_out2576_out1            : std_logic;
  SIGNAL Logical_Operator_out2577_out1            : std_logic;
  SIGNAL Logical_Operator_out2578_out1            : std_logic;
  SIGNAL Logical_Operator_out2579_out1            : std_logic;
  SIGNAL Logical_Operator_out2580_out1            : std_logic;
  SIGNAL Logical_Operator_out2581_out1            : std_logic;
  SIGNAL Logical_Operator_out2582_out1            : std_logic;
  SIGNAL Logical_Operator_out2583_out1            : std_logic;
  SIGNAL Logical_Operator_out2584_out1            : std_logic;
  SIGNAL Logical_Operator_out2585_out1            : std_logic;
  SIGNAL Logical_Operator_out2586_out1            : std_logic;
  SIGNAL Logical_Operator_out2587_out1            : std_logic;
  SIGNAL Logical_Operator_out2588_out1            : std_logic;
  SIGNAL Logical_Operator_out2589_out1            : std_logic;
  SIGNAL Logical_Operator_out2590_out1            : std_logic;
  SIGNAL Logical_Operator_out2591_out1            : std_logic;
  SIGNAL Logical_Operator_out2592_out1            : std_logic;
  SIGNAL Logical_Operator_out2593_out1            : std_logic;
  SIGNAL Logical_Operator_out2594_out1            : std_logic;
  SIGNAL Logical_Operator_out2595_out1            : std_logic;
  SIGNAL Logical_Operator_out2596_out1            : std_logic;
  SIGNAL Logical_Operator_out2597_out1            : std_logic;
  SIGNAL Logical_Operator_out2598_out1            : std_logic;
  SIGNAL Logical_Operator_out2599_out1            : std_logic;
  SIGNAL Logical_Operator_out2600_out1            : std_logic;
  SIGNAL Logical_Operator_out2601_out1            : std_logic;
  SIGNAL Logical_Operator_out2602_out1            : std_logic;
  SIGNAL Logical_Operator_out2603_out1            : std_logic;
  SIGNAL Logical_Operator_out2604_out1            : std_logic;
  SIGNAL Logical_Operator_out2605_out1            : std_logic;
  SIGNAL Logical_Operator_out2606_out1            : std_logic;
  SIGNAL Logical_Operator_out2607_out1            : std_logic;
  SIGNAL Logical_Operator_out2608_out1            : std_logic;
  SIGNAL Logical_Operator_out2609_out1            : std_logic;
  SIGNAL Logical_Operator_out2610_out1            : std_logic;
  SIGNAL Logical_Operator_out2611_out1            : std_logic;
  SIGNAL Logical_Operator_out2612_out1            : std_logic;
  SIGNAL Logical_Operator_out2613_out1            : std_logic;
  SIGNAL Logical_Operator_out2614_out1            : std_logic;
  SIGNAL Logical_Operator_out2615_out1            : std_logic;
  SIGNAL Logical_Operator_out2616_out1            : std_logic;
  SIGNAL Logical_Operator_out2617_out1            : std_logic;
  SIGNAL Logical_Operator_out2618_out1            : std_logic;
  SIGNAL Logical_Operator_out2619_out1            : std_logic;
  SIGNAL Logical_Operator_out2620_out1            : std_logic;
  SIGNAL Logical_Operator_out2621_out1            : std_logic;
  SIGNAL Logical_Operator_out2622_out1            : std_logic;
  SIGNAL Logical_Operator_out2623_out1            : std_logic;
  SIGNAL Logical_Operator_out2624_out1            : std_logic;
  SIGNAL Logical_Operator_out2625_out1            : std_logic;
  SIGNAL Logical_Operator_out2626_out1            : std_logic;
  SIGNAL Logical_Operator_out2627_out1            : std_logic;
  SIGNAL Logical_Operator_out2628_out1            : std_logic;
  SIGNAL Logical_Operator_out2629_out1            : std_logic;
  SIGNAL Logical_Operator_out2630_out1            : std_logic;
  SIGNAL Logical_Operator_out2631_out1            : std_logic;
  SIGNAL Logical_Operator_out2632_out1            : std_logic;
  SIGNAL Logical_Operator_out2633_out1            : std_logic;
  SIGNAL Logical_Operator_out2634_out1            : std_logic;
  SIGNAL Logical_Operator_out2635_out1            : std_logic;
  SIGNAL Logical_Operator_out2636_out1            : std_logic;
  SIGNAL Logical_Operator_out2637_out1            : std_logic;
  SIGNAL Logical_Operator_out2638_out1            : std_logic;
  SIGNAL Logical_Operator_out2639_out1            : std_logic;
  SIGNAL Logical_Operator_out2640_out1            : std_logic;
  SIGNAL Logical_Operator_out2641_out1            : std_logic;
  SIGNAL Logical_Operator_out2642_out1            : std_logic;
  SIGNAL Logical_Operator_out2643_out1            : std_logic;
  SIGNAL Logical_Operator_out2644_out1            : std_logic;
  SIGNAL Logical_Operator_out2645_out1            : std_logic;
  SIGNAL Logical_Operator_out2646_out1            : std_logic;
  SIGNAL Logical_Operator_out2647_out1            : std_logic;
  SIGNAL Logical_Operator_out2648_out1            : std_logic;
  SIGNAL Logical_Operator_out2649_out1            : std_logic;
  SIGNAL Logical_Operator_out2650_out1            : std_logic;
  SIGNAL Logical_Operator_out2651_out1            : std_logic;
  SIGNAL Logical_Operator_out2652_out1            : std_logic;
  SIGNAL Logical_Operator_out2653_out1            : std_logic;
  SIGNAL Logical_Operator_out2654_out1            : std_logic;
  SIGNAL Logical_Operator_out2655_out1            : std_logic;
  SIGNAL Logical_Operator_out2656_out1            : std_logic;
  SIGNAL Logical_Operator_out2657_out1            : std_logic;
  SIGNAL Logical_Operator_out2658_out1            : std_logic;
  SIGNAL Logical_Operator_out2659_out1            : std_logic;
  SIGNAL Logical_Operator_out2660_out1            : std_logic;
  SIGNAL Logical_Operator_out2661_out1            : std_logic;
  SIGNAL Logical_Operator_out2662_out1            : std_logic;
  SIGNAL Logical_Operator_out2663_out1            : std_logic;
  SIGNAL Logical_Operator_out2664_out1            : std_logic;
  SIGNAL Logical_Operator_out2665_out1            : std_logic;
  SIGNAL Logical_Operator_out2666_out1            : std_logic;
  SIGNAL Logical_Operator_out2667_out1            : std_logic;
  SIGNAL Logical_Operator_out2668_out1            : std_logic;
  SIGNAL Logical_Operator_out2669_out1            : std_logic;
  SIGNAL Logical_Operator_out2670_out1            : std_logic;
  SIGNAL Logical_Operator_out2671_out1            : std_logic;
  SIGNAL Logical_Operator_out2672_out1            : std_logic;
  SIGNAL Logical_Operator_out2673_out1            : std_logic;
  SIGNAL Logical_Operator_out2674_out1            : std_logic;
  SIGNAL Logical_Operator_out2675_out1            : std_logic;
  SIGNAL Logical_Operator_out2676_out1            : std_logic;
  SIGNAL Logical_Operator_out2677_out1            : std_logic;
  SIGNAL Logical_Operator_out2678_out1            : std_logic;
  SIGNAL Logical_Operator_out2679_out1            : std_logic;
  SIGNAL Logical_Operator_out2680_out1            : std_logic;
  SIGNAL Logical_Operator_out2681_out1            : std_logic;
  SIGNAL Logical_Operator_out2682_out1            : std_logic;
  SIGNAL Logical_Operator_out2683_out1            : std_logic;
  SIGNAL Logical_Operator_out2684_out1            : std_logic;
  SIGNAL Logical_Operator_out2685_out1            : std_logic;
  SIGNAL Logical_Operator_out2686_out1            : std_logic;
  SIGNAL Logical_Operator_out2687_out1            : std_logic;
  SIGNAL Logical_Operator_out2688_out1            : std_logic;
  SIGNAL Logical_Operator_out2689_out1            : std_logic;
  SIGNAL Logical_Operator_out2690_out1            : std_logic;
  SIGNAL Logical_Operator_out2691_out1            : std_logic;
  SIGNAL Logical_Operator_out2692_out1            : std_logic;
  SIGNAL Logical_Operator_out2693_out1            : std_logic;
  SIGNAL Logical_Operator_out2694_out1            : std_logic;
  SIGNAL Logical_Operator_out2695_out1            : std_logic;
  SIGNAL Logical_Operator_out2696_out1            : std_logic;
  SIGNAL Logical_Operator_out2697_out1            : std_logic;
  SIGNAL Logical_Operator_out2698_out1            : std_logic;
  SIGNAL Logical_Operator_out2699_out1            : std_logic;
  SIGNAL Logical_Operator_out2700_out1            : std_logic;
  SIGNAL Logical_Operator_out2701_out1            : std_logic;
  SIGNAL Logical_Operator_out2702_out1            : std_logic;
  SIGNAL Logical_Operator_out2703_out1            : std_logic;
  SIGNAL Logical_Operator_out2704_out1            : std_logic;
  SIGNAL Logical_Operator_out2705_out1            : std_logic;
  SIGNAL Logical_Operator_out2706_out1            : std_logic;
  SIGNAL Logical_Operator_out2707_out1            : std_logic;
  SIGNAL Logical_Operator_out2708_out1            : std_logic;
  SIGNAL Logical_Operator_out2709_out1            : std_logic;
  SIGNAL Logical_Operator_out2710_out1            : std_logic;
  SIGNAL Logical_Operator_out2711_out1            : std_logic;
  SIGNAL Logical_Operator_out2712_out1            : std_logic;
  SIGNAL Logical_Operator_out2713_out1            : std_logic;
  SIGNAL Logical_Operator_out2714_out1            : std_logic;
  SIGNAL Logical_Operator_out2715_out1            : std_logic;
  SIGNAL Logical_Operator_out2716_out1            : std_logic;
  SIGNAL Logical_Operator_out2717_out1            : std_logic;
  SIGNAL Logical_Operator_out2718_out1            : std_logic;
  SIGNAL Logical_Operator_out2719_out1            : std_logic;
  SIGNAL Logical_Operator_out2720_out1            : std_logic;
  SIGNAL Logical_Operator_out2721_out1            : std_logic;
  SIGNAL Logical_Operator_out2722_out1            : std_logic;
  SIGNAL Logical_Operator_out2723_out1            : std_logic;
  SIGNAL Logical_Operator_out2724_out1            : std_logic;
  SIGNAL Logical_Operator_out2725_out1            : std_logic;
  SIGNAL Logical_Operator_out2726_out1            : std_logic;
  SIGNAL Logical_Operator_out2727_out1            : std_logic;
  SIGNAL Logical_Operator_out2728_out1            : std_logic;
  SIGNAL Logical_Operator_out2729_out1            : std_logic;
  SIGNAL Logical_Operator_out2730_out1            : std_logic;
  SIGNAL Logical_Operator_out2731_out1            : std_logic;
  SIGNAL Logical_Operator_out2732_out1            : std_logic;
  SIGNAL Logical_Operator_out2733_out1            : std_logic;
  SIGNAL Logical_Operator_out2734_out1            : std_logic;
  SIGNAL Logical_Operator_out2735_out1            : std_logic;
  SIGNAL Logical_Operator_out2736_out1            : std_logic;
  SIGNAL Logical_Operator_out2737_out1            : std_logic;
  SIGNAL Logical_Operator_out2738_out1            : std_logic;
  SIGNAL Logical_Operator_out2739_out1            : std_logic;
  SIGNAL Logical_Operator_out2740_out1            : std_logic;
  SIGNAL Logical_Operator_out2741_out1            : std_logic;
  SIGNAL Logical_Operator_out2742_out1            : std_logic;
  SIGNAL Logical_Operator_out2743_out1            : std_logic;
  SIGNAL Logical_Operator_out2744_out1            : std_logic;
  SIGNAL Logical_Operator_out2745_out1            : std_logic;
  SIGNAL Logical_Operator_out2746_out1            : std_logic;
  SIGNAL Logical_Operator_out2747_out1            : std_logic;
  SIGNAL Logical_Operator_out2748_out1            : std_logic;
  SIGNAL Logical_Operator_out2749_out1            : std_logic;
  SIGNAL Logical_Operator_out2750_out1            : std_logic;
  SIGNAL Logical_Operator_out2751_out1            : std_logic;
  SIGNAL Logical_Operator_out2752_out1            : std_logic;
  SIGNAL Logical_Operator_out2753_out1            : std_logic;
  SIGNAL Logical_Operator_out2754_out1            : std_logic;
  SIGNAL Logical_Operator_out2755_out1            : std_logic;
  SIGNAL Logical_Operator_out2756_out1            : std_logic;
  SIGNAL Logical_Operator_out2757_out1            : std_logic;
  SIGNAL Logical_Operator_out2758_out1            : std_logic;
  SIGNAL Logical_Operator_out2759_out1            : std_logic;
  SIGNAL Logical_Operator_out2760_out1            : std_logic;
  SIGNAL Logical_Operator_out2761_out1            : std_logic;
  SIGNAL Logical_Operator_out2762_out1            : std_logic;
  SIGNAL Logical_Operator_out2763_out1            : std_logic;
  SIGNAL Logical_Operator_out2764_out1            : std_logic;
  SIGNAL Logical_Operator_out2765_out1            : std_logic;
  SIGNAL Logical_Operator_out2766_out1            : std_logic;
  SIGNAL Logical_Operator_out2767_out1            : std_logic;
  SIGNAL Logical_Operator_out2768_out1            : std_logic;
  SIGNAL Logical_Operator_out2769_out1            : std_logic;
  SIGNAL Logical_Operator_out2770_out1            : std_logic;
  SIGNAL Logical_Operator_out2771_out1            : std_logic;
  SIGNAL Logical_Operator_out2772_out1            : std_logic;
  SIGNAL Logical_Operator_out2773_out1            : std_logic;
  SIGNAL Logical_Operator_out2774_out1            : std_logic;
  SIGNAL Logical_Operator_out2775_out1            : std_logic;
  SIGNAL Logical_Operator_out2776_out1            : std_logic;
  SIGNAL Logical_Operator_out2777_out1            : std_logic;
  SIGNAL Logical_Operator_out2778_out1            : std_logic;
  SIGNAL Logical_Operator_out2779_out1            : std_logic;
  SIGNAL Logical_Operator_out2780_out1            : std_logic;
  SIGNAL Logical_Operator_out2781_out1            : std_logic;
  SIGNAL Logical_Operator_out2782_out1            : std_logic;
  SIGNAL Logical_Operator_out2783_out1            : std_logic;
  SIGNAL Logical_Operator_out2784_out1            : std_logic;
  SIGNAL Logical_Operator_out2785_out1            : std_logic;
  SIGNAL Logical_Operator_out2786_out1            : std_logic;
  SIGNAL Logical_Operator_out2787_out1            : std_logic;
  SIGNAL Logical_Operator_out2788_out1            : std_logic;
  SIGNAL Logical_Operator_out2789_out1            : std_logic;
  SIGNAL Logical_Operator_out2790_out1            : std_logic;
  SIGNAL Logical_Operator_out2791_out1            : std_logic;
  SIGNAL Logical_Operator_out2792_out1            : std_logic;
  SIGNAL Logical_Operator_out2793_out1            : std_logic;
  SIGNAL Logical_Operator_out2794_out1            : std_logic;
  SIGNAL Logical_Operator_out2795_out1            : std_logic;
  SIGNAL Logical_Operator_out2796_out1            : std_logic;
  SIGNAL Logical_Operator_out2797_out1            : std_logic;
  SIGNAL Logical_Operator_out2798_out1            : std_logic;
  SIGNAL Logical_Operator_out2799_out1            : std_logic;
  SIGNAL Logical_Operator_out2800_out1            : std_logic;
  SIGNAL Logical_Operator_out2801_out1            : std_logic;
  SIGNAL Logical_Operator_out2802_out1            : std_logic;
  SIGNAL Logical_Operator_out2803_out1            : std_logic;
  SIGNAL Logical_Operator_out2804_out1            : std_logic;
  SIGNAL Logical_Operator_out2805_out1            : std_logic;
  SIGNAL Logical_Operator_out2806_out1            : std_logic;
  SIGNAL Logical_Operator_out2807_out1            : std_logic;
  SIGNAL Logical_Operator_out2808_out1            : std_logic;
  SIGNAL Logical_Operator_out2809_out1            : std_logic;
  SIGNAL Logical_Operator_out2810_out1            : std_logic;
  SIGNAL Logical_Operator_out2811_out1            : std_logic;
  SIGNAL Logical_Operator_out2812_out1            : std_logic;
  SIGNAL Logical_Operator_out2813_out1            : std_logic;
  SIGNAL Logical_Operator_out2814_out1            : std_logic;
  SIGNAL Logical_Operator_out2815_out1            : std_logic;
  SIGNAL Logical_Operator_out2816_out1            : std_logic;
  SIGNAL Logical_Operator_out2817_out1            : std_logic;
  SIGNAL Logical_Operator_out2818_out1            : std_logic;
  SIGNAL Logical_Operator_out2819_out1            : std_logic;
  SIGNAL Logical_Operator_out2820_out1            : std_logic;
  SIGNAL Logical_Operator_out2821_out1            : std_logic;
  SIGNAL Logical_Operator_out2822_out1            : std_logic;
  SIGNAL Logical_Operator_out2823_out1            : std_logic;
  SIGNAL Logical_Operator_out2824_out1            : std_logic;
  SIGNAL Logical_Operator_out2825_out1            : std_logic;
  SIGNAL Logical_Operator_out2826_out1            : std_logic;
  SIGNAL Logical_Operator_out2827_out1            : std_logic;
  SIGNAL Logical_Operator_out2828_out1            : std_logic;
  SIGNAL Logical_Operator_out2829_out1            : std_logic;
  SIGNAL Logical_Operator_out2830_out1            : std_logic;
  SIGNAL Logical_Operator_out2831_out1            : std_logic;
  SIGNAL Logical_Operator_out2832_out1            : std_logic;
  SIGNAL Logical_Operator_out2833_out1            : std_logic;
  SIGNAL Logical_Operator_out2834_out1            : std_logic;
  SIGNAL Logical_Operator_out2835_out1            : std_logic;
  SIGNAL Logical_Operator_out2836_out1            : std_logic;
  SIGNAL Logical_Operator_out2837_out1            : std_logic;
  SIGNAL Logical_Operator_out2838_out1            : std_logic;
  SIGNAL Logical_Operator_out2839_out1            : std_logic;
  SIGNAL Logical_Operator_out2840_out1            : std_logic;
  SIGNAL Logical_Operator_out2841_out1            : std_logic;
  SIGNAL Logical_Operator_out2842_out1            : std_logic;
  SIGNAL Logical_Operator_out2843_out1            : std_logic;
  SIGNAL Logical_Operator_out2844_out1            : std_logic;
  SIGNAL Logical_Operator_out2845_out1            : std_logic;
  SIGNAL Logical_Operator_out2846_out1            : std_logic;
  SIGNAL Logical_Operator_out2847_out1            : std_logic;
  SIGNAL Logical_Operator_out2848_out1            : std_logic;
  SIGNAL Logical_Operator_out2849_out1            : std_logic;
  SIGNAL Logical_Operator_out2850_out1            : std_logic;
  SIGNAL Logical_Operator_out2851_out1            : std_logic;
  SIGNAL Logical_Operator_out2852_out1            : std_logic;
  SIGNAL Logical_Operator_out2853_out1            : std_logic;
  SIGNAL Logical_Operator_out2854_out1            : std_logic;
  SIGNAL Logical_Operator_out2855_out1            : std_logic;
  SIGNAL Logical_Operator_out2856_out1            : std_logic;
  SIGNAL Logical_Operator_out2857_out1            : std_logic;
  SIGNAL Logical_Operator_out2858_out1            : std_logic;
  SIGNAL Logical_Operator_out2859_out1            : std_logic;
  SIGNAL Logical_Operator_out2860_out1            : std_logic;
  SIGNAL Logical_Operator_out2861_out1            : std_logic;
  SIGNAL Logical_Operator_out2862_out1            : std_logic;
  SIGNAL Logical_Operator_out2863_out1            : std_logic;
  SIGNAL Logical_Operator_out2864_out1            : std_logic;
  SIGNAL Logical_Operator_out2865_out1            : std_logic;
  SIGNAL Logical_Operator_out2866_out1            : std_logic;
  SIGNAL Logical_Operator_out2867_out1            : std_logic;
  SIGNAL Logical_Operator_out2868_out1            : std_logic;
  SIGNAL Logical_Operator_out2869_out1            : std_logic;
  SIGNAL Logical_Operator_out2870_out1            : std_logic;
  SIGNAL Logical_Operator_out2871_out1            : std_logic;
  SIGNAL Logical_Operator_out2872_out1            : std_logic;
  SIGNAL Logical_Operator_out2873_out1            : std_logic;
  SIGNAL Logical_Operator_out2874_out1            : std_logic;
  SIGNAL Logical_Operator_out2875_out1            : std_logic;
  SIGNAL Logical_Operator_out2876_out1            : std_logic;
  SIGNAL Logical_Operator_out2877_out1            : std_logic;
  SIGNAL Logical_Operator_out2878_out1            : std_logic;
  SIGNAL Logical_Operator_out2879_out1            : std_logic;
  SIGNAL Logical_Operator_out2880_out1            : std_logic;
  SIGNAL Logical_Operator_out2881_out1            : std_logic;
  SIGNAL Logical_Operator_out2882_out1            : std_logic;
  SIGNAL Logical_Operator_out2883_out1            : std_logic;
  SIGNAL Logical_Operator_out2884_out1            : std_logic;
  SIGNAL Logical_Operator_out2885_out1            : std_logic;
  SIGNAL Logical_Operator_out2886_out1            : std_logic;
  SIGNAL Logical_Operator_out2887_out1            : std_logic;
  SIGNAL Logical_Operator_out2888_out1            : std_logic;
  SIGNAL Logical_Operator_out2889_out1            : std_logic;
  SIGNAL Logical_Operator_out2890_out1            : std_logic;
  SIGNAL Logical_Operator_out2891_out1            : std_logic;
  SIGNAL Logical_Operator_out2892_out1            : std_logic;
  SIGNAL Logical_Operator_out2893_out1            : std_logic;
  SIGNAL Logical_Operator_out2894_out1            : std_logic;
  SIGNAL Logical_Operator_out2895_out1            : std_logic;
  SIGNAL Logical_Operator_out2896_out1            : std_logic;
  SIGNAL Logical_Operator_out2897_out1            : std_logic;
  SIGNAL Logical_Operator_out2898_out1            : std_logic;
  SIGNAL Logical_Operator_out2899_out1            : std_logic;
  SIGNAL Logical_Operator_out2900_out1            : std_logic;
  SIGNAL Logical_Operator_out2901_out1            : std_logic;
  SIGNAL Logical_Operator_out2902_out1            : std_logic;
  SIGNAL Logical_Operator_out2903_out1            : std_logic;
  SIGNAL Logical_Operator_out2904_out1            : std_logic;
  SIGNAL Logical_Operator_out2905_out1            : std_logic;
  SIGNAL Logical_Operator_out2906_out1            : std_logic;
  SIGNAL Logical_Operator_out2907_out1            : std_logic;
  SIGNAL Logical_Operator_out2908_out1            : std_logic;
  SIGNAL Logical_Operator_out2909_out1            : std_logic;
  SIGNAL Logical_Operator_out2910_out1            : std_logic;
  SIGNAL Logical_Operator_out2911_out1            : std_logic;
  SIGNAL Logical_Operator_out2912_out1            : std_logic;
  SIGNAL Logical_Operator_out2913_out1            : std_logic;
  SIGNAL Logical_Operator_out2914_out1            : std_logic;
  SIGNAL Logical_Operator_out2915_out1            : std_logic;
  SIGNAL Logical_Operator_out2916_out1            : std_logic;
  SIGNAL Logical_Operator_out2917_out1            : std_logic;
  SIGNAL Logical_Operator_out2918_out1            : std_logic;
  SIGNAL Logical_Operator_out2919_out1            : std_logic;
  SIGNAL Logical_Operator_out2920_out1            : std_logic;
  SIGNAL Logical_Operator_out2921_out1            : std_logic;
  SIGNAL Logical_Operator_out2922_out1            : std_logic;
  SIGNAL Logical_Operator_out2923_out1            : std_logic;
  SIGNAL Logical_Operator_out2924_out1            : std_logic;
  SIGNAL Logical_Operator_out2925_out1            : std_logic;
  SIGNAL Logical_Operator_out2926_out1            : std_logic;
  SIGNAL Logical_Operator_out2927_out1            : std_logic;
  SIGNAL Logical_Operator_out2928_out1            : std_logic;
  SIGNAL Logical_Operator_out2929_out1            : std_logic;
  SIGNAL Logical_Operator_out2930_out1            : std_logic;
  SIGNAL Logical_Operator_out2931_out1            : std_logic;
  SIGNAL Logical_Operator_out2932_out1            : std_logic;
  SIGNAL Logical_Operator_out2933_out1            : std_logic;
  SIGNAL Logical_Operator_out2934_out1            : std_logic;
  SIGNAL Logical_Operator_out2935_out1            : std_logic;
  SIGNAL Logical_Operator_out2936_out1            : std_logic;
  SIGNAL Logical_Operator_out2937_out1            : std_logic;
  SIGNAL Logical_Operator_out2938_out1            : std_logic;
  SIGNAL Logical_Operator_out2939_out1            : std_logic;
  SIGNAL Logical_Operator_out2940_out1            : std_logic;
  SIGNAL Logical_Operator_out2941_out1            : std_logic;
  SIGNAL Logical_Operator_out2942_out1            : std_logic;
  SIGNAL Logical_Operator_out2943_out1            : std_logic;
  SIGNAL Logical_Operator_out2944_out1            : std_logic;
  SIGNAL Logical_Operator_out2945_out1            : std_logic;
  SIGNAL Logical_Operator_out2946_out1            : std_logic;
  SIGNAL Logical_Operator_out2947_out1            : std_logic;
  SIGNAL Logical_Operator_out2948_out1            : std_logic;
  SIGNAL Logical_Operator_out2949_out1            : std_logic;
  SIGNAL Logical_Operator_out2950_out1            : std_logic;
  SIGNAL Logical_Operator_out2951_out1            : std_logic;
  SIGNAL Logical_Operator_out2952_out1            : std_logic;
  SIGNAL Logical_Operator_out2953_out1            : std_logic;
  SIGNAL Logical_Operator_out2954_out1            : std_logic;
  SIGNAL Logical_Operator_out2955_out1            : std_logic;
  SIGNAL Logical_Operator_out2956_out1            : std_logic;
  SIGNAL Logical_Operator_out2957_out1            : std_logic;
  SIGNAL Logical_Operator_out2958_out1            : std_logic;
  SIGNAL Logical_Operator_out2959_out1            : std_logic;
  SIGNAL Logical_Operator_out2960_out1            : std_logic;
  SIGNAL Logical_Operator_out2961_out1            : std_logic;
  SIGNAL Logical_Operator_out2962_out1            : std_logic;
  SIGNAL Logical_Operator_out2963_out1            : std_logic;
  SIGNAL Logical_Operator_out2964_out1            : std_logic;
  SIGNAL Logical_Operator_out2965_out1            : std_logic;
  SIGNAL Logical_Operator_out2966_out1            : std_logic;
  SIGNAL Logical_Operator_out2967_out1            : std_logic;
  SIGNAL Logical_Operator_out2968_out1            : std_logic;
  SIGNAL Logical_Operator_out2969_out1            : std_logic;
  SIGNAL Logical_Operator_out2970_out1            : std_logic;
  SIGNAL Logical_Operator_out2971_out1            : std_logic;
  SIGNAL Logical_Operator_out2972_out1            : std_logic;
  SIGNAL Logical_Operator_out2973_out1            : std_logic;
  SIGNAL Logical_Operator_out2974_out1            : std_logic;
  SIGNAL Logical_Operator_out2975_out1            : std_logic;
  SIGNAL Logical_Operator_out2976_out1            : std_logic;
  SIGNAL Logical_Operator_out2977_out1            : std_logic;
  SIGNAL Logical_Operator_out2978_out1            : std_logic;
  SIGNAL Logical_Operator_out2979_out1            : std_logic;
  SIGNAL Logical_Operator_out2980_out1            : std_logic;
  SIGNAL Logical_Operator_out2981_out1            : std_logic;
  SIGNAL Logical_Operator_out2982_out1            : std_logic;
  SIGNAL Logical_Operator_out2983_out1            : std_logic;
  SIGNAL Logical_Operator_out2984_out1            : std_logic;
  SIGNAL Logical_Operator_out2985_out1            : std_logic;
  SIGNAL Logical_Operator_out2986_out1            : std_logic;
  SIGNAL Logical_Operator_out2987_out1            : std_logic;
  SIGNAL Logical_Operator_out2988_out1            : std_logic;
  SIGNAL Logical_Operator_out2989_out1            : std_logic;
  SIGNAL Logical_Operator_out2990_out1            : std_logic;
  SIGNAL Logical_Operator_out2991_out1            : std_logic;
  SIGNAL Logical_Operator_out2992_out1            : std_logic;
  SIGNAL Logical_Operator_out2993_out1            : std_logic;
  SIGNAL Logical_Operator_out2994_out1            : std_logic;
  SIGNAL Logical_Operator_out2995_out1            : std_logic;
  SIGNAL Logical_Operator_out2996_out1            : std_logic;
  SIGNAL Logical_Operator_out2997_out1            : std_logic;
  SIGNAL Logical_Operator_out2998_out1            : std_logic;
  SIGNAL Logical_Operator_out2999_out1            : std_logic;
  SIGNAL Logical_Operator_out3000_out1            : std_logic;
  SIGNAL Logical_Operator_out3001_out1            : std_logic;
  SIGNAL Logical_Operator_out3002_out1            : std_logic;
  SIGNAL Logical_Operator_out3003_out1            : std_logic;
  SIGNAL Logical_Operator_out3004_out1            : std_logic;
  SIGNAL Logical_Operator_out3005_out1            : std_logic;
  SIGNAL Logical_Operator_out3006_out1            : std_logic;
  SIGNAL Logical_Operator_out3007_out1            : std_logic;
  SIGNAL Logical_Operator_out3008_out1            : std_logic;
  SIGNAL Logical_Operator_out3009_out1            : std_logic;
  SIGNAL Logical_Operator_out3010_out1            : std_logic;
  SIGNAL Logical_Operator_out3011_out1            : std_logic;
  SIGNAL Logical_Operator_out3012_out1            : std_logic;
  SIGNAL Logical_Operator_out3013_out1            : std_logic;
  SIGNAL Logical_Operator_out3014_out1            : std_logic;
  SIGNAL Logical_Operator_out3015_out1            : std_logic;
  SIGNAL Logical_Operator_out3016_out1            : std_logic;
  SIGNAL Logical_Operator_out3017_out1            : std_logic;
  SIGNAL Logical_Operator_out3018_out1            : std_logic;
  SIGNAL Logical_Operator_out3019_out1            : std_logic;
  SIGNAL Logical_Operator_out3020_out1            : std_logic;
  SIGNAL Logical_Operator_out3021_out1            : std_logic;
  SIGNAL Logical_Operator_out3022_out1            : std_logic;
  SIGNAL Logical_Operator_out3023_out1            : std_logic;
  SIGNAL Logical_Operator_out3024_out1            : std_logic;
  SIGNAL Logical_Operator_out3025_out1            : std_logic;
  SIGNAL Logical_Operator_out3026_out1            : std_logic;
  SIGNAL Logical_Operator_out3027_out1            : std_logic;
  SIGNAL Logical_Operator_out3028_out1            : std_logic;
  SIGNAL Logical_Operator_out3029_out1            : std_logic;
  SIGNAL Logical_Operator_out3030_out1            : std_logic;
  SIGNAL Logical_Operator_out3031_out1            : std_logic;
  SIGNAL Logical_Operator_out3032_out1            : std_logic;
  SIGNAL Logical_Operator_out3033_out1            : std_logic;
  SIGNAL Logical_Operator_out3034_out1            : std_logic;
  SIGNAL Logical_Operator_out3035_out1            : std_logic;
  SIGNAL Logical_Operator_out3036_out1            : std_logic;
  SIGNAL Logical_Operator_out3037_out1            : std_logic;
  SIGNAL Logical_Operator_out3038_out1            : std_logic;
  SIGNAL Logical_Operator_out3039_out1            : std_logic;
  SIGNAL Logical_Operator_out3040_out1            : std_logic;
  SIGNAL Logical_Operator_out3041_out1            : std_logic;
  SIGNAL Logical_Operator_out3042_out1            : std_logic;
  SIGNAL Logical_Operator_out3043_out1            : std_logic;
  SIGNAL Logical_Operator_out3044_out1            : std_logic;
  SIGNAL Logical_Operator_out3045_out1            : std_logic;
  SIGNAL Logical_Operator_out3046_out1            : std_logic;
  SIGNAL Logical_Operator_out3047_out1            : std_logic;
  SIGNAL Logical_Operator_out3048_out1            : std_logic;
  SIGNAL Logical_Operator_out3049_out1            : std_logic;
  SIGNAL Logical_Operator_out3050_out1            : std_logic;
  SIGNAL Logical_Operator_out3051_out1            : std_logic;
  SIGNAL Logical_Operator_out3052_out1            : std_logic;
  SIGNAL Logical_Operator_out3053_out1            : std_logic;
  SIGNAL Logical_Operator_out3054_out1            : std_logic;
  SIGNAL Logical_Operator_out3055_out1            : std_logic;
  SIGNAL Logical_Operator_out3056_out1            : std_logic;
  SIGNAL Logical_Operator_out3057_out1            : std_logic;
  SIGNAL Logical_Operator_out3058_out1            : std_logic;
  SIGNAL Logical_Operator_out3059_out1            : std_logic;
  SIGNAL Logical_Operator_out3060_out1            : std_logic;
  SIGNAL Logical_Operator_out3061_out1            : std_logic;
  SIGNAL Logical_Operator_out3062_out1            : std_logic;
  SIGNAL Logical_Operator_out3063_out1            : std_logic;
  SIGNAL Logical_Operator_out3064_out1            : std_logic;
  SIGNAL Logical_Operator_out3065_out1            : std_logic;
  SIGNAL Logical_Operator_out3066_out1            : std_logic;
  SIGNAL Logical_Operator_out3067_out1            : std_logic;
  SIGNAL Logical_Operator_out3068_out1            : std_logic;
  SIGNAL Logical_Operator_out3069_out1            : std_logic;
  SIGNAL Logical_Operator_out3070_out1            : std_logic;
  SIGNAL Logical_Operator_out3071_out1            : std_logic;
  SIGNAL Logical_Operator_out3072_out1            : std_logic;
  SIGNAL Logical_Operator_out3073_out1            : std_logic;
  SIGNAL Logical_Operator_out3074_out1            : std_logic;
  SIGNAL Logical_Operator_out3075_out1            : std_logic;
  SIGNAL Logical_Operator_out3076_out1            : std_logic;
  SIGNAL Logical_Operator_out3077_out1            : std_logic;
  SIGNAL Logical_Operator_out3078_out1            : std_logic;
  SIGNAL Logical_Operator_out3079_out1            : std_logic;
  SIGNAL Logical_Operator_out3080_out1            : std_logic;
  SIGNAL Logical_Operator_out3081_out1            : std_logic;
  SIGNAL Logical_Operator_out3082_out1            : std_logic;
  SIGNAL Logical_Operator_out3083_out1            : std_logic;
  SIGNAL Logical_Operator_out3084_out1            : std_logic;
  SIGNAL Logical_Operator_out3085_out1            : std_logic;
  SIGNAL Logical_Operator_out3086_out1            : std_logic;
  SIGNAL Logical_Operator_out3087_out1            : std_logic;
  SIGNAL Logical_Operator_out3088_out1            : std_logic;
  SIGNAL Logical_Operator_out3089_out1            : std_logic;
  SIGNAL Logical_Operator_out3090_out1            : std_logic;
  SIGNAL Logical_Operator_out3091_out1            : std_logic;
  SIGNAL Logical_Operator_out3092_out1            : std_logic;
  SIGNAL Logical_Operator_out3093_out1            : std_logic;
  SIGNAL Logical_Operator_out3094_out1            : std_logic;
  SIGNAL Logical_Operator_out3095_out1            : std_logic;
  SIGNAL Logical_Operator_out3096_out1            : std_logic;
  SIGNAL Logical_Operator_out3097_out1            : std_logic;
  SIGNAL Logical_Operator_out3098_out1            : std_logic;
  SIGNAL Logical_Operator_out3099_out1            : std_logic;
  SIGNAL Logical_Operator_out3100_out1            : std_logic;
  SIGNAL Logical_Operator_out3101_out1            : std_logic;
  SIGNAL Logical_Operator_out3102_out1            : std_logic;
  SIGNAL Logical_Operator_out3103_out1            : std_logic;
  SIGNAL Logical_Operator_out3104_out1            : std_logic;
  SIGNAL Logical_Operator_out3105_out1            : std_logic;
  SIGNAL Logical_Operator_out3106_out1            : std_logic;
  SIGNAL Logical_Operator_out3107_out1            : std_logic;
  SIGNAL Logical_Operator_out3108_out1            : std_logic;
  SIGNAL Logical_Operator_out3109_out1            : std_logic;
  SIGNAL Logical_Operator_out3110_out1            : std_logic;
  SIGNAL Logical_Operator_out3111_out1            : std_logic;
  SIGNAL Logical_Operator_out3112_out1            : std_logic;
  SIGNAL Logical_Operator_out3113_out1            : std_logic;
  SIGNAL Logical_Operator_out3114_out1            : std_logic;
  SIGNAL Logical_Operator_out3115_out1            : std_logic;
  SIGNAL Logical_Operator_out3116_out1            : std_logic;
  SIGNAL Logical_Operator_out3117_out1            : std_logic;
  SIGNAL Logical_Operator_out3118_out1            : std_logic;
  SIGNAL Logical_Operator_out3119_out1            : std_logic;
  SIGNAL Logical_Operator_out3120_out1            : std_logic;
  SIGNAL Logical_Operator_out3121_out1            : std_logic;
  SIGNAL Logical_Operator_out3122_out1            : std_logic;
  SIGNAL Logical_Operator_out3123_out1            : std_logic;
  SIGNAL Logical_Operator_out3124_out1            : std_logic;
  SIGNAL Logical_Operator_out3125_out1            : std_logic;
  SIGNAL Logical_Operator_out3126_out1            : std_logic;
  SIGNAL Logical_Operator_out3127_out1            : std_logic;
  SIGNAL Logical_Operator_out3128_out1            : std_logic;
  SIGNAL Logical_Operator_out3129_out1            : std_logic;
  SIGNAL Logical_Operator_out3130_out1            : std_logic;
  SIGNAL Logical_Operator_out3131_out1            : std_logic;
  SIGNAL Logical_Operator_out3132_out1            : std_logic;
  SIGNAL Logical_Operator_out3133_out1            : std_logic;
  SIGNAL Logical_Operator_out3134_out1            : std_logic;
  SIGNAL Logical_Operator_out3135_out1            : std_logic;
  SIGNAL Logical_Operator_out3136_out1            : std_logic;
  SIGNAL Logical_Operator_out3137_out1            : std_logic;
  SIGNAL Logical_Operator_out3138_out1            : std_logic;
  SIGNAL Logical_Operator_out3139_out1            : std_logic;
  SIGNAL Logical_Operator_out3140_out1            : std_logic;
  SIGNAL Logical_Operator_out3141_out1            : std_logic;
  SIGNAL Logical_Operator_out3142_out1            : std_logic;
  SIGNAL Logical_Operator_out3143_out1            : std_logic;
  SIGNAL Logical_Operator_out3144_out1            : std_logic;
  SIGNAL Logical_Operator_out3145_out1            : std_logic;
  SIGNAL Logical_Operator_out3146_out1            : std_logic;
  SIGNAL Logical_Operator_out3147_out1            : std_logic;
  SIGNAL Logical_Operator_out3148_out1            : std_logic;
  SIGNAL Logical_Operator_out3149_out1            : std_logic;
  SIGNAL Logical_Operator_out3150_out1            : std_logic;
  SIGNAL Logical_Operator_out3151_out1            : std_logic;
  SIGNAL Logical_Operator_out3152_out1            : std_logic;
  SIGNAL Logical_Operator_out3153_out1            : std_logic;
  SIGNAL Logical_Operator_out3154_out1            : std_logic;
  SIGNAL Logical_Operator_out3155_out1            : std_logic;
  SIGNAL Logical_Operator_out3156_out1            : std_logic;
  SIGNAL Logical_Operator_out3157_out1            : std_logic;
  SIGNAL Logical_Operator_out3158_out1            : std_logic;
  SIGNAL Logical_Operator_out3159_out1            : std_logic;
  SIGNAL Logical_Operator_out3160_out1            : std_logic;
  SIGNAL Logical_Operator_out3161_out1            : std_logic;
  SIGNAL Logical_Operator_out3162_out1            : std_logic;
  SIGNAL Logical_Operator_out3163_out1            : std_logic;
  SIGNAL Logical_Operator_out3164_out1            : std_logic;
  SIGNAL Logical_Operator_out3165_out1            : std_logic;
  SIGNAL Logical_Operator_out3166_out1            : std_logic;
  SIGNAL Logical_Operator_out3167_out1            : std_logic;
  SIGNAL Logical_Operator_out3168_out1            : std_logic;
  SIGNAL Logical_Operator_out3169_out1            : std_logic;
  SIGNAL Logical_Operator_out3170_out1            : std_logic;
  SIGNAL Logical_Operator_out3171_out1            : std_logic;
  SIGNAL Logical_Operator_out3172_out1            : std_logic;
  SIGNAL Logical_Operator_out3173_out1            : std_logic;
  SIGNAL Logical_Operator_out3174_out1            : std_logic;
  SIGNAL Logical_Operator_out3175_out1            : std_logic;
  SIGNAL Logical_Operator_out3176_out1            : std_logic;
  SIGNAL Logical_Operator_out3177_out1            : std_logic;
  SIGNAL Logical_Operator_out3178_out1            : std_logic;
  SIGNAL Logical_Operator_out3179_out1            : std_logic;
  SIGNAL Logical_Operator_out3180_out1            : std_logic;
  SIGNAL Logical_Operator_out3181_out1            : std_logic;
  SIGNAL Logical_Operator_out3182_out1            : std_logic;
  SIGNAL Logical_Operator_out3183_out1            : std_logic;
  SIGNAL Logical_Operator_out3184_out1            : std_logic;
  SIGNAL Logical_Operator_out3185_out1            : std_logic;
  SIGNAL Logical_Operator_out3186_out1            : std_logic;
  SIGNAL Logical_Operator_out3187_out1            : std_logic;
  SIGNAL Logical_Operator_out3188_out1            : std_logic;
  SIGNAL Logical_Operator_out3189_out1            : std_logic;
  SIGNAL Logical_Operator_out3190_out1            : std_logic;
  SIGNAL Logical_Operator_out3191_out1            : std_logic;
  SIGNAL Logical_Operator_out3192_out1            : std_logic;
  SIGNAL Logical_Operator_out3193_out1            : std_logic;
  SIGNAL Logical_Operator_out3194_out1            : std_logic;
  SIGNAL Logical_Operator_out3195_out1            : std_logic;
  SIGNAL Logical_Operator_out3196_out1            : std_logic;
  SIGNAL Logical_Operator_out3197_out1            : std_logic;
  SIGNAL Logical_Operator_out3198_out1            : std_logic;
  SIGNAL Logical_Operator_out3199_out1            : std_logic;
  SIGNAL Logical_Operator_out3200_out1            : std_logic;
  SIGNAL Logical_Operator_out3201_out1            : std_logic;
  SIGNAL Logical_Operator_out3202_out1            : std_logic;
  SIGNAL Logical_Operator_out3203_out1            : std_logic;
  SIGNAL Logical_Operator_out3204_out1            : std_logic;
  SIGNAL Logical_Operator_out3205_out1            : std_logic;
  SIGNAL Logical_Operator_out3206_out1            : std_logic;
  SIGNAL Logical_Operator_out3207_out1            : std_logic;
  SIGNAL Logical_Operator_out3208_out1            : std_logic;
  SIGNAL Logical_Operator_out3209_out1            : std_logic;
  SIGNAL Logical_Operator_out3210_out1            : std_logic;
  SIGNAL Logical_Operator_out3211_out1            : std_logic;
  SIGNAL Logical_Operator_out3212_out1            : std_logic;
  SIGNAL Logical_Operator_out3213_out1            : std_logic;
  SIGNAL Logical_Operator_out3214_out1            : std_logic;
  SIGNAL Logical_Operator_out3215_out1            : std_logic;
  SIGNAL Logical_Operator_out3216_out1            : std_logic;
  SIGNAL Logical_Operator_out3217_out1            : std_logic;
  SIGNAL Logical_Operator_out3218_out1            : std_logic;
  SIGNAL Logical_Operator_out3219_out1            : std_logic;
  SIGNAL Logical_Operator_out3220_out1            : std_logic;
  SIGNAL Logical_Operator_out3221_out1            : std_logic;
  SIGNAL Logical_Operator_out3222_out1            : std_logic;
  SIGNAL Logical_Operator_out3223_out1            : std_logic;
  SIGNAL Logical_Operator_out3224_out1            : std_logic;
  SIGNAL Logical_Operator_out3225_out1            : std_logic;
  SIGNAL Logical_Operator_out3226_out1            : std_logic;
  SIGNAL Logical_Operator_out3227_out1            : std_logic;
  SIGNAL Logical_Operator_out3228_out1            : std_logic;
  SIGNAL Logical_Operator_out3229_out1            : std_logic;
  SIGNAL Logical_Operator_out3230_out1            : std_logic;
  SIGNAL Logical_Operator_out3231_out1            : std_logic;
  SIGNAL Logical_Operator_out3232_out1            : std_logic;
  SIGNAL Logical_Operator_out3233_out1            : std_logic;
  SIGNAL Logical_Operator_out3234_out1            : std_logic;
  SIGNAL Logical_Operator_out3235_out1            : std_logic;
  SIGNAL Logical_Operator_out3236_out1            : std_logic;
  SIGNAL Logical_Operator_out3237_out1            : std_logic;
  SIGNAL Logical_Operator_out3238_out1            : std_logic;
  SIGNAL Logical_Operator_out3239_out1            : std_logic;
  SIGNAL Logical_Operator_out3240_out1            : std_logic;
  SIGNAL Logical_Operator_out3241_out1            : std_logic;
  SIGNAL Logical_Operator_out3242_out1            : std_logic;
  SIGNAL Logical_Operator_out3243_out1            : std_logic;
  SIGNAL Logical_Operator_out3244_out1            : std_logic;
  SIGNAL Logical_Operator_out3245_out1            : std_logic;
  SIGNAL Logical_Operator_out3246_out1            : std_logic;
  SIGNAL Logical_Operator_out3247_out1            : std_logic;
  SIGNAL Logical_Operator_out3248_out1            : std_logic;
  SIGNAL Logical_Operator_out3249_out1            : std_logic;
  SIGNAL Logical_Operator_out3250_out1            : std_logic;
  SIGNAL Logical_Operator_out3251_out1            : std_logic;
  SIGNAL Logical_Operator_out3252_out1            : std_logic;
  SIGNAL Logical_Operator_out3253_out1            : std_logic;
  SIGNAL Logical_Operator_out3254_out1            : std_logic;
  SIGNAL Logical_Operator_out3255_out1            : std_logic;
  SIGNAL Logical_Operator_out3256_out1            : std_logic;
  SIGNAL Logical_Operator_out3257_out1            : std_logic;
  SIGNAL Logical_Operator_out3258_out1            : std_logic;
  SIGNAL Logical_Operator_out3259_out1            : std_logic;
  SIGNAL Logical_Operator_out3260_out1            : std_logic;
  SIGNAL Logical_Operator_out3261_out1            : std_logic;
  SIGNAL Logical_Operator_out3262_out1            : std_logic;
  SIGNAL Logical_Operator_out3263_out1            : std_logic;
  SIGNAL Logical_Operator_out3264_out1            : std_logic;
  SIGNAL Logical_Operator_out3265_out1            : std_logic;
  SIGNAL Logical_Operator_out3266_out1            : std_logic;
  SIGNAL Logical_Operator_out3267_out1            : std_logic;
  SIGNAL Logical_Operator_out3268_out1            : std_logic;
  SIGNAL Logical_Operator_out3269_out1            : std_logic;
  SIGNAL Logical_Operator_out3270_out1            : std_logic;
  SIGNAL Logical_Operator_out3271_out1            : std_logic;
  SIGNAL Logical_Operator_out3272_out1            : std_logic;
  SIGNAL Logical_Operator_out3273_out1            : std_logic;
  SIGNAL Logical_Operator_out3274_out1            : std_logic;
  SIGNAL Logical_Operator_out3275_out1            : std_logic;
  SIGNAL Logical_Operator_out3276_out1            : std_logic;
  SIGNAL Logical_Operator_out3277_out1            : std_logic;
  SIGNAL Logical_Operator_out3278_out1            : std_logic;
  SIGNAL Logical_Operator_out3279_out1            : std_logic;
  SIGNAL Logical_Operator_out3280_out1            : std_logic;
  SIGNAL Logical_Operator_out3281_out1            : std_logic;
  SIGNAL Logical_Operator_out3282_out1            : std_logic;
  SIGNAL Logical_Operator_out3283_out1            : std_logic;
  SIGNAL Logical_Operator_out3284_out1            : std_logic;
  SIGNAL Logical_Operator_out3285_out1            : std_logic;
  SIGNAL Logical_Operator_out3286_out1            : std_logic;
  SIGNAL Logical_Operator_out3287_out1            : std_logic;
  SIGNAL Logical_Operator_out3288_out1            : std_logic;
  SIGNAL Logical_Operator_out3289_out1            : std_logic;
  SIGNAL Logical_Operator_out3290_out1            : std_logic;
  SIGNAL Logical_Operator_out3291_out1            : std_logic;
  SIGNAL Logical_Operator_out3292_out1            : std_logic;
  SIGNAL Logical_Operator_out3293_out1            : std_logic;
  SIGNAL Logical_Operator_out3294_out1            : std_logic;
  SIGNAL Logical_Operator_out3295_out1            : std_logic;
  SIGNAL Logical_Operator_out3296_out1            : std_logic;
  SIGNAL Logical_Operator_out3297_out1            : std_logic;
  SIGNAL Logical_Operator_out3298_out1            : std_logic;
  SIGNAL Logical_Operator_out3299_out1            : std_logic;
  SIGNAL Logical_Operator_out3300_out1            : std_logic;
  SIGNAL Logical_Operator_out3301_out1            : std_logic;
  SIGNAL Logical_Operator_out3302_out1            : std_logic;
  SIGNAL Logical_Operator_out3303_out1            : std_logic;
  SIGNAL Logical_Operator_out3304_out1            : std_logic;
  SIGNAL Logical_Operator_out3305_out1            : std_logic;
  SIGNAL Logical_Operator_out3306_out1            : std_logic;
  SIGNAL Logical_Operator_out3307_out1            : std_logic;
  SIGNAL Logical_Operator_out3308_out1            : std_logic;
  SIGNAL Logical_Operator_out3309_out1            : std_logic;
  SIGNAL Logical_Operator_out3310_out1            : std_logic;
  SIGNAL Logical_Operator_out3311_out1            : std_logic;
  SIGNAL Logical_Operator_out3312_out1            : std_logic;
  SIGNAL Logical_Operator_out3313_out1            : std_logic;
  SIGNAL Logical_Operator_out3314_out1            : std_logic;
  SIGNAL Logical_Operator_out3315_out1            : std_logic;
  SIGNAL Logical_Operator_out3316_out1            : std_logic;
  SIGNAL Logical_Operator_out3317_out1            : std_logic;
  SIGNAL Logical_Operator_out3318_out1            : std_logic;
  SIGNAL Logical_Operator_out3319_out1            : std_logic;
  SIGNAL Logical_Operator_out3320_out1            : std_logic;
  SIGNAL Logical_Operator_out3321_out1            : std_logic;
  SIGNAL Logical_Operator_out3322_out1            : std_logic;
  SIGNAL Logical_Operator_out3323_out1            : std_logic;
  SIGNAL Logical_Operator_out3324_out1            : std_logic;
  SIGNAL Logical_Operator_out3325_out1            : std_logic;
  SIGNAL Logical_Operator_out3326_out1            : std_logic;
  SIGNAL Logical_Operator_out3327_out1            : std_logic;
  SIGNAL Logical_Operator_out3328_out1            : std_logic;
  SIGNAL Logical_Operator_out3329_out1            : std_logic;
  SIGNAL Logical_Operator_out3330_out1            : std_logic;
  SIGNAL Logical_Operator_out3331_out1            : std_logic;
  SIGNAL Logical_Operator_out3332_out1            : std_logic;
  SIGNAL Logical_Operator_out3333_out1            : std_logic;
  SIGNAL Logical_Operator_out3334_out1            : std_logic;
  SIGNAL Logical_Operator_out3335_out1            : std_logic;
  SIGNAL Logical_Operator_out3336_out1            : std_logic;
  SIGNAL Logical_Operator_out3337_out1            : std_logic;
  SIGNAL Logical_Operator_out3338_out1            : std_logic;
  SIGNAL Logical_Operator_out3339_out1            : std_logic;
  SIGNAL Logical_Operator_out3340_out1            : std_logic;
  SIGNAL Logical_Operator_out3341_out1            : std_logic;
  SIGNAL Logical_Operator_out3342_out1            : std_logic;
  SIGNAL Logical_Operator_out3343_out1            : std_logic;
  SIGNAL Logical_Operator_out3344_out1            : std_logic;
  SIGNAL Logical_Operator_out3345_out1            : std_logic;
  SIGNAL Logical_Operator_out3346_out1            : std_logic;
  SIGNAL Logical_Operator_out3347_out1            : std_logic;
  SIGNAL Logical_Operator_out3348_out1            : std_logic;
  SIGNAL Logical_Operator_out3349_out1            : std_logic;
  SIGNAL Logical_Operator_out3350_out1            : std_logic;
  SIGNAL Logical_Operator_out3351_out1            : std_logic;
  SIGNAL Logical_Operator_out3352_out1            : std_logic;
  SIGNAL Logical_Operator_out3353_out1            : std_logic;
  SIGNAL Logical_Operator_out3354_out1            : std_logic;
  SIGNAL Logical_Operator_out3355_out1            : std_logic;
  SIGNAL Logical_Operator_out3356_out1            : std_logic;
  SIGNAL Logical_Operator_out3357_out1            : std_logic;
  SIGNAL Logical_Operator_out3358_out1            : std_logic;
  SIGNAL Logical_Operator_out3359_out1            : std_logic;
  SIGNAL Logical_Operator_out3360_out1            : std_logic;
  SIGNAL Logical_Operator_out3361_out1            : std_logic;
  SIGNAL Logical_Operator_out3362_out1            : std_logic;
  SIGNAL Logical_Operator_out3363_out1            : std_logic;
  SIGNAL Logical_Operator_out3364_out1            : std_logic;
  SIGNAL Logical_Operator_out3365_out1            : std_logic;
  SIGNAL Logical_Operator_out3366_out1            : std_logic;
  SIGNAL Logical_Operator_out3367_out1            : std_logic;
  SIGNAL Logical_Operator_out3368_out1            : std_logic;
  SIGNAL Logical_Operator_out3369_out1            : std_logic;
  SIGNAL Logical_Operator_out3370_out1            : std_logic;
  SIGNAL Logical_Operator_out3371_out1            : std_logic;
  SIGNAL Logical_Operator_out3372_out1            : std_logic;
  SIGNAL Logical_Operator_out3373_out1            : std_logic;
  SIGNAL Logical_Operator_out3374_out1            : std_logic;
  SIGNAL Logical_Operator_out3375_out1            : std_logic;
  SIGNAL Logical_Operator_out3376_out1            : std_logic;
  SIGNAL Logical_Operator_out3377_out1            : std_logic;
  SIGNAL Logical_Operator_out3378_out1            : std_logic;
  SIGNAL Logical_Operator_out3379_out1            : std_logic;
  SIGNAL Logical_Operator_out3380_out1            : std_logic;
  SIGNAL Logical_Operator_out3381_out1            : std_logic;
  SIGNAL Logical_Operator_out3382_out1            : std_logic;
  SIGNAL Logical_Operator_out3383_out1            : std_logic;
  SIGNAL Logical_Operator_out3384_out1            : std_logic;
  SIGNAL Logical_Operator_out3385_out1            : std_logic;
  SIGNAL Logical_Operator_out3386_out1            : std_logic;
  SIGNAL Logical_Operator_out3387_out1            : std_logic;
  SIGNAL Logical_Operator_out3388_out1            : std_logic;
  SIGNAL Logical_Operator_out3389_out1            : std_logic;
  SIGNAL Logical_Operator_out3390_out1            : std_logic;
  SIGNAL Logical_Operator_out3391_out1            : std_logic;
  SIGNAL Logical_Operator_out3392_out1            : std_logic;
  SIGNAL Logical_Operator_out3393_out1            : std_logic;
  SIGNAL Logical_Operator_out3394_out1            : std_logic;
  SIGNAL Logical_Operator_out3395_out1            : std_logic;
  SIGNAL Logical_Operator_out3396_out1            : std_logic;
  SIGNAL Logical_Operator_out3397_out1            : std_logic;
  SIGNAL Logical_Operator_out3398_out1            : std_logic;
  SIGNAL Logical_Operator_out3399_out1            : std_logic;
  SIGNAL Logical_Operator_out3400_out1            : std_logic;
  SIGNAL Logical_Operator_out3401_out1            : std_logic;
  SIGNAL Logical_Operator_out3402_out1            : std_logic;
  SIGNAL Logical_Operator_out3403_out1            : std_logic;
  SIGNAL Logical_Operator_out3404_out1            : std_logic;
  SIGNAL Logical_Operator_out3405_out1            : std_logic;
  SIGNAL Logical_Operator_out3406_out1            : std_logic;
  SIGNAL Logical_Operator_out3407_out1            : std_logic;
  SIGNAL Logical_Operator_out3408_out1            : std_logic;
  SIGNAL Logical_Operator_out3409_out1            : std_logic;
  SIGNAL Logical_Operator_out3410_out1            : std_logic;
  SIGNAL Logical_Operator_out3411_out1            : std_logic;
  SIGNAL Logical_Operator_out3412_out1            : std_logic;
  SIGNAL Logical_Operator_out3413_out1            : std_logic;
  SIGNAL Logical_Operator_out3414_out1            : std_logic;
  SIGNAL Logical_Operator_out3415_out1            : std_logic;
  SIGNAL Logical_Operator_out3416_out1            : std_logic;
  SIGNAL Logical_Operator_out3417_out1            : std_logic;
  SIGNAL Logical_Operator_out3418_out1            : std_logic;
  SIGNAL Logical_Operator_out3419_out1            : std_logic;
  SIGNAL Logical_Operator_out3420_out1            : std_logic;
  SIGNAL Logical_Operator_out3421_out1            : std_logic;
  SIGNAL Logical_Operator_out3422_out1            : std_logic;
  SIGNAL Logical_Operator_out3423_out1            : std_logic;
  SIGNAL Logical_Operator_out3424_out1            : std_logic;
  SIGNAL Logical_Operator_out3425_out1            : std_logic;
  SIGNAL Logical_Operator_out3426_out1            : std_logic;
  SIGNAL Logical_Operator_out3427_out1            : std_logic;
  SIGNAL Logical_Operator_out3428_out1            : std_logic;
  SIGNAL Logical_Operator_out3429_out1            : std_logic;
  SIGNAL Logical_Operator_out3430_out1            : std_logic;
  SIGNAL Logical_Operator_out3431_out1            : std_logic;
  SIGNAL Logical_Operator_out3432_out1            : std_logic;
  SIGNAL Logical_Operator_out3433_out1            : std_logic;
  SIGNAL Logical_Operator_out3434_out1            : std_logic;
  SIGNAL Logical_Operator_out3435_out1            : std_logic;
  SIGNAL Logical_Operator_out3436_out1            : std_logic;
  SIGNAL Logical_Operator_out3437_out1            : std_logic;
  SIGNAL Logical_Operator_out3438_out1            : std_logic;
  SIGNAL Logical_Operator_out3439_out1            : std_logic;
  SIGNAL Logical_Operator_out3440_out1            : std_logic;
  SIGNAL Logical_Operator_out3441_out1            : std_logic;
  SIGNAL Logical_Operator_out3442_out1            : std_logic;
  SIGNAL Logical_Operator_out3443_out1            : std_logic;
  SIGNAL Logical_Operator_out3444_out1            : std_logic;
  SIGNAL Logical_Operator_out3445_out1            : std_logic;
  SIGNAL Logical_Operator_out3446_out1            : std_logic;
  SIGNAL Logical_Operator_out3447_out1            : std_logic;
  SIGNAL Logical_Operator_out3448_out1            : std_logic;
  SIGNAL Logical_Operator_out3449_out1            : std_logic;
  SIGNAL Logical_Operator_out3450_out1            : std_logic;
  SIGNAL Logical_Operator_out3451_out1            : std_logic;
  SIGNAL Logical_Operator_out3452_out1            : std_logic;
  SIGNAL Logical_Operator_out3453_out1            : std_logic;
  SIGNAL Logical_Operator_out3454_out1            : std_logic;
  SIGNAL Logical_Operator_out3455_out1            : std_logic;
  SIGNAL Logical_Operator_out3456_out1            : std_logic;
  SIGNAL Logical_Operator_out3457_out1            : std_logic;
  SIGNAL Logical_Operator_out3458_out1            : std_logic;
  SIGNAL Logical_Operator_out3459_out1            : std_logic;
  SIGNAL Logical_Operator_out3460_out1            : std_logic;
  SIGNAL Logical_Operator_out3461_out1            : std_logic;
  SIGNAL Logical_Operator_out3462_out1            : std_logic;
  SIGNAL Logical_Operator_out3463_out1            : std_logic;
  SIGNAL Logical_Operator_out3464_out1            : std_logic;
  SIGNAL Logical_Operator_out3465_out1            : std_logic;
  SIGNAL Logical_Operator_out3466_out1            : std_logic;
  SIGNAL Logical_Operator_out3467_out1            : std_logic;
  SIGNAL Logical_Operator_out3468_out1            : std_logic;
  SIGNAL Logical_Operator_out3469_out1            : std_logic;
  SIGNAL Logical_Operator_out3470_out1            : std_logic;
  SIGNAL Logical_Operator_out3471_out1            : std_logic;
  SIGNAL Logical_Operator_out3472_out1            : std_logic;
  SIGNAL Logical_Operator_out3473_out1            : std_logic;
  SIGNAL Logical_Operator_out3474_out1            : std_logic;
  SIGNAL Logical_Operator_out3475_out1            : std_logic;
  SIGNAL Logical_Operator_out3476_out1            : std_logic;
  SIGNAL Logical_Operator_out3477_out1            : std_logic;
  SIGNAL Logical_Operator_out3478_out1            : std_logic;
  SIGNAL Logical_Operator_out3479_out1            : std_logic;
  SIGNAL Logical_Operator_out3480_out1            : std_logic;
  SIGNAL Logical_Operator_out3481_out1            : std_logic;
  SIGNAL Logical_Operator_out3482_out1            : std_logic;
  SIGNAL Logical_Operator_out3483_out1            : std_logic;
  SIGNAL Logical_Operator_out3484_out1            : std_logic;
  SIGNAL Logical_Operator_out3485_out1            : std_logic;
  SIGNAL Logical_Operator_out3486_out1            : std_logic;
  SIGNAL Logical_Operator_out3487_out1            : std_logic;
  SIGNAL Logical_Operator_out3488_out1            : std_logic;
  SIGNAL Logical_Operator_out3489_out1            : std_logic;
  SIGNAL Logical_Operator_out3490_out1            : std_logic;
  SIGNAL Logical_Operator_out3491_out1            : std_logic;
  SIGNAL Logical_Operator_out3492_out1            : std_logic;
  SIGNAL Logical_Operator_out3493_out1            : std_logic;
  SIGNAL Logical_Operator_out3494_out1            : std_logic;
  SIGNAL Logical_Operator_out3495_out1            : std_logic;
  SIGNAL Logical_Operator_out3496_out1            : std_logic;
  SIGNAL Logical_Operator_out3497_out1            : std_logic;
  SIGNAL Logical_Operator_out3498_out1            : std_logic;
  SIGNAL Logical_Operator_out3499_out1            : std_logic;
  SIGNAL Logical_Operator_out3500_out1            : std_logic;
  SIGNAL Logical_Operator_out3501_out1            : std_logic;
  SIGNAL Logical_Operator_out3502_out1            : std_logic;
  SIGNAL Logical_Operator_out3503_out1            : std_logic;
  SIGNAL Logical_Operator_out3504_out1            : std_logic;
  SIGNAL Logical_Operator_out3505_out1            : std_logic;
  SIGNAL Logical_Operator_out3506_out1            : std_logic;
  SIGNAL Logical_Operator_out3507_out1            : std_logic;
  SIGNAL Logical_Operator_out3508_out1            : std_logic;
  SIGNAL Logical_Operator_out3509_out1            : std_logic;
  SIGNAL Logical_Operator_out3510_out1            : std_logic;
  SIGNAL Logical_Operator_out3511_out1            : std_logic;
  SIGNAL Logical_Operator_out3512_out1            : std_logic;
  SIGNAL Logical_Operator_out3513_out1            : std_logic;
  SIGNAL Logical_Operator_out3514_out1            : std_logic;
  SIGNAL Logical_Operator_out3515_out1            : std_logic;
  SIGNAL Logical_Operator_out3516_out1            : std_logic;
  SIGNAL Logical_Operator_out3517_out1            : std_logic;
  SIGNAL Logical_Operator_out3518_out1            : std_logic;
  SIGNAL Logical_Operator_out3519_out1            : std_logic;
  SIGNAL Logical_Operator_out3520_out1            : std_logic;
  SIGNAL Logical_Operator_out3521_out1            : std_logic;
  SIGNAL Logical_Operator_out3522_out1            : std_logic;
  SIGNAL Logical_Operator_out3523_out1            : std_logic;
  SIGNAL Logical_Operator_out3524_out1            : std_logic;
  SIGNAL Logical_Operator_out3525_out1            : std_logic;
  SIGNAL Logical_Operator_out3526_out1            : std_logic;
  SIGNAL Logical_Operator_out3527_out1            : std_logic;
  SIGNAL Logical_Operator_out3528_out1            : std_logic;
  SIGNAL Logical_Operator_out3529_out1            : std_logic;
  SIGNAL Logical_Operator_out3530_out1            : std_logic;
  SIGNAL Logical_Operator_out3531_out1            : std_logic;
  SIGNAL Logical_Operator_out3532_out1            : std_logic;
  SIGNAL Logical_Operator_out3533_out1            : std_logic;
  SIGNAL Logical_Operator_out3534_out1            : std_logic;
  SIGNAL Logical_Operator_out3535_out1            : std_logic;
  SIGNAL Logical_Operator_out3536_out1            : std_logic;
  SIGNAL Logical_Operator_out3537_out1            : std_logic;
  SIGNAL Logical_Operator_out3538_out1            : std_logic;
  SIGNAL Logical_Operator_out3539_out1            : std_logic;
  SIGNAL Logical_Operator_out3540_out1            : std_logic;
  SIGNAL Logical_Operator_out3541_out1            : std_logic;
  SIGNAL Logical_Operator_out3542_out1            : std_logic;
  SIGNAL Logical_Operator_out3543_out1            : std_logic;
  SIGNAL Logical_Operator_out3544_out1            : std_logic;
  SIGNAL Logical_Operator_out3545_out1            : std_logic;
  SIGNAL Logical_Operator_out3546_out1            : std_logic;
  SIGNAL Logical_Operator_out3547_out1            : std_logic;
  SIGNAL Logical_Operator_out3548_out1            : std_logic;
  SIGNAL Logical_Operator_out3549_out1            : std_logic;
  SIGNAL Logical_Operator_out3550_out1            : std_logic;
  SIGNAL Logical_Operator_out3551_out1            : std_logic;
  SIGNAL Logical_Operator_out3552_out1            : std_logic;
  SIGNAL Logical_Operator_out3553_out1            : std_logic;
  SIGNAL Logical_Operator_out3554_out1            : std_logic;
  SIGNAL Logical_Operator_out3555_out1            : std_logic;
  SIGNAL Logical_Operator_out3556_out1            : std_logic;
  SIGNAL Logical_Operator_out3557_out1            : std_logic;
  SIGNAL Logical_Operator_out3558_out1            : std_logic;
  SIGNAL Logical_Operator_out3559_out1            : std_logic;
  SIGNAL Logical_Operator_out3560_out1            : std_logic;
  SIGNAL Logical_Operator_out3561_out1            : std_logic;
  SIGNAL Logical_Operator_out3562_out1            : std_logic;
  SIGNAL Logical_Operator_out3563_out1            : std_logic;
  SIGNAL Logical_Operator_out3564_out1            : std_logic;
  SIGNAL Logical_Operator_out3565_out1            : std_logic;
  SIGNAL Logical_Operator_out3566_out1            : std_logic;
  SIGNAL Logical_Operator_out3567_out1            : std_logic;
  SIGNAL Logical_Operator_out3568_out1            : std_logic;
  SIGNAL Logical_Operator_out3569_out1            : std_logic;
  SIGNAL Logical_Operator_out3570_out1            : std_logic;
  SIGNAL Logical_Operator_out3571_out1            : std_logic;
  SIGNAL Logical_Operator_out3572_out1            : std_logic;
  SIGNAL Logical_Operator_out3573_out1            : std_logic;
  SIGNAL Logical_Operator_out3574_out1            : std_logic;
  SIGNAL Logical_Operator_out3575_out1            : std_logic;
  SIGNAL Logical_Operator_out3576_out1            : std_logic;
  SIGNAL Logical_Operator_out3577_out1            : std_logic;
  SIGNAL Logical_Operator_out3578_out1            : std_logic;
  SIGNAL Logical_Operator_out3579_out1            : std_logic;
  SIGNAL Logical_Operator_out3580_out1            : std_logic;
  SIGNAL Logical_Operator_out3581_out1            : std_logic;
  SIGNAL Logical_Operator_out3582_out1            : std_logic;
  SIGNAL Logical_Operator_out3583_out1            : std_logic;
  SIGNAL Logical_Operator_out3584_out1            : std_logic;
  SIGNAL Logical_Operator_out3585_out1            : std_logic;
  SIGNAL Logical_Operator_out3586_out1            : std_logic;
  SIGNAL Logical_Operator_out3587_out1            : std_logic;
  SIGNAL Logical_Operator_out3588_out1            : std_logic;
  SIGNAL Logical_Operator_out3589_out1            : std_logic;
  SIGNAL Logical_Operator_out3590_out1            : std_logic;
  SIGNAL Logical_Operator_out3591_out1            : std_logic;
  SIGNAL Logical_Operator_out3592_out1            : std_logic;
  SIGNAL Logical_Operator_out3593_out1            : std_logic;
  SIGNAL Logical_Operator_out3594_out1            : std_logic;
  SIGNAL Logical_Operator_out3595_out1            : std_logic;
  SIGNAL Logical_Operator_out3596_out1            : std_logic;
  SIGNAL Logical_Operator_out3597_out1            : std_logic;
  SIGNAL Logical_Operator_out3598_out1            : std_logic;
  SIGNAL Logical_Operator_out3599_out1            : std_logic;
  SIGNAL Logical_Operator_out3600_out1            : std_logic;
  SIGNAL Logical_Operator_out3601_out1            : std_logic;
  SIGNAL Logical_Operator_out3602_out1            : std_logic;
  SIGNAL Logical_Operator_out3603_out1            : std_logic;
  SIGNAL Logical_Operator_out3604_out1            : std_logic;
  SIGNAL Logical_Operator_out3605_out1            : std_logic;
  SIGNAL Logical_Operator_out3606_out1            : std_logic;
  SIGNAL Logical_Operator_out3607_out1            : std_logic;
  SIGNAL Logical_Operator_out3608_out1            : std_logic;
  SIGNAL Logical_Operator_out3609_out1            : std_logic;
  SIGNAL Logical_Operator_out3610_out1            : std_logic;
  SIGNAL Logical_Operator_out3611_out1            : std_logic;
  SIGNAL Logical_Operator_out3612_out1            : std_logic;
  SIGNAL Logical_Operator_out3613_out1            : std_logic;
  SIGNAL Logical_Operator_out3614_out1            : std_logic;
  SIGNAL Logical_Operator_out3615_out1            : std_logic;
  SIGNAL Logical_Operator_out3616_out1            : std_logic;
  SIGNAL Logical_Operator_out3617_out1            : std_logic;
  SIGNAL Logical_Operator_out3618_out1            : std_logic;
  SIGNAL Logical_Operator_out3619_out1            : std_logic;
  SIGNAL Logical_Operator_out3620_out1            : std_logic;
  SIGNAL Logical_Operator_out3621_out1            : std_logic;
  SIGNAL Logical_Operator_out3622_out1            : std_logic;
  SIGNAL Logical_Operator_out3623_out1            : std_logic;
  SIGNAL Logical_Operator_out3624_out1            : std_logic;
  SIGNAL Logical_Operator_out3625_out1            : std_logic;
  SIGNAL Logical_Operator_out3626_out1            : std_logic;
  SIGNAL Logical_Operator_out3627_out1            : std_logic;
  SIGNAL Logical_Operator_out3628_out1            : std_logic;
  SIGNAL Logical_Operator_out3629_out1            : std_logic;
  SIGNAL Logical_Operator_out3630_out1            : std_logic;
  SIGNAL Logical_Operator_out3631_out1            : std_logic;
  SIGNAL Logical_Operator_out3632_out1            : std_logic;
  SIGNAL Logical_Operator_out3633_out1            : std_logic;
  SIGNAL Logical_Operator_out3634_out1            : std_logic;
  SIGNAL Logical_Operator_out3635_out1            : std_logic;
  SIGNAL Logical_Operator_out3636_out1            : std_logic;
  SIGNAL Logical_Operator_out3637_out1            : std_logic;
  SIGNAL Logical_Operator_out3638_out1            : std_logic;
  SIGNAL Logical_Operator_out3639_out1            : std_logic;
  SIGNAL Logical_Operator_out3640_out1            : std_logic;
  SIGNAL Logical_Operator_out3641_out1            : std_logic;
  SIGNAL Logical_Operator_out3642_out1            : std_logic;
  SIGNAL Logical_Operator_out3643_out1            : std_logic;
  SIGNAL Logical_Operator_out3644_out1            : std_logic;
  SIGNAL Logical_Operator_out3645_out1            : std_logic;
  SIGNAL Logical_Operator_out3646_out1            : std_logic;
  SIGNAL Logical_Operator_out3647_out1            : std_logic;
  SIGNAL Logical_Operator_out3648_out1            : std_logic;
  SIGNAL Logical_Operator_out3649_out1            : std_logic;
  SIGNAL Logical_Operator_out3650_out1            : std_logic;
  SIGNAL Logical_Operator_out3651_out1            : std_logic;
  SIGNAL Logical_Operator_out3652_out1            : std_logic;
  SIGNAL Logical_Operator_out3653_out1            : std_logic;
  SIGNAL Logical_Operator_out3654_out1            : std_logic;
  SIGNAL Logical_Operator_out3655_out1            : std_logic;
  SIGNAL Logical_Operator_out3656_out1            : std_logic;
  SIGNAL Logical_Operator_out3657_out1            : std_logic;
  SIGNAL Logical_Operator_out3658_out1            : std_logic;
  SIGNAL Logical_Operator_out3659_out1            : std_logic;
  SIGNAL Logical_Operator_out3660_out1            : std_logic;
  SIGNAL Logical_Operator_out3661_out1            : std_logic;
  SIGNAL Logical_Operator_out3662_out1            : std_logic;
  SIGNAL Logical_Operator_out3663_out1            : std_logic;
  SIGNAL Logical_Operator_out3664_out1            : std_logic;
  SIGNAL Logical_Operator_out3665_out1            : std_logic;
  SIGNAL Logical_Operator_out3666_out1            : std_logic;
  SIGNAL Logical_Operator_out3667_out1            : std_logic;
  SIGNAL Logical_Operator_out3668_out1            : std_logic;
  SIGNAL Logical_Operator_out3669_out1            : std_logic;
  SIGNAL Logical_Operator_out3670_out1            : std_logic;
  SIGNAL Logical_Operator_out3671_out1            : std_logic;
  SIGNAL Logical_Operator_out3672_out1            : std_logic;
  SIGNAL Logical_Operator_out3673_out1            : std_logic;
  SIGNAL Logical_Operator_out3674_out1            : std_logic;
  SIGNAL Logical_Operator_out3675_out1            : std_logic;
  SIGNAL Logical_Operator_out3676_out1            : std_logic;
  SIGNAL Logical_Operator_out3677_out1            : std_logic;
  SIGNAL Logical_Operator_out3678_out1            : std_logic;
  SIGNAL Logical_Operator_out3679_out1            : std_logic;
  SIGNAL Logical_Operator_out3680_out1            : std_logic;
  SIGNAL Logical_Operator_out3681_out1            : std_logic;
  SIGNAL Logical_Operator_out3682_out1            : std_logic;
  SIGNAL Logical_Operator_out3683_out1            : std_logic;
  SIGNAL Logical_Operator_out3684_out1            : std_logic;
  SIGNAL Logical_Operator_out3685_out1            : std_logic;
  SIGNAL Logical_Operator_out3686_out1            : std_logic;
  SIGNAL Logical_Operator_out3687_out1            : std_logic;
  SIGNAL Logical_Operator_out3688_out1            : std_logic;
  SIGNAL Logical_Operator_out3689_out1            : std_logic;
  SIGNAL Logical_Operator_out3690_out1            : std_logic;
  SIGNAL Logical_Operator_out3691_out1            : std_logic;
  SIGNAL Logical_Operator_out3692_out1            : std_logic;
  SIGNAL Logical_Operator_out3693_out1            : std_logic;
  SIGNAL Logical_Operator_out3694_out1            : std_logic;
  SIGNAL Logical_Operator_out3695_out1            : std_logic;
  SIGNAL Logical_Operator_out3696_out1            : std_logic;
  SIGNAL Logical_Operator_out3697_out1            : std_logic;
  SIGNAL Logical_Operator_out3698_out1            : std_logic;
  SIGNAL Logical_Operator_out3699_out1            : std_logic;
  SIGNAL Logical_Operator_out3700_out1            : std_logic;
  SIGNAL Logical_Operator_out3701_out1            : std_logic;
  SIGNAL Logical_Operator_out3702_out1            : std_logic;
  SIGNAL Logical_Operator_out3703_out1            : std_logic;
  SIGNAL Logical_Operator_out3704_out1            : std_logic;
  SIGNAL Logical_Operator_out3705_out1            : std_logic;
  SIGNAL Logical_Operator_out3706_out1            : std_logic;
  SIGNAL Logical_Operator_out3707_out1            : std_logic;
  SIGNAL Logical_Operator_out3708_out1            : std_logic;
  SIGNAL Logical_Operator_out3709_out1            : std_logic;
  SIGNAL Logical_Operator_out3710_out1            : std_logic;
  SIGNAL Logical_Operator_out3711_out1            : std_logic;
  SIGNAL Logical_Operator_out3712_out1            : std_logic;
  SIGNAL Logical_Operator_out3713_out1            : std_logic;
  SIGNAL Logical_Operator_out3714_out1            : std_logic;
  SIGNAL Logical_Operator_out3715_out1            : std_logic;
  SIGNAL Logical_Operator_out3716_out1            : std_logic;
  SIGNAL Logical_Operator_out3717_out1            : std_logic;
  SIGNAL Logical_Operator_out3718_out1            : std_logic;
  SIGNAL Logical_Operator_out3719_out1            : std_logic;
  SIGNAL Logical_Operator_out3720_out1            : std_logic;
  SIGNAL Logical_Operator_out3721_out1            : std_logic;
  SIGNAL Logical_Operator_out3722_out1            : std_logic;
  SIGNAL Logical_Operator_out3723_out1            : std_logic;
  SIGNAL Logical_Operator_out3724_out1            : std_logic;
  SIGNAL Logical_Operator_out3725_out1            : std_logic;
  SIGNAL Logical_Operator_out3726_out1            : std_logic;
  SIGNAL Logical_Operator_out3727_out1            : std_logic;
  SIGNAL Logical_Operator_out3728_out1            : std_logic;
  SIGNAL Logical_Operator_out3729_out1            : std_logic;
  SIGNAL Logical_Operator_out3730_out1            : std_logic;
  SIGNAL Logical_Operator_out3731_out1            : std_logic;
  SIGNAL Logical_Operator_out3732_out1            : std_logic;
  SIGNAL Logical_Operator_out3733_out1            : std_logic;
  SIGNAL Logical_Operator_out3734_out1            : std_logic;
  SIGNAL Logical_Operator_out3735_out1            : std_logic;
  SIGNAL Logical_Operator_out3736_out1            : std_logic;
  SIGNAL Logical_Operator_out3737_out1            : std_logic;
  SIGNAL Logical_Operator_out3738_out1            : std_logic;
  SIGNAL Logical_Operator_out3739_out1            : std_logic;
  SIGNAL Logical_Operator_out3740_out1            : std_logic;
  SIGNAL Logical_Operator_out3741_out1            : std_logic;
  SIGNAL Logical_Operator_out3742_out1            : std_logic;
  SIGNAL Logical_Operator_out3743_out1            : std_logic;
  SIGNAL Logical_Operator_out3744_out1            : std_logic;
  SIGNAL Logical_Operator_out3745_out1            : std_logic;
  SIGNAL Logical_Operator_out3746_out1            : std_logic;
  SIGNAL Logical_Operator_out3747_out1            : std_logic;
  SIGNAL Logical_Operator_out3748_out1            : std_logic;
  SIGNAL Logical_Operator_out3749_out1            : std_logic;
  SIGNAL Logical_Operator_out3750_out1            : std_logic;
  SIGNAL Logical_Operator_out3751_out1            : std_logic;
  SIGNAL Logical_Operator_out3752_out1            : std_logic;
  SIGNAL Logical_Operator_out3753_out1            : std_logic;
  SIGNAL Logical_Operator_out3754_out1            : std_logic;
  SIGNAL Logical_Operator_out3755_out1            : std_logic;
  SIGNAL Logical_Operator_out3756_out1            : std_logic;
  SIGNAL Logical_Operator_out3757_out1            : std_logic;
  SIGNAL Logical_Operator_out3758_out1            : std_logic;
  SIGNAL Logical_Operator_out3759_out1            : std_logic;
  SIGNAL Logical_Operator_out3760_out1            : std_logic;
  SIGNAL Logical_Operator_out3761_out1            : std_logic;
  SIGNAL Logical_Operator_out3762_out1            : std_logic;
  SIGNAL Logical_Operator_out3763_out1            : std_logic;
  SIGNAL Logical_Operator_out3764_out1            : std_logic;
  SIGNAL Logical_Operator_out3765_out1            : std_logic;
  SIGNAL Logical_Operator_out3766_out1            : std_logic;
  SIGNAL Logical_Operator_out3767_out1            : std_logic;
  SIGNAL Logical_Operator_out3768_out1            : std_logic;
  SIGNAL Logical_Operator_out3769_out1            : std_logic;
  SIGNAL Logical_Operator_out3770_out1            : std_logic;
  SIGNAL Logical_Operator_out3771_out1            : std_logic;
  SIGNAL Logical_Operator_out3772_out1            : std_logic;
  SIGNAL Logical_Operator_out3773_out1            : std_logic;
  SIGNAL Logical_Operator_out3774_out1            : std_logic;
  SIGNAL Logical_Operator_out3775_out1            : std_logic;
  SIGNAL Logical_Operator_out3776_out1            : std_logic;
  SIGNAL Logical_Operator_out3777_out1            : std_logic;
  SIGNAL Logical_Operator_out3778_out1            : std_logic;
  SIGNAL Logical_Operator_out3779_out1            : std_logic;
  SIGNAL Logical_Operator_out3780_out1            : std_logic;
  SIGNAL Logical_Operator_out3781_out1            : std_logic;
  SIGNAL Logical_Operator_out3782_out1            : std_logic;
  SIGNAL Logical_Operator_out3783_out1            : std_logic;
  SIGNAL Logical_Operator_out3784_out1            : std_logic;
  SIGNAL Logical_Operator_out3785_out1            : std_logic;
  SIGNAL Logical_Operator_out3786_out1            : std_logic;
  SIGNAL Logical_Operator_out3787_out1            : std_logic;
  SIGNAL Logical_Operator_out3788_out1            : std_logic;
  SIGNAL Logical_Operator_out3789_out1            : std_logic;
  SIGNAL Logical_Operator_out3790_out1            : std_logic;
  SIGNAL Logical_Operator_out3791_out1            : std_logic;
  SIGNAL Logical_Operator_out3792_out1            : std_logic;
  SIGNAL Logical_Operator_out3793_out1            : std_logic;
  SIGNAL Logical_Operator_out3794_out1            : std_logic;
  SIGNAL Logical_Operator_out3795_out1            : std_logic;
  SIGNAL Logical_Operator_out3796_out1            : std_logic;
  SIGNAL Logical_Operator_out3797_out1            : std_logic;
  SIGNAL Logical_Operator_out3798_out1            : std_logic;
  SIGNAL Logical_Operator_out3799_out1            : std_logic;
  SIGNAL Logical_Operator_out3800_out1            : std_logic;
  SIGNAL Logical_Operator_out3801_out1            : std_logic;
  SIGNAL Logical_Operator_out3802_out1            : std_logic;
  SIGNAL Logical_Operator_out3803_out1            : std_logic;
  SIGNAL Logical_Operator_out3804_out1            : std_logic;
  SIGNAL Logical_Operator_out3805_out1            : std_logic;
  SIGNAL Logical_Operator_out3806_out1            : std_logic;
  SIGNAL Logical_Operator_out3807_out1            : std_logic;
  SIGNAL Logical_Operator_out3808_out1            : std_logic;
  SIGNAL Logical_Operator_out3809_out1            : std_logic;
  SIGNAL Logical_Operator_out3810_out1            : std_logic;
  SIGNAL Logical_Operator_out3811_out1            : std_logic;
  SIGNAL Logical_Operator_out3812_out1            : std_logic;
  SIGNAL Logical_Operator_out3813_out1            : std_logic;
  SIGNAL Logical_Operator_out3814_out1            : std_logic;
  SIGNAL Logical_Operator_out3815_out1            : std_logic;
  SIGNAL Logical_Operator_out3816_out1            : std_logic;
  SIGNAL Logical_Operator_out3817_out1            : std_logic;
  SIGNAL Logical_Operator_out3818_out1            : std_logic;
  SIGNAL Logical_Operator_out3819_out1            : std_logic;
  SIGNAL Logical_Operator_out3820_out1            : std_logic;
  SIGNAL Logical_Operator_out3821_out1            : std_logic;
  SIGNAL Logical_Operator_out3822_out1            : std_logic;
  SIGNAL Logical_Operator_out3823_out1            : std_logic;
  SIGNAL Logical_Operator_out3824_out1            : std_logic;
  SIGNAL Logical_Operator_out3825_out1            : std_logic;
  SIGNAL Logical_Operator_out3826_out1            : std_logic;
  SIGNAL Logical_Operator_out3827_out1            : std_logic;
  SIGNAL Logical_Operator_out3828_out1            : std_logic;
  SIGNAL Logical_Operator_out3829_out1            : std_logic;
  SIGNAL Logical_Operator_out3830_out1            : std_logic;
  SIGNAL Logical_Operator_out3831_out1            : std_logic;
  SIGNAL Logical_Operator_out3832_out1            : std_logic;
  SIGNAL Logical_Operator_out3833_out1            : std_logic;
  SIGNAL Logical_Operator_out3834_out1            : std_logic;
  SIGNAL Logical_Operator_out3835_out1            : std_logic;
  SIGNAL Logical_Operator_out3836_out1            : std_logic;
  SIGNAL Logical_Operator_out3837_out1            : std_logic;
  SIGNAL Logical_Operator_out3838_out1            : std_logic;
  SIGNAL Logical_Operator_out3839_out1            : std_logic;
  SIGNAL Logical_Operator_out3840_out1            : std_logic;
  SIGNAL Logical_Operator_out3841_out1            : std_logic;
  SIGNAL Logical_Operator_out3842_out1            : std_logic;
  SIGNAL Logical_Operator_out3843_out1            : std_logic;
  SIGNAL Logical_Operator_out3844_out1            : std_logic;
  SIGNAL Logical_Operator_out3845_out1            : std_logic;
  SIGNAL Logical_Operator_out3846_out1            : std_logic;
  SIGNAL Logical_Operator_out3847_out1            : std_logic;
  SIGNAL Logical_Operator_out3848_out1            : std_logic;
  SIGNAL Logical_Operator_out3849_out1            : std_logic;
  SIGNAL Logical_Operator_out3850_out1            : std_logic;
  SIGNAL Logical_Operator_out3851_out1            : std_logic;
  SIGNAL Logical_Operator_out3852_out1            : std_logic;
  SIGNAL Logical_Operator_out3853_out1            : std_logic;
  SIGNAL Logical_Operator_out3854_out1            : std_logic;
  SIGNAL Logical_Operator_out3855_out1            : std_logic;
  SIGNAL Logical_Operator_out3856_out1            : std_logic;
  SIGNAL Logical_Operator_out3857_out1            : std_logic;
  SIGNAL Logical_Operator_out3858_out1            : std_logic;
  SIGNAL Logical_Operator_out3859_out1            : std_logic;
  SIGNAL Logical_Operator_out3860_out1            : std_logic;
  SIGNAL Logical_Operator_out3861_out1            : std_logic;
  SIGNAL Logical_Operator_out3862_out1            : std_logic;
  SIGNAL Logical_Operator_out3863_out1            : std_logic;
  SIGNAL Logical_Operator_out3864_out1            : std_logic;
  SIGNAL Logical_Operator_out3865_out1            : std_logic;
  SIGNAL Logical_Operator_out3866_out1            : std_logic;
  SIGNAL Logical_Operator_out3867_out1            : std_logic;
  SIGNAL Logical_Operator_out3868_out1            : std_logic;
  SIGNAL Logical_Operator_out3869_out1            : std_logic;
  SIGNAL Logical_Operator_out3870_out1            : std_logic;
  SIGNAL Logical_Operator_out3871_out1            : std_logic;
  SIGNAL Logical_Operator_out3872_out1            : std_logic;
  SIGNAL Logical_Operator_out3873_out1            : std_logic;
  SIGNAL Logical_Operator_out3874_out1            : std_logic;
  SIGNAL Logical_Operator_out3875_out1            : std_logic;
  SIGNAL Logical_Operator_out3876_out1            : std_logic;
  SIGNAL Logical_Operator_out3877_out1            : std_logic;
  SIGNAL Logical_Operator_out3878_out1            : std_logic;
  SIGNAL Logical_Operator_out3879_out1            : std_logic;
  SIGNAL Logical_Operator_out3880_out1            : std_logic;
  SIGNAL Logical_Operator_out3881_out1            : std_logic;
  SIGNAL Logical_Operator_out3882_out1            : std_logic;
  SIGNAL Logical_Operator_out3883_out1            : std_logic;
  SIGNAL Logical_Operator_out3884_out1            : std_logic;
  SIGNAL Logical_Operator_out3885_out1            : std_logic;
  SIGNAL Logical_Operator_out3886_out1            : std_logic;
  SIGNAL Logical_Operator_out3887_out1            : std_logic;
  SIGNAL Logical_Operator_out3888_out1            : std_logic;
  SIGNAL Logical_Operator_out3889_out1            : std_logic;
  SIGNAL Logical_Operator_out3890_out1            : std_logic;
  SIGNAL Logical_Operator_out3891_out1            : std_logic;
  SIGNAL Logical_Operator_out3892_out1            : std_logic;
  SIGNAL Logical_Operator_out3893_out1            : std_logic;
  SIGNAL Logical_Operator_out3894_out1            : std_logic;
  SIGNAL Logical_Operator_out3895_out1            : std_logic;
  SIGNAL Logical_Operator_out3896_out1            : std_logic;
  SIGNAL Logical_Operator_out3897_out1            : std_logic;
  SIGNAL Logical_Operator_out3898_out1            : std_logic;
  SIGNAL Logical_Operator_out3899_out1            : std_logic;
  SIGNAL Logical_Operator_out3900_out1            : std_logic;
  SIGNAL Logical_Operator_out3901_out1            : std_logic;
  SIGNAL Logical_Operator_out3902_out1            : std_logic;
  SIGNAL Logical_Operator_out3903_out1            : std_logic;
  SIGNAL Logical_Operator_out3904_out1            : std_logic;
  SIGNAL Logical_Operator_out3905_out1            : std_logic;
  SIGNAL Logical_Operator_out3906_out1            : std_logic;
  SIGNAL Logical_Operator_out3907_out1            : std_logic;
  SIGNAL Logical_Operator_out3908_out1            : std_logic;
  SIGNAL Logical_Operator_out3909_out1            : std_logic;
  SIGNAL Logical_Operator_out3910_out1            : std_logic;
  SIGNAL Logical_Operator_out3911_out1            : std_logic;
  SIGNAL Logical_Operator_out3912_out1            : std_logic;
  SIGNAL Logical_Operator_out3913_out1            : std_logic;
  SIGNAL Logical_Operator_out3914_out1            : std_logic;
  SIGNAL Logical_Operator_out3915_out1            : std_logic;
  SIGNAL Logical_Operator_out3916_out1            : std_logic;
  SIGNAL Logical_Operator_out3917_out1            : std_logic;
  SIGNAL Logical_Operator_out3918_out1            : std_logic;
  SIGNAL Logical_Operator_out3919_out1            : std_logic;
  SIGNAL Logical_Operator_out3920_out1            : std_logic;
  SIGNAL Logical_Operator_out3921_out1            : std_logic;
  SIGNAL Logical_Operator_out3922_out1            : std_logic;
  SIGNAL Logical_Operator_out3923_out1            : std_logic;
  SIGNAL Logical_Operator_out3924_out1            : std_logic;
  SIGNAL Logical_Operator_out3925_out1            : std_logic;
  SIGNAL Logical_Operator_out3926_out1            : std_logic;
  SIGNAL Logical_Operator_out3927_out1            : std_logic;
  SIGNAL Logical_Operator_out3928_out1            : std_logic;
  SIGNAL Logical_Operator_out3929_out1            : std_logic;
  SIGNAL Logical_Operator_out3930_out1            : std_logic;
  SIGNAL Logical_Operator_out3931_out1            : std_logic;
  SIGNAL Logical_Operator_out3932_out1            : std_logic;
  SIGNAL Logical_Operator_out3933_out1            : std_logic;
  SIGNAL Logical_Operator_out3934_out1            : std_logic;
  SIGNAL Logical_Operator_out3935_out1            : std_logic;
  SIGNAL Logical_Operator_out3936_out1            : std_logic;
  SIGNAL Logical_Operator_out3937_out1            : std_logic;
  SIGNAL Logical_Operator_out3938_out1            : std_logic;
  SIGNAL Logical_Operator_out3939_out1            : std_logic;
  SIGNAL Logical_Operator_out3940_out1            : std_logic;
  SIGNAL Logical_Operator_out3941_out1            : std_logic;
  SIGNAL Logical_Operator_out3942_out1            : std_logic;
  SIGNAL Logical_Operator_out3943_out1            : std_logic;
  SIGNAL Logical_Operator_out3944_out1            : std_logic;
  SIGNAL Logical_Operator_out3945_out1            : std_logic;
  SIGNAL Logical_Operator_out3946_out1            : std_logic;
  SIGNAL Logical_Operator_out3947_out1            : std_logic;
  SIGNAL Logical_Operator_out3948_out1            : std_logic;
  SIGNAL Logical_Operator_out3949_out1            : std_logic;
  SIGNAL Logical_Operator_out3950_out1            : std_logic;
  SIGNAL Logical_Operator_out3951_out1            : std_logic;
  SIGNAL Logical_Operator_out3952_out1            : std_logic;
  SIGNAL Logical_Operator_out3953_out1            : std_logic;
  SIGNAL Logical_Operator_out3954_out1            : std_logic;
  SIGNAL Logical_Operator_out3955_out1            : std_logic;
  SIGNAL Logical_Operator_out3956_out1            : std_logic;
  SIGNAL Logical_Operator_out3957_out1            : std_logic;
  SIGNAL Logical_Operator_out3958_out1            : std_logic;
  SIGNAL Logical_Operator_out3959_out1            : std_logic;
  SIGNAL Logical_Operator_out3960_out1            : std_logic;
  SIGNAL Logical_Operator_out3961_out1            : std_logic;
  SIGNAL Logical_Operator_out3962_out1            : std_logic;
  SIGNAL Logical_Operator_out3963_out1            : std_logic;
  SIGNAL Logical_Operator_out3964_out1            : std_logic;
  SIGNAL Logical_Operator_out3965_out1            : std_logic;
  SIGNAL Logical_Operator_out3966_out1            : std_logic;
  SIGNAL Logical_Operator_out3967_out1            : std_logic;
  SIGNAL Logical_Operator_out3968_out1            : std_logic;
  SIGNAL Logical_Operator_out3969_out1            : std_logic;
  SIGNAL Logical_Operator_out3970_out1            : std_logic;
  SIGNAL Logical_Operator_out3971_out1            : std_logic;
  SIGNAL Logical_Operator_out3972_out1            : std_logic;
  SIGNAL Logical_Operator_out3973_out1            : std_logic;
  SIGNAL Logical_Operator_out3974_out1            : std_logic;
  SIGNAL Logical_Operator_out3975_out1            : std_logic;
  SIGNAL Logical_Operator_out3976_out1            : std_logic;
  SIGNAL Logical_Operator_out3977_out1            : std_logic;
  SIGNAL Logical_Operator_out3978_out1            : std_logic;
  SIGNAL Logical_Operator_out3979_out1            : std_logic;
  SIGNAL Logical_Operator_out3980_out1            : std_logic;
  SIGNAL Logical_Operator_out3981_out1            : std_logic;
  SIGNAL Logical_Operator_out3982_out1            : std_logic;
  SIGNAL Logical_Operator_out3983_out1            : std_logic;
  SIGNAL Logical_Operator_out3984_out1            : std_logic;
  SIGNAL Logical_Operator_out3985_out1            : std_logic;
  SIGNAL Logical_Operator_out3986_out1            : std_logic;
  SIGNAL Logical_Operator_out3987_out1            : std_logic;
  SIGNAL Logical_Operator_out3988_out1            : std_logic;
  SIGNAL Logical_Operator_out3989_out1            : std_logic;
  SIGNAL Logical_Operator_out3990_out1            : std_logic;
  SIGNAL Logical_Operator_out3991_out1            : std_logic;
  SIGNAL Logical_Operator_out3992_out1            : std_logic;
  SIGNAL Logical_Operator_out3993_out1            : std_logic;
  SIGNAL Logical_Operator_out3994_out1            : std_logic;
  SIGNAL Logical_Operator_out3995_out1            : std_logic;
  SIGNAL Logical_Operator_out3996_out1            : std_logic;
  SIGNAL Logical_Operator_out3997_out1            : std_logic;
  SIGNAL Logical_Operator_out3998_out1            : std_logic;
  SIGNAL Logical_Operator_out3999_out1            : std_logic;
  SIGNAL Logical_Operator_out4000_out1            : std_logic;
  SIGNAL Logical_Operator_out4001_out1            : std_logic;
  SIGNAL Logical_Operator_out4002_out1            : std_logic;
  SIGNAL Logical_Operator_out4003_out1            : std_logic;
  SIGNAL Logical_Operator_out4004_out1            : std_logic;
  SIGNAL Logical_Operator_out4005_out1            : std_logic;
  SIGNAL Logical_Operator_out4006_out1            : std_logic;
  SIGNAL Logical_Operator_out4007_out1            : std_logic;
  SIGNAL Logical_Operator_out4008_out1            : std_logic;
  SIGNAL Logical_Operator_out4009_out1            : std_logic;
  SIGNAL Logical_Operator_out4010_out1            : std_logic;
  SIGNAL Logical_Operator_out4011_out1            : std_logic;
  SIGNAL Logical_Operator_out4012_out1            : std_logic;
  SIGNAL Logical_Operator_out4013_out1            : std_logic;
  SIGNAL Logical_Operator_out4014_out1            : std_logic;
  SIGNAL Logical_Operator_out4015_out1            : std_logic;
  SIGNAL Logical_Operator_out4016_out1            : std_logic;
  SIGNAL Logical_Operator_out4017_out1            : std_logic;
  SIGNAL Logical_Operator_out4018_out1            : std_logic;
  SIGNAL Logical_Operator_out4019_out1            : std_logic;
  SIGNAL Logical_Operator_out4020_out1            : std_logic;
  SIGNAL Logical_Operator_out4021_out1            : std_logic;
  SIGNAL Logical_Operator_out4022_out1            : std_logic;
  SIGNAL Logical_Operator_out4023_out1            : std_logic;
  SIGNAL Logical_Operator_out4024_out1            : std_logic;
  SIGNAL Logical_Operator_out4025_out1            : std_logic;
  SIGNAL Logical_Operator_out4026_out1            : std_logic;
  SIGNAL Logical_Operator_out4027_out1            : std_logic;
  SIGNAL Logical_Operator_out4028_out1            : std_logic;
  SIGNAL Logical_Operator_out4029_out1            : std_logic;
  SIGNAL Logical_Operator_out4030_out1            : std_logic;
  SIGNAL Logical_Operator_out4031_out1            : std_logic;
  SIGNAL Logical_Operator_out4032_out1            : std_logic;
  SIGNAL Logical_Operator_out4033_out1            : std_logic;
  SIGNAL Logical_Operator_out4034_out1            : std_logic;
  SIGNAL Logical_Operator_out4035_out1            : std_logic;
  SIGNAL Logical_Operator_out4036_out1            : std_logic;
  SIGNAL Logical_Operator_out4037_out1            : std_logic;
  SIGNAL Logical_Operator_out4038_out1            : std_logic;
  SIGNAL Logical_Operator_out4039_out1            : std_logic;
  SIGNAL Logical_Operator_out4040_out1            : std_logic;
  SIGNAL Logical_Operator_out4041_out1            : std_logic;
  SIGNAL Logical_Operator_out4042_out1            : std_logic;
  SIGNAL Logical_Operator_out4043_out1            : std_logic;
  SIGNAL Logical_Operator_out4044_out1            : std_logic;
  SIGNAL Logical_Operator_out4045_out1            : std_logic;
  SIGNAL Logical_Operator_out4046_out1            : std_logic;
  SIGNAL Logical_Operator_out4047_out1            : std_logic;
  SIGNAL Logical_Operator_out4048_out1            : std_logic;
  SIGNAL Logical_Operator_out4049_out1            : std_logic;
  SIGNAL Logical_Operator_out4050_out1            : std_logic;
  SIGNAL Logical_Operator_out4051_out1            : std_logic;
  SIGNAL Logical_Operator_out4052_out1            : std_logic;
  SIGNAL Logical_Operator_out4053_out1            : std_logic;
  SIGNAL Logical_Operator_out4054_out1            : std_logic;
  SIGNAL Logical_Operator_out4055_out1            : std_logic;
  SIGNAL Logical_Operator_out4056_out1            : std_logic;
  SIGNAL Logical_Operator_out4057_out1            : std_logic;
  SIGNAL Logical_Operator_out4058_out1            : std_logic;
  SIGNAL Logical_Operator_out4059_out1            : std_logic;
  SIGNAL Logical_Operator_out4060_out1            : std_logic;
  SIGNAL Logical_Operator_out4061_out1            : std_logic;
  SIGNAL Logical_Operator_out4062_out1            : std_logic;
  SIGNAL Logical_Operator_out4063_out1            : std_logic;
  SIGNAL Logical_Operator_out4064_out1            : std_logic;
  SIGNAL Logical_Operator_out4065_out1            : std_logic;
  SIGNAL Logical_Operator_out4066_out1            : std_logic;
  SIGNAL Logical_Operator_out4067_out1            : std_logic;
  SIGNAL Logical_Operator_out4068_out1            : std_logic;
  SIGNAL Logical_Operator_out4069_out1            : std_logic;
  SIGNAL Logical_Operator_out4070_out1            : std_logic;
  SIGNAL Logical_Operator_out4071_out1            : std_logic;
  SIGNAL Logical_Operator_out4072_out1            : std_logic;
  SIGNAL Logical_Operator_out4073_out1            : std_logic;
  SIGNAL Logical_Operator_out4074_out1            : std_logic;
  SIGNAL Logical_Operator_out4075_out1            : std_logic;
  SIGNAL Logical_Operator_out4076_out1            : std_logic;
  SIGNAL Logical_Operator_out4077_out1            : std_logic;
  SIGNAL Logical_Operator_out4078_out1            : std_logic;
  SIGNAL Logical_Operator_out4079_out1            : std_logic;
  SIGNAL Logical_Operator_out4080_out1            : std_logic;
  SIGNAL Logical_Operator_out4081_out1            : std_logic;
  SIGNAL Logical_Operator_out4082_out1            : std_logic;
  SIGNAL Logical_Operator_out4083_out1            : std_logic;
  SIGNAL Logical_Operator_out4084_out1            : std_logic;
  SIGNAL Logical_Operator_out4085_out1            : std_logic;
  SIGNAL Logical_Operator_out4086_out1            : std_logic;
  SIGNAL Logical_Operator_out4087_out1            : std_logic;
  SIGNAL Logical_Operator_out4088_out1            : std_logic;
  SIGNAL Logical_Operator_out4089_out1            : std_logic;
  SIGNAL Logical_Operator_out4090_out1            : std_logic;
  SIGNAL Logical_Operator_out4091_out1            : std_logic;
  SIGNAL Logical_Operator_out4092_out1            : std_logic;
  SIGNAL Logical_Operator_out4093_out1            : std_logic;
  SIGNAL Logical_Operator_out4094_out1            : std_logic;
  SIGNAL Logical_Operator_out4095_out1            : std_logic;
  SIGNAL Logical_Operator_out4096_out1            : std_logic;
  SIGNAL Logical_Operator_out4097_out1            : std_logic;
  SIGNAL Logical_Operator_out4098_out1            : std_logic;
  SIGNAL Logical_Operator_out4099_out1            : std_logic;
  SIGNAL Logical_Operator_out4100_out1            : std_logic;
  SIGNAL Logical_Operator_out4101_out1            : std_logic;
  SIGNAL Logical_Operator_out4102_out1            : std_logic;
  SIGNAL Logical_Operator_out4103_out1            : std_logic;
  SIGNAL Logical_Operator_out4104_out1            : std_logic;
  SIGNAL Logical_Operator_out4105_out1            : std_logic;
  SIGNAL Logical_Operator_out4106_out1            : std_logic;
  SIGNAL Logical_Operator_out4107_out1            : std_logic;
  SIGNAL Logical_Operator_out4108_out1            : std_logic;
  SIGNAL Logical_Operator_out4109_out1            : std_logic;
  SIGNAL Logical_Operator_out4110_out1            : std_logic;
  SIGNAL Logical_Operator_out4111_out1            : std_logic;
  SIGNAL Logical_Operator_out4112_out1            : std_logic;
  SIGNAL Logical_Operator_out4113_out1            : std_logic;
  SIGNAL Logical_Operator_out4114_out1            : std_logic;
  SIGNAL Logical_Operator_out4115_out1            : std_logic;
  SIGNAL Logical_Operator_out4116_out1            : std_logic;
  SIGNAL Logical_Operator_out4117_out1            : std_logic;
  SIGNAL Logical_Operator_out4118_out1            : std_logic;
  SIGNAL Logical_Operator_out4119_out1            : std_logic;
  SIGNAL Logical_Operator_out4120_out1            : std_logic;
  SIGNAL Logical_Operator_out4121_out1            : std_logic;
  SIGNAL Logical_Operator_out4122_out1            : std_logic;
  SIGNAL Logical_Operator_out4123_out1            : std_logic;
  SIGNAL Logical_Operator_out4124_out1            : std_logic;
  SIGNAL Logical_Operator_out4125_out1            : std_logic;
  SIGNAL Logical_Operator_out4126_out1            : std_logic;
  SIGNAL Logical_Operator_out4127_out1            : std_logic;
  SIGNAL Logical_Operator_out4128_out1            : std_logic;
  SIGNAL Logical_Operator_out4129_out1            : std_logic;
  SIGNAL Logical_Operator_out4130_out1            : std_logic;
  SIGNAL Logical_Operator_out4131_out1            : std_logic;
  SIGNAL Logical_Operator_out4132_out1            : std_logic;
  SIGNAL Logical_Operator_out4133_out1            : std_logic;
  SIGNAL Logical_Operator_out4134_out1            : std_logic;
  SIGNAL Logical_Operator_out4135_out1            : std_logic;
  SIGNAL Logical_Operator_out4136_out1            : std_logic;
  SIGNAL Logical_Operator_out4137_out1            : std_logic;
  SIGNAL Logical_Operator_out4138_out1            : std_logic;
  SIGNAL Logical_Operator_out4139_out1            : std_logic;
  SIGNAL Logical_Operator_out4140_out1            : std_logic;
  SIGNAL Logical_Operator_out4141_out1            : std_logic;
  SIGNAL Logical_Operator_out4142_out1            : std_logic;
  SIGNAL Logical_Operator_out4143_out1            : std_logic;
  SIGNAL Logical_Operator_out4144_out1            : std_logic;
  SIGNAL Logical_Operator_out4145_out1            : std_logic;
  SIGNAL Logical_Operator_out4146_out1            : std_logic;
  SIGNAL Logical_Operator_out4147_out1            : std_logic;
  SIGNAL Logical_Operator_out4148_out1            : std_logic;
  SIGNAL Logical_Operator_out4149_out1            : std_logic;
  SIGNAL Logical_Operator_out4150_out1            : std_logic;
  SIGNAL Logical_Operator_out4151_out1            : std_logic;
  SIGNAL Logical_Operator_out4152_out1            : std_logic;
  SIGNAL Logical_Operator_out4153_out1            : std_logic;
  SIGNAL Logical_Operator_out4154_out1            : std_logic;
  SIGNAL Logical_Operator_out4155_out1            : std_logic;
  SIGNAL Logical_Operator_out4156_out1            : std_logic;
  SIGNAL Logical_Operator_out4157_out1            : std_logic;
  SIGNAL Logical_Operator_out4158_out1            : std_logic;
  SIGNAL Logical_Operator_out4159_out1            : std_logic;
  SIGNAL Logical_Operator_out4160_out1            : std_logic;
  SIGNAL Logical_Operator_out4161_out1            : std_logic;
  SIGNAL Logical_Operator_out4162_out1            : std_logic;
  SIGNAL Logical_Operator_out4163_out1            : std_logic;
  SIGNAL Logical_Operator_out4164_out1            : std_logic;
  SIGNAL Logical_Operator_out4165_out1            : std_logic;
  SIGNAL Logical_Operator_out4166_out1            : std_logic;
  SIGNAL Logical_Operator_out4167_out1            : std_logic;
  SIGNAL Logical_Operator_out4168_out1            : std_logic;
  SIGNAL Logical_Operator_out4169_out1            : std_logic;
  SIGNAL Logical_Operator_out4170_out1            : std_logic;
  SIGNAL Logical_Operator_out4171_out1            : std_logic;
  SIGNAL Logical_Operator_out4172_out1            : std_logic;
  SIGNAL Logical_Operator_out4173_out1            : std_logic;
  SIGNAL Logical_Operator_out4174_out1            : std_logic;
  SIGNAL Logical_Operator_out4175_out1            : std_logic;
  SIGNAL Logical_Operator_out4176_out1            : std_logic;
  SIGNAL Logical_Operator_out4177_out1            : std_logic;
  SIGNAL Logical_Operator_out4178_out1            : std_logic;
  SIGNAL Logical_Operator_out4179_out1            : std_logic;
  SIGNAL Logical_Operator_out4180_out1            : std_logic;
  SIGNAL Logical_Operator_out4181_out1            : std_logic;
  SIGNAL Logical_Operator_out4182_out1            : std_logic;
  SIGNAL Logical_Operator_out4183_out1            : std_logic;
  SIGNAL Logical_Operator_out4184_out1            : std_logic;
  SIGNAL Logical_Operator_out4185_out1            : std_logic;
  SIGNAL Logical_Operator_out4186_out1            : std_logic;
  SIGNAL Logical_Operator_out4187_out1            : std_logic;
  SIGNAL Logical_Operator_out4188_out1            : std_logic;
  SIGNAL Logical_Operator_out4189_out1            : std_logic;
  SIGNAL Logical_Operator_out4190_out1            : std_logic;
  SIGNAL Logical_Operator_out4191_out1            : std_logic;
  SIGNAL Logical_Operator_out4192_out1            : std_logic;
  SIGNAL Logical_Operator_out4193_out1            : std_logic;
  SIGNAL Logical_Operator_out4194_out1            : std_logic;
  SIGNAL Logical_Operator_out4195_out1            : std_logic;
  SIGNAL Logical_Operator_out4196_out1            : std_logic;
  SIGNAL Logical_Operator_out4197_out1            : std_logic;
  SIGNAL Logical_Operator_out4198_out1            : std_logic;
  SIGNAL Logical_Operator_out4199_out1            : std_logic;
  SIGNAL Logical_Operator_out4200_out1            : std_logic;
  SIGNAL Logical_Operator_out4201_out1            : std_logic;
  SIGNAL Logical_Operator_out4202_out1            : std_logic;
  SIGNAL Logical_Operator_out4203_out1            : std_logic;
  SIGNAL Logical_Operator_out4204_out1            : std_logic;
  SIGNAL Logical_Operator_out4205_out1            : std_logic;
  SIGNAL Logical_Operator_out4206_out1            : std_logic;
  SIGNAL Logical_Operator_out4207_out1            : std_logic;
  SIGNAL Logical_Operator_out4208_out1            : std_logic;
  SIGNAL Logical_Operator_out4209_out1            : std_logic;
  SIGNAL Logical_Operator_out4210_out1            : std_logic;
  SIGNAL Logical_Operator_out4211_out1            : std_logic;
  SIGNAL Logical_Operator_out4212_out1            : std_logic;
  SIGNAL Logical_Operator_out4213_out1            : std_logic;
  SIGNAL Logical_Operator_out4214_out1            : std_logic;
  SIGNAL Logical_Operator_out4215_out1            : std_logic;
  SIGNAL Logical_Operator_out4216_out1            : std_logic;
  SIGNAL Logical_Operator_out4217_out1            : std_logic;
  SIGNAL Logical_Operator_out4218_out1            : std_logic;
  SIGNAL Logical_Operator_out4219_out1            : std_logic;
  SIGNAL Logical_Operator_out4220_out1            : std_logic;
  SIGNAL Logical_Operator_out4221_out1            : std_logic;
  SIGNAL Logical_Operator_out4222_out1            : std_logic;
  SIGNAL Logical_Operator_out4223_out1            : std_logic;
  SIGNAL Logical_Operator_out4224_out1            : std_logic;
  SIGNAL Logical_Operator_out4225_out1            : std_logic;
  SIGNAL Logical_Operator_out4226_out1            : std_logic;
  SIGNAL Logical_Operator_out4227_out1            : std_logic;
  SIGNAL Logical_Operator_out4228_out1            : std_logic;
  SIGNAL Logical_Operator_out4229_out1            : std_logic;
  SIGNAL Logical_Operator_out4230_out1            : std_logic;
  SIGNAL Logical_Operator_out4231_out1            : std_logic;
  SIGNAL Logical_Operator_out4232_out1            : std_logic;
  SIGNAL Logical_Operator_out4233_out1            : std_logic;
  SIGNAL Logical_Operator_out4234_out1            : std_logic;
  SIGNAL Logical_Operator_out4235_out1            : std_logic;
  SIGNAL Logical_Operator_out4236_out1            : std_logic;
  SIGNAL Logical_Operator_out4237_out1            : std_logic;
  SIGNAL Logical_Operator_out4238_out1            : std_logic;
  SIGNAL Logical_Operator_out4239_out1            : std_logic;
  SIGNAL Logical_Operator_out4240_out1            : std_logic;
  SIGNAL Logical_Operator_out4241_out1            : std_logic;
  SIGNAL Logical_Operator_out4242_out1            : std_logic;
  SIGNAL Logical_Operator_out4243_out1            : std_logic;
  SIGNAL Logical_Operator_out4244_out1            : std_logic;
  SIGNAL Logical_Operator_out4245_out1            : std_logic;
  SIGNAL Logical_Operator_out4246_out1            : std_logic;
  SIGNAL Logical_Operator_out4247_out1            : std_logic;
  SIGNAL Logical_Operator_out4248_out1            : std_logic;
  SIGNAL Logical_Operator_out4249_out1            : std_logic;
  SIGNAL Logical_Operator_out4250_out1            : std_logic;
  SIGNAL Logical_Operator_out4251_out1            : std_logic;
  SIGNAL Logical_Operator_out4252_out1            : std_logic;
  SIGNAL Logical_Operator_out4253_out1            : std_logic;
  SIGNAL Logical_Operator_out4254_out1            : std_logic;
  SIGNAL Logical_Operator_out4255_out1            : std_logic;
  SIGNAL Logical_Operator_out4256_out1            : std_logic;
  SIGNAL Logical_Operator_out4257_out1            : std_logic;
  SIGNAL Logical_Operator_out4258_out1            : std_logic;
  SIGNAL Logical_Operator_out4259_out1            : std_logic;
  SIGNAL Logical_Operator_out4260_out1            : std_logic;
  SIGNAL Logical_Operator_out4261_out1            : std_logic;
  SIGNAL Logical_Operator_out4262_out1            : std_logic;
  SIGNAL Logical_Operator_out4263_out1            : std_logic;
  SIGNAL Logical_Operator_out4264_out1            : std_logic;
  SIGNAL Logical_Operator_out4265_out1            : std_logic;
  SIGNAL Logical_Operator_out4266_out1            : std_logic;
  SIGNAL Logical_Operator_out4267_out1            : std_logic;
  SIGNAL Logical_Operator_out4268_out1            : std_logic;
  SIGNAL Logical_Operator_out4269_out1            : std_logic;
  SIGNAL Logical_Operator_out4270_out1            : std_logic;
  SIGNAL Logical_Operator_out4271_out1            : std_logic;
  SIGNAL Logical_Operator_out4272_out1            : std_logic;
  SIGNAL Logical_Operator_out4273_out1            : std_logic;
  SIGNAL Logical_Operator_out4274_out1            : std_logic;
  SIGNAL Logical_Operator_out4275_out1            : std_logic;
  SIGNAL Logical_Operator_out4276_out1            : std_logic;
  SIGNAL Logical_Operator_out4277_out1            : std_logic;
  SIGNAL Logical_Operator_out4278_out1            : std_logic;
  SIGNAL Logical_Operator_out4279_out1            : std_logic;
  SIGNAL Logical_Operator_out4280_out1            : std_logic;
  SIGNAL Logical_Operator_out4281_out1            : std_logic;
  SIGNAL Logical_Operator_out4282_out1            : std_logic;
  SIGNAL Logical_Operator_out4283_out1            : std_logic;
  SIGNAL Logical_Operator_out4284_out1            : std_logic;
  SIGNAL Logical_Operator_out4285_out1            : std_logic;
  SIGNAL Logical_Operator_out4286_out1            : std_logic;
  SIGNAL Logical_Operator_out4287_out1            : std_logic;
  SIGNAL Logical_Operator_out4288_out1            : std_logic;
  SIGNAL Logical_Operator_out4289_out1            : std_logic;
  SIGNAL Logical_Operator_out4290_out1            : std_logic;
  SIGNAL Logical_Operator_out4291_out1            : std_logic;
  SIGNAL Logical_Operator_out4292_out1            : std_logic;
  SIGNAL Logical_Operator_out4293_out1            : std_logic;
  SIGNAL Logical_Operator_out4294_out1            : std_logic;
  SIGNAL Logical_Operator_out4295_out1            : std_logic;
  SIGNAL Logical_Operator_out4296_out1            : std_logic;
  SIGNAL Logical_Operator_out4297_out1            : std_logic;
  SIGNAL Logical_Operator_out4298_out1            : std_logic;
  SIGNAL Logical_Operator_out4299_out1            : std_logic;
  SIGNAL Logical_Operator_out4300_out1            : std_logic;
  SIGNAL Logical_Operator_out4301_out1            : std_logic;
  SIGNAL Logical_Operator_out4302_out1            : std_logic;
  SIGNAL Logical_Operator_out4303_out1            : std_logic;
  SIGNAL Logical_Operator_out4304_out1            : std_logic;
  SIGNAL Logical_Operator_out4305_out1            : std_logic;
  SIGNAL Logical_Operator_out4306_out1            : std_logic;
  SIGNAL Logical_Operator_out4307_out1            : std_logic;
  SIGNAL Logical_Operator_out4308_out1            : std_logic;
  SIGNAL Logical_Operator_out4309_out1            : std_logic;
  SIGNAL Logical_Operator_out4310_out1            : std_logic;
  SIGNAL Logical_Operator_out4311_out1            : std_logic;
  SIGNAL Logical_Operator_out4312_out1            : std_logic;
  SIGNAL Logical_Operator_out4313_out1            : std_logic;
  SIGNAL Logical_Operator_out4314_out1            : std_logic;
  SIGNAL Logical_Operator_out4315_out1            : std_logic;
  SIGNAL Logical_Operator_out4316_out1            : std_logic;
  SIGNAL Logical_Operator_out4317_out1            : std_logic;
  SIGNAL Logical_Operator_out4318_out1            : std_logic;
  SIGNAL Logical_Operator_out4319_out1            : std_logic;
  SIGNAL Logical_Operator_out4320_out1            : std_logic;
  SIGNAL Logical_Operator_out4321_out1            : std_logic;
  SIGNAL Logical_Operator_out4322_out1            : std_logic;
  SIGNAL Logical_Operator_out4323_out1            : std_logic;
  SIGNAL Logical_Operator_out4324_out1            : std_logic;
  SIGNAL Logical_Operator_out4325_out1            : std_logic;
  SIGNAL Logical_Operator_out4326_out1            : std_logic;
  SIGNAL Logical_Operator_out4327_out1            : std_logic;
  SIGNAL Logical_Operator_out4328_out1            : std_logic;
  SIGNAL Logical_Operator_out4329_out1            : std_logic;
  SIGNAL Logical_Operator_out4330_out1            : std_logic;
  SIGNAL Logical_Operator_out4331_out1            : std_logic;
  SIGNAL Logical_Operator_out4332_out1            : std_logic;
  SIGNAL Logical_Operator_out4333_out1            : std_logic;
  SIGNAL Logical_Operator_out4334_out1            : std_logic;
  SIGNAL Logical_Operator_out4335_out1            : std_logic;
  SIGNAL Logical_Operator_out4336_out1            : std_logic;
  SIGNAL Logical_Operator_out4337_out1            : std_logic;
  SIGNAL Logical_Operator_out4338_out1            : std_logic;
  SIGNAL Logical_Operator_out4339_out1            : std_logic;
  SIGNAL Logical_Operator_out4340_out1            : std_logic;
  SIGNAL Logical_Operator_out4341_out1            : std_logic;
  SIGNAL Logical_Operator_out4342_out1            : std_logic;
  SIGNAL Logical_Operator_out4343_out1            : std_logic;
  SIGNAL Logical_Operator_out4344_out1            : std_logic;
  SIGNAL Logical_Operator_out4345_out1            : std_logic;
  SIGNAL Logical_Operator_out4346_out1            : std_logic;
  SIGNAL Logical_Operator_out4347_out1            : std_logic;
  SIGNAL Logical_Operator_out4348_out1            : std_logic;
  SIGNAL Logical_Operator_out4349_out1            : std_logic;
  SIGNAL Logical_Operator_out4350_out1            : std_logic;
  SIGNAL Logical_Operator_out4351_out1            : std_logic;
  SIGNAL Logical_Operator_out4352_out1            : std_logic;
  SIGNAL Logical_Operator_out4353_out1            : std_logic;
  SIGNAL Logical_Operator_out4354_out1            : std_logic;
  SIGNAL Logical_Operator_out4355_out1            : std_logic;
  SIGNAL Logical_Operator_out4356_out1            : std_logic;
  SIGNAL Logical_Operator_out4357_out1            : std_logic;
  SIGNAL Logical_Operator_out4358_out1            : std_logic;
  SIGNAL Logical_Operator_out4359_out1            : std_logic;
  SIGNAL Logical_Operator_out4360_out1            : std_logic;
  SIGNAL Logical_Operator_out4361_out1            : std_logic;
  SIGNAL Logical_Operator_out4362_out1            : std_logic;
  SIGNAL Logical_Operator_out4363_out1            : std_logic;
  SIGNAL Logical_Operator_out4364_out1            : std_logic;
  SIGNAL Logical_Operator_out4365_out1            : std_logic;
  SIGNAL Logical_Operator_out4366_out1            : std_logic;
  SIGNAL Logical_Operator_out4367_out1            : std_logic;
  SIGNAL Logical_Operator_out4368_out1            : std_logic;
  SIGNAL Logical_Operator_out4369_out1            : std_logic;
  SIGNAL Logical_Operator_out4370_out1            : std_logic;
  SIGNAL Logical_Operator_out4371_out1            : std_logic;
  SIGNAL Logical_Operator_out4372_out1            : std_logic;
  SIGNAL Logical_Operator_out4373_out1            : std_logic;
  SIGNAL Logical_Operator_out4374_out1            : std_logic;
  SIGNAL Logical_Operator_out4375_out1            : std_logic;
  SIGNAL Logical_Operator_out4376_out1            : std_logic;
  SIGNAL Logical_Operator_out4377_out1            : std_logic;
  SIGNAL Logical_Operator_out4378_out1            : std_logic;
  SIGNAL Logical_Operator_out4379_out1            : std_logic;
  SIGNAL Logical_Operator_out4380_out1            : std_logic;
  SIGNAL Logical_Operator_out4381_out1            : std_logic;
  SIGNAL Logical_Operator_out4382_out1            : std_logic;
  SIGNAL Logical_Operator_out4383_out1            : std_logic;
  SIGNAL Logical_Operator_out4384_out1            : std_logic;
  SIGNAL Logical_Operator_out4385_out1            : std_logic;
  SIGNAL Logical_Operator_out4386_out1            : std_logic;
  SIGNAL Logical_Operator_out4387_out1            : std_logic;
  SIGNAL Logical_Operator_out4388_out1            : std_logic;
  SIGNAL Logical_Operator_out4389_out1            : std_logic;
  SIGNAL Logical_Operator_out4390_out1            : std_logic;
  SIGNAL Logical_Operator_out4391_out1            : std_logic;
  SIGNAL Logical_Operator_out4392_out1            : std_logic;
  SIGNAL Logical_Operator_out4393_out1            : std_logic;
  SIGNAL Logical_Operator_out4394_out1            : std_logic;
  SIGNAL Logical_Operator_out4395_out1            : std_logic;
  SIGNAL Logical_Operator_out4396_out1            : std_logic;
  SIGNAL Logical_Operator_out4397_out1            : std_logic;
  SIGNAL Logical_Operator_out4398_out1            : std_logic;
  SIGNAL Logical_Operator_out4399_out1            : std_logic;
  SIGNAL Logical_Operator_out4400_out1            : std_logic;
  SIGNAL Logical_Operator_out4401_out1            : std_logic;
  SIGNAL Logical_Operator_out4402_out1            : std_logic;
  SIGNAL Logical_Operator_out4403_out1            : std_logic;
  SIGNAL Logical_Operator_out4404_out1            : std_logic;
  SIGNAL Logical_Operator_out4405_out1            : std_logic;
  SIGNAL Logical_Operator_out4406_out1            : std_logic;
  SIGNAL Logical_Operator_out4407_out1            : std_logic;
  SIGNAL Logical_Operator_out4408_out1            : std_logic;
  SIGNAL Logical_Operator_out4409_out1            : std_logic;
  SIGNAL Logical_Operator_out4410_out1            : std_logic;
  SIGNAL Logical_Operator_out4411_out1            : std_logic;
  SIGNAL Logical_Operator_out4412_out1            : std_logic;
  SIGNAL Logical_Operator_out4413_out1            : std_logic;
  SIGNAL Logical_Operator_out4414_out1            : std_logic;
  SIGNAL Logical_Operator_out4415_out1            : std_logic;
  SIGNAL Logical_Operator_out4416_out1            : std_logic;
  SIGNAL Logical_Operator_out4417_out1            : std_logic;
  SIGNAL Logical_Operator_out4418_out1            : std_logic;
  SIGNAL Logical_Operator_out4419_out1            : std_logic;
  SIGNAL Logical_Operator_out4420_out1            : std_logic;
  SIGNAL Logical_Operator_out4421_out1            : std_logic;
  SIGNAL Logical_Operator_out4422_out1            : std_logic;
  SIGNAL Logical_Operator_out4423_out1            : std_logic;
  SIGNAL Logical_Operator_out4424_out1            : std_logic;
  SIGNAL Logical_Operator_out4425_out1            : std_logic;
  SIGNAL Logical_Operator_out4426_out1            : std_logic;
  SIGNAL Logical_Operator_out4427_out1            : std_logic;
  SIGNAL Logical_Operator_out4428_out1            : std_logic;
  SIGNAL Logical_Operator_out4429_out1            : std_logic;
  SIGNAL Logical_Operator_out4430_out1            : std_logic;
  SIGNAL Logical_Operator_out4431_out1            : std_logic;
  SIGNAL Logical_Operator_out4432_out1            : std_logic;
  SIGNAL Logical_Operator_out4433_out1            : std_logic;
  SIGNAL Logical_Operator_out4434_out1            : std_logic;
  SIGNAL Logical_Operator_out4435_out1            : std_logic;
  SIGNAL Logical_Operator_out4436_out1            : std_logic;
  SIGNAL Logical_Operator_out4437_out1            : std_logic;
  SIGNAL Logical_Operator_out4438_out1            : std_logic;
  SIGNAL Logical_Operator_out4439_out1            : std_logic;
  SIGNAL Logical_Operator_out4440_out1            : std_logic;
  SIGNAL Logical_Operator_out4441_out1            : std_logic;
  SIGNAL Logical_Operator_out4442_out1            : std_logic;
  SIGNAL Logical_Operator_out4443_out1            : std_logic;
  SIGNAL Logical_Operator_out4444_out1            : std_logic;
  SIGNAL Logical_Operator_out4445_out1            : std_logic;
  SIGNAL Logical_Operator_out4446_out1            : std_logic;
  SIGNAL Logical_Operator_out4447_out1            : std_logic;
  SIGNAL Logical_Operator_out4448_out1            : std_logic;
  SIGNAL Logical_Operator_out4449_out1            : std_logic;
  SIGNAL Logical_Operator_out4450_out1            : std_logic;
  SIGNAL Logical_Operator_out4451_out1            : std_logic;
  SIGNAL Logical_Operator_out4452_out1            : std_logic;
  SIGNAL Logical_Operator_out4453_out1            : std_logic;
  SIGNAL Logical_Operator_out4454_out1            : std_logic;
  SIGNAL Logical_Operator_out4455_out1            : std_logic;
  SIGNAL Logical_Operator_out4456_out1            : std_logic;
  SIGNAL Logical_Operator_out4457_out1            : std_logic;
  SIGNAL Logical_Operator_out4458_out1            : std_logic;
  SIGNAL Logical_Operator_out4459_out1            : std_logic;
  SIGNAL Logical_Operator_out4460_out1            : std_logic;
  SIGNAL Logical_Operator_out4461_out1            : std_logic;
  SIGNAL Logical_Operator_out4462_out1            : std_logic;
  SIGNAL Logical_Operator_out4463_out1            : std_logic;
  SIGNAL Logical_Operator_out4464_out1            : std_logic;
  SIGNAL Logical_Operator_out4465_out1            : std_logic;
  SIGNAL Logical_Operator_out4466_out1            : std_logic;
  SIGNAL Logical_Operator_out4467_out1            : std_logic;
  SIGNAL Logical_Operator_out4468_out1            : std_logic;
  SIGNAL Logical_Operator_out4469_out1            : std_logic;
  SIGNAL Logical_Operator_out4470_out1            : std_logic;
  SIGNAL Logical_Operator_out4471_out1            : std_logic;
  SIGNAL Logical_Operator_out4472_out1            : std_logic;
  SIGNAL Logical_Operator_out4473_out1            : std_logic;
  SIGNAL Logical_Operator_out4474_out1            : std_logic;
  SIGNAL Logical_Operator_out4475_out1            : std_logic;
  SIGNAL Logical_Operator_out4476_out1            : std_logic;
  SIGNAL Logical_Operator_out4477_out1            : std_logic;
  SIGNAL Logical_Operator_out4478_out1            : std_logic;
  SIGNAL Logical_Operator_out4479_out1            : std_logic;
  SIGNAL Logical_Operator_out4480_out1            : std_logic;
  SIGNAL Logical_Operator_out4481_out1            : std_logic;
  SIGNAL Logical_Operator_out4482_out1            : std_logic;
  SIGNAL Logical_Operator_out4483_out1            : std_logic;
  SIGNAL Logical_Operator_out4484_out1            : std_logic;
  SIGNAL Logical_Operator_out4485_out1            : std_logic;
  SIGNAL Logical_Operator_out4486_out1            : std_logic;
  SIGNAL Logical_Operator_out4487_out1            : std_logic;
  SIGNAL Logical_Operator_out4488_out1            : std_logic;
  SIGNAL Logical_Operator_out4489_out1            : std_logic;
  SIGNAL Logical_Operator_out4490_out1            : std_logic;
  SIGNAL Logical_Operator_out4491_out1            : std_logic;
  SIGNAL Logical_Operator_out4492_out1            : std_logic;
  SIGNAL Logical_Operator_out4493_out1            : std_logic;
  SIGNAL Logical_Operator_out4494_out1            : std_logic;
  SIGNAL Logical_Operator_out4495_out1            : std_logic;
  SIGNAL Logical_Operator_out4496_out1            : std_logic;
  SIGNAL Logical_Operator_out4497_out1            : std_logic;
  SIGNAL Logical_Operator_out4498_out1            : std_logic;
  SIGNAL Logical_Operator_out4499_out1            : std_logic;
  SIGNAL Logical_Operator_out4500_out1            : std_logic;
  SIGNAL Logical_Operator_out4501_out1            : std_logic;
  SIGNAL Logical_Operator_out4502_out1            : std_logic;
  SIGNAL Logical_Operator_out4503_out1            : std_logic;
  SIGNAL Logical_Operator_out4504_out1            : std_logic;
  SIGNAL Logical_Operator_out4505_out1            : std_logic;
  SIGNAL Logical_Operator_out4506_out1            : std_logic;
  SIGNAL Logical_Operator_out4507_out1            : std_logic;
  SIGNAL Logical_Operator_out4508_out1            : std_logic;
  SIGNAL Logical_Operator_out4509_out1            : std_logic;
  SIGNAL Logical_Operator_out4510_out1            : std_logic;
  SIGNAL Logical_Operator_out4511_out1            : std_logic;
  SIGNAL Logical_Operator_out4512_out1            : std_logic;
  SIGNAL Logical_Operator_out4513_out1            : std_logic;
  SIGNAL Logical_Operator_out4514_out1            : std_logic;
  SIGNAL Logical_Operator_out4515_out1            : std_logic;
  SIGNAL Logical_Operator_out4516_out1            : std_logic;
  SIGNAL Logical_Operator_out4517_out1            : std_logic;
  SIGNAL Logical_Operator_out4518_out1            : std_logic;
  SIGNAL Logical_Operator_out4519_out1            : std_logic;
  SIGNAL Logical_Operator_out4520_out1            : std_logic;
  SIGNAL Logical_Operator_out4521_out1            : std_logic;
  SIGNAL Logical_Operator_out4522_out1            : std_logic;
  SIGNAL Logical_Operator_out4523_out1            : std_logic;
  SIGNAL Logical_Operator_out4524_out1            : std_logic;
  SIGNAL Logical_Operator_out4525_out1            : std_logic;
  SIGNAL Logical_Operator_out4526_out1            : std_logic;
  SIGNAL Logical_Operator_out4527_out1            : std_logic;
  SIGNAL Logical_Operator_out4528_out1            : std_logic;
  SIGNAL Logical_Operator_out4529_out1            : std_logic;
  SIGNAL Logical_Operator_out4530_out1            : std_logic;
  SIGNAL Logical_Operator_out4531_out1            : std_logic;
  SIGNAL Logical_Operator_out4532_out1            : std_logic;
  SIGNAL Logical_Operator_out4533_out1            : std_logic;
  SIGNAL Logical_Operator_out4534_out1            : std_logic;
  SIGNAL Logical_Operator_out4535_out1            : std_logic;
  SIGNAL Logical_Operator_out4536_out1            : std_logic;
  SIGNAL Logical_Operator_out4537_out1            : std_logic;
  SIGNAL Logical_Operator_out4538_out1            : std_logic;
  SIGNAL Logical_Operator_out4539_out1            : std_logic;
  SIGNAL Logical_Operator_out4540_out1            : std_logic;
  SIGNAL Logical_Operator_out4541_out1            : std_logic;
  SIGNAL Logical_Operator_out4542_out1            : std_logic;
  SIGNAL Logical_Operator_out4543_out1            : std_logic;
  SIGNAL Logical_Operator_out4544_out1            : std_logic;
  SIGNAL Logical_Operator_out4545_out1            : std_logic;
  SIGNAL Logical_Operator_out4546_out1            : std_logic;
  SIGNAL Logical_Operator_out4547_out1            : std_logic;
  SIGNAL Logical_Operator_out4548_out1            : std_logic;
  SIGNAL Logical_Operator_out4549_out1            : std_logic;
  SIGNAL Logical_Operator_out4550_out1            : std_logic;
  SIGNAL Logical_Operator_out4551_out1            : std_logic;
  SIGNAL Logical_Operator_out4552_out1            : std_logic;
  SIGNAL Logical_Operator_out4553_out1            : std_logic;
  SIGNAL Logical_Operator_out4554_out1            : std_logic;
  SIGNAL Logical_Operator_out4555_out1            : std_logic;
  SIGNAL Logical_Operator_out4556_out1            : std_logic;
  SIGNAL Logical_Operator_out4557_out1            : std_logic;
  SIGNAL Logical_Operator_out4558_out1            : std_logic;
  SIGNAL Logical_Operator_out4559_out1            : std_logic;
  SIGNAL Logical_Operator_out4560_out1            : std_logic;
  SIGNAL Logical_Operator_out4561_out1            : std_logic;
  SIGNAL Logical_Operator_out4562_out1            : std_logic;
  SIGNAL Logical_Operator_out4563_out1            : std_logic;
  SIGNAL Logical_Operator_out4564_out1            : std_logic;
  SIGNAL Logical_Operator_out4565_out1            : std_logic;
  SIGNAL Logical_Operator_out4566_out1            : std_logic;
  SIGNAL Logical_Operator_out4567_out1            : std_logic;
  SIGNAL Logical_Operator_out4568_out1            : std_logic;
  SIGNAL Logical_Operator_out4569_out1            : std_logic;
  SIGNAL Logical_Operator_out4570_out1            : std_logic;
  SIGNAL Logical_Operator_out4571_out1            : std_logic;
  SIGNAL Logical_Operator_out4572_out1            : std_logic;
  SIGNAL Logical_Operator_out4573_out1            : std_logic;
  SIGNAL Logical_Operator_out4574_out1            : std_logic;
  SIGNAL Logical_Operator_out4575_out1            : std_logic;
  SIGNAL Logical_Operator_out4576_out1            : std_logic;
  SIGNAL Logical_Operator_out4577_out1            : std_logic;
  SIGNAL Logical_Operator_out4578_out1            : std_logic;
  SIGNAL Logical_Operator_out4579_out1            : std_logic;
  SIGNAL Logical_Operator_out4580_out1            : std_logic;
  SIGNAL Logical_Operator_out4581_out1            : std_logic;
  SIGNAL Logical_Operator_out4582_out1            : std_logic;
  SIGNAL Logical_Operator_out4583_out1            : std_logic;
  SIGNAL Logical_Operator_out4584_out1            : std_logic;
  SIGNAL Logical_Operator_out4585_out1            : std_logic;
  SIGNAL Logical_Operator_out4586_out1            : std_logic;
  SIGNAL Logical_Operator_out4587_out1            : std_logic;
  SIGNAL Logical_Operator_out4588_out1            : std_logic;
  SIGNAL Logical_Operator_out4589_out1            : std_logic;
  SIGNAL Logical_Operator_out4590_out1            : std_logic;
  SIGNAL Logical_Operator_out4591_out1            : std_logic;
  SIGNAL Logical_Operator_out4592_out1            : std_logic;
  SIGNAL Logical_Operator_out4593_out1            : std_logic;
  SIGNAL Logical_Operator_out4594_out1            : std_logic;
  SIGNAL Logical_Operator_out4595_out1            : std_logic;
  SIGNAL Logical_Operator_out4596_out1            : std_logic;
  SIGNAL Logical_Operator_out4597_out1            : std_logic;
  SIGNAL Logical_Operator_out4598_out1            : std_logic;
  SIGNAL Logical_Operator_out4599_out1            : std_logic;
  SIGNAL Logical_Operator_out4600_out1            : std_logic;
  SIGNAL Logical_Operator_out4601_out1            : std_logic;
  SIGNAL Logical_Operator_out4602_out1            : std_logic;
  SIGNAL Logical_Operator_out4603_out1            : std_logic;
  SIGNAL Logical_Operator_out4604_out1            : std_logic;
  SIGNAL Logical_Operator_out4605_out1            : std_logic;
  SIGNAL Logical_Operator_out4606_out1            : std_logic;
  SIGNAL Logical_Operator_out4607_out1            : std_logic;
  SIGNAL Logical_Operator_out4608_out1            : std_logic;
  SIGNAL Logical_Operator_out4609_out1            : std_logic;
  SIGNAL Logical_Operator_out4610_out1            : std_logic;
  SIGNAL Logical_Operator_out4611_out1            : std_logic;
  SIGNAL Logical_Operator_out4612_out1            : std_logic;
  SIGNAL Logical_Operator_out4613_out1            : std_logic;
  SIGNAL Logical_Operator_out4614_out1            : std_logic;
  SIGNAL Logical_Operator_out4615_out1            : std_logic;
  SIGNAL Logical_Operator_out4616_out1            : std_logic;
  SIGNAL Logical_Operator_out4617_out1            : std_logic;
  SIGNAL Logical_Operator_out4618_out1            : std_logic;
  SIGNAL Logical_Operator_out4619_out1            : std_logic;
  SIGNAL Logical_Operator_out4620_out1            : std_logic;
  SIGNAL Logical_Operator_out4621_out1            : std_logic;
  SIGNAL Logical_Operator_out4622_out1            : std_logic;
  SIGNAL Logical_Operator_out4623_out1            : std_logic;
  SIGNAL Logical_Operator_out4624_out1            : std_logic;
  SIGNAL Logical_Operator_out4625_out1            : std_logic;
  SIGNAL Logical_Operator_out4626_out1            : std_logic;
  SIGNAL Logical_Operator_out4627_out1            : std_logic;
  SIGNAL Logical_Operator_out4628_out1            : std_logic;
  SIGNAL Logical_Operator_out4629_out1            : std_logic;
  SIGNAL Logical_Operator_out4630_out1            : std_logic;
  SIGNAL Logical_Operator_out4631_out1            : std_logic;
  SIGNAL Logical_Operator_out4632_out1            : std_logic;
  SIGNAL Logical_Operator_out4633_out1            : std_logic;
  SIGNAL Logical_Operator_out4634_out1            : std_logic;
  SIGNAL Logical_Operator_out4635_out1            : std_logic;
  SIGNAL Logical_Operator_out4636_out1            : std_logic;
  SIGNAL Logical_Operator_out4637_out1            : std_logic;
  SIGNAL Logical_Operator_out4638_out1            : std_logic;
  SIGNAL Logical_Operator_out4639_out1            : std_logic;
  SIGNAL Logical_Operator_out4640_out1            : std_logic;
  SIGNAL Logical_Operator_out4641_out1            : std_logic;
  SIGNAL Logical_Operator_out4642_out1            : std_logic;
  SIGNAL Logical_Operator_out4643_out1            : std_logic;
  SIGNAL Logical_Operator_out4644_out1            : std_logic;
  SIGNAL Logical_Operator_out4645_out1            : std_logic;
  SIGNAL Logical_Operator_out4646_out1            : std_logic;
  SIGNAL Logical_Operator_out4647_out1            : std_logic;
  SIGNAL Logical_Operator_out4648_out1            : std_logic;
  SIGNAL Logical_Operator_out4649_out1            : std_logic;
  SIGNAL Logical_Operator_out4650_out1            : std_logic;
  SIGNAL Logical_Operator_out4651_out1            : std_logic;
  SIGNAL Logical_Operator_out4652_out1            : std_logic;
  SIGNAL Logical_Operator_out4653_out1            : std_logic;
  SIGNAL Logical_Operator_out4654_out1            : std_logic;
  SIGNAL Logical_Operator_out4655_out1            : std_logic;
  SIGNAL Logical_Operator_out4656_out1            : std_logic;
  SIGNAL Logical_Operator_out4657_out1            : std_logic;
  SIGNAL Logical_Operator_out4658_out1            : std_logic;
  SIGNAL Logical_Operator_out4659_out1            : std_logic;
  SIGNAL Logical_Operator_out4660_out1            : std_logic;
  SIGNAL Logical_Operator_out4661_out1            : std_logic;
  SIGNAL Logical_Operator_out4662_out1            : std_logic;
  SIGNAL Logical_Operator_out4663_out1            : std_logic;
  SIGNAL Logical_Operator_out4664_out1            : std_logic;
  SIGNAL Logical_Operator_out4665_out1            : std_logic;
  SIGNAL Logical_Operator_out4666_out1            : std_logic;
  SIGNAL Logical_Operator_out4667_out1            : std_logic;
  SIGNAL Logical_Operator_out4668_out1            : std_logic;
  SIGNAL Logical_Operator_out4669_out1            : std_logic;
  SIGNAL Logical_Operator_out4670_out1            : std_logic;
  SIGNAL Logical_Operator_out4671_out1            : std_logic;
  SIGNAL Logical_Operator_out4672_out1            : std_logic;
  SIGNAL Logical_Operator_out4673_out1            : std_logic;
  SIGNAL Logical_Operator_out4674_out1            : std_logic;
  SIGNAL Logical_Operator_out4675_out1            : std_logic;
  SIGNAL Logical_Operator_out4676_out1            : std_logic;
  SIGNAL Logical_Operator_out4677_out1            : std_logic;
  SIGNAL Logical_Operator_out4678_out1            : std_logic;
  SIGNAL Logical_Operator_out4679_out1            : std_logic;
  SIGNAL Logical_Operator_out4680_out1            : std_logic;
  SIGNAL Logical_Operator_out4681_out1            : std_logic;
  SIGNAL Logical_Operator_out4682_out1            : std_logic;
  SIGNAL Logical_Operator_out4683_out1            : std_logic;
  SIGNAL Logical_Operator_out4684_out1            : std_logic;
  SIGNAL Logical_Operator_out4685_out1            : std_logic;
  SIGNAL Logical_Operator_out4686_out1            : std_logic;
  SIGNAL Logical_Operator_out4687_out1            : std_logic;
  SIGNAL Logical_Operator_out4688_out1            : std_logic;
  SIGNAL Logical_Operator_out4689_out1            : std_logic;
  SIGNAL Logical_Operator_out4690_out1            : std_logic;
  SIGNAL Logical_Operator_out4691_out1            : std_logic;
  SIGNAL Logical_Operator_out4692_out1            : std_logic;
  SIGNAL Logical_Operator_out4693_out1            : std_logic;
  SIGNAL Logical_Operator_out4694_out1            : std_logic;
  SIGNAL Logical_Operator_out4695_out1            : std_logic;
  SIGNAL Logical_Operator_out4696_out1            : std_logic;
  SIGNAL Logical_Operator_out4697_out1            : std_logic;
  SIGNAL Logical_Operator_out4698_out1            : std_logic;
  SIGNAL Logical_Operator_out4699_out1            : std_logic;
  SIGNAL Logical_Operator_out4700_out1            : std_logic;
  SIGNAL Logical_Operator_out4701_out1            : std_logic;
  SIGNAL Logical_Operator_out4702_out1            : std_logic;
  SIGNAL Logical_Operator_out4703_out1            : std_logic;
  SIGNAL Logical_Operator_out4704_out1            : std_logic;
  SIGNAL Logical_Operator_out4705_out1            : std_logic;
  SIGNAL Logical_Operator_out4706_out1            : std_logic;
  SIGNAL Logical_Operator_out4707_out1            : std_logic;
  SIGNAL Logical_Operator_out4708_out1            : std_logic;
  SIGNAL Logical_Operator_out4709_out1            : std_logic;
  SIGNAL Logical_Operator_out4710_out1            : std_logic;
  SIGNAL Logical_Operator_out4711_out1            : std_logic;
  SIGNAL Logical_Operator_out4712_out1            : std_logic;
  SIGNAL Logical_Operator_out4713_out1            : std_logic;
  SIGNAL Logical_Operator_out4714_out1            : std_logic;
  SIGNAL Logical_Operator_out4715_out1            : std_logic;
  SIGNAL Logical_Operator_out4716_out1            : std_logic;
  SIGNAL Logical_Operator_out4717_out1            : std_logic;
  SIGNAL Logical_Operator_out4718_out1            : std_logic;
  SIGNAL Logical_Operator_out4719_out1            : std_logic;
  SIGNAL Logical_Operator_out4720_out1            : std_logic;
  SIGNAL Logical_Operator_out4721_out1            : std_logic;
  SIGNAL Logical_Operator_out4722_out1            : std_logic;
  SIGNAL Logical_Operator_out4723_out1            : std_logic;
  SIGNAL Logical_Operator_out4724_out1            : std_logic;
  SIGNAL Logical_Operator_out4725_out1            : std_logic;
  SIGNAL Logical_Operator_out4726_out1            : std_logic;
  SIGNAL Logical_Operator_out4727_out1            : std_logic;
  SIGNAL Logical_Operator_out4728_out1            : std_logic;
  SIGNAL Logical_Operator_out4729_out1            : std_logic;
  SIGNAL Logical_Operator_out4730_out1            : std_logic;
  SIGNAL Logical_Operator_out4731_out1            : std_logic;
  SIGNAL Logical_Operator_out4732_out1            : std_logic;
  SIGNAL Logical_Operator_out4733_out1            : std_logic;
  SIGNAL Logical_Operator_out4734_out1            : std_logic;
  SIGNAL Logical_Operator_out4735_out1            : std_logic;
  SIGNAL Logical_Operator_out4736_out1            : std_logic;
  SIGNAL Logical_Operator_out4737_out1            : std_logic;
  SIGNAL Logical_Operator_out4738_out1            : std_logic;
  SIGNAL Logical_Operator_out4739_out1            : std_logic;
  SIGNAL Logical_Operator_out4740_out1            : std_logic;
  SIGNAL Logical_Operator_out4741_out1            : std_logic;
  SIGNAL Logical_Operator_out4742_out1            : std_logic;
  SIGNAL Logical_Operator_out4743_out1            : std_logic;
  SIGNAL Logical_Operator_out4744_out1            : std_logic;
  SIGNAL Logical_Operator_out4745_out1            : std_logic;
  SIGNAL Logical_Operator_out4746_out1            : std_logic;
  SIGNAL Logical_Operator_out4747_out1            : std_logic;
  SIGNAL Logical_Operator_out4748_out1            : std_logic;
  SIGNAL Logical_Operator_out4749_out1            : std_logic;
  SIGNAL Logical_Operator_out4750_out1            : std_logic;
  SIGNAL Logical_Operator_out4751_out1            : std_logic;
  SIGNAL Logical_Operator_out4752_out1            : std_logic;
  SIGNAL Logical_Operator_out4753_out1            : std_logic;
  SIGNAL Logical_Operator_out4754_out1            : std_logic;
  SIGNAL Logical_Operator_out4755_out1            : std_logic;
  SIGNAL Logical_Operator_out4756_out1            : std_logic;
  SIGNAL Logical_Operator_out4757_out1            : std_logic;
  SIGNAL Logical_Operator_out4758_out1            : std_logic;
  SIGNAL Logical_Operator_out4759_out1            : std_logic;
  SIGNAL Logical_Operator_out4760_out1            : std_logic;
  SIGNAL Logical_Operator_out4761_out1            : std_logic;
  SIGNAL Logical_Operator_out4762_out1            : std_logic;
  SIGNAL Logical_Operator_out4763_out1            : std_logic;
  SIGNAL Logical_Operator_out4764_out1            : std_logic;
  SIGNAL Logical_Operator_out4765_out1            : std_logic;
  SIGNAL Logical_Operator_out4766_out1            : std_logic;
  SIGNAL Logical_Operator_out4767_out1            : std_logic;
  SIGNAL Logical_Operator_out4768_out1            : std_logic;
  SIGNAL Logical_Operator_out4769_out1            : std_logic;
  SIGNAL Logical_Operator_out4770_out1            : std_logic;
  SIGNAL Logical_Operator_out4771_out1            : std_logic;
  SIGNAL Logical_Operator_out4772_out1            : std_logic;
  SIGNAL Logical_Operator_out4773_out1            : std_logic;
  SIGNAL Logical_Operator_out4774_out1            : std_logic;
  SIGNAL Logical_Operator_out4775_out1            : std_logic;
  SIGNAL Logical_Operator_out4776_out1            : std_logic;
  SIGNAL Logical_Operator_out4777_out1            : std_logic;
  SIGNAL Logical_Operator_out4778_out1            : std_logic;
  SIGNAL Logical_Operator_out4779_out1            : std_logic;
  SIGNAL Logical_Operator_out4780_out1            : std_logic;
  SIGNAL Logical_Operator_out4781_out1            : std_logic;
  SIGNAL Logical_Operator_out4782_out1            : std_logic;
  SIGNAL Logical_Operator_out4783_out1            : std_logic;
  SIGNAL Logical_Operator_out4784_out1            : std_logic;
  SIGNAL Logical_Operator_out4785_out1            : std_logic;
  SIGNAL Logical_Operator_out4786_out1            : std_logic;
  SIGNAL Logical_Operator_out4787_out1            : std_logic;
  SIGNAL Logical_Operator_out4788_out1            : std_logic;
  SIGNAL Logical_Operator_out4789_out1            : std_logic;
  SIGNAL Logical_Operator_out4790_out1            : std_logic;
  SIGNAL Logical_Operator_out4791_out1            : std_logic;
  SIGNAL Logical_Operator_out4792_out1            : std_logic;
  SIGNAL Logical_Operator_out4793_out1            : std_logic;
  SIGNAL Logical_Operator_out4794_out1            : std_logic;
  SIGNAL Logical_Operator_out4795_out1            : std_logic;
  SIGNAL Logical_Operator_out4796_out1            : std_logic;
  SIGNAL Logical_Operator_out4797_out1            : std_logic;
  SIGNAL Logical_Operator_out4798_out1            : std_logic;
  SIGNAL Logical_Operator_out4799_out1            : std_logic;
  SIGNAL Logical_Operator_out4800_out1            : std_logic;
  SIGNAL Logical_Operator_out4801_out1            : std_logic;
  SIGNAL Logical_Operator_out4802_out1            : std_logic;
  SIGNAL Logical_Operator_out4803_out1            : std_logic;
  SIGNAL Logical_Operator_out4804_out1            : std_logic;
  SIGNAL Logical_Operator_out4805_out1            : std_logic;
  SIGNAL Logical_Operator_out4806_out1            : std_logic;
  SIGNAL Logical_Operator_out4807_out1            : std_logic;
  SIGNAL Logical_Operator_out4808_out1            : std_logic;
  SIGNAL Logical_Operator_out4809_out1            : std_logic;
  SIGNAL Logical_Operator_out4810_out1            : std_logic;
  SIGNAL Logical_Operator_out4811_out1            : std_logic;
  SIGNAL Logical_Operator_out4812_out1            : std_logic;
  SIGNAL Logical_Operator_out4813_out1            : std_logic;
  SIGNAL Logical_Operator_out4814_out1            : std_logic;
  SIGNAL Logical_Operator_out4815_out1            : std_logic;
  SIGNAL Logical_Operator_out4816_out1            : std_logic;
  SIGNAL Logical_Operator_out4817_out1            : std_logic;
  SIGNAL Logical_Operator_out4818_out1            : std_logic;
  SIGNAL Logical_Operator_out4819_out1            : std_logic;
  SIGNAL Logical_Operator_out4820_out1            : std_logic;
  SIGNAL Logical_Operator_out4821_out1            : std_logic;
  SIGNAL Logical_Operator_out4822_out1            : std_logic;
  SIGNAL Logical_Operator_out4823_out1            : std_logic;
  SIGNAL Logical_Operator_out4824_out1            : std_logic;
  SIGNAL Logical_Operator_out4825_out1            : std_logic;
  SIGNAL Logical_Operator_out4826_out1            : std_logic;
  SIGNAL Logical_Operator_out4827_out1            : std_logic;
  SIGNAL Logical_Operator_out4828_out1            : std_logic;
  SIGNAL Logical_Operator_out4829_out1            : std_logic;
  SIGNAL Logical_Operator_out4830_out1            : std_logic;
  SIGNAL Logical_Operator_out4831_out1            : std_logic;
  SIGNAL Logical_Operator_out4832_out1            : std_logic;
  SIGNAL Logical_Operator_out4833_out1            : std_logic;
  SIGNAL Logical_Operator_out4834_out1            : std_logic;
  SIGNAL Logical_Operator_out4835_out1            : std_logic;
  SIGNAL Logical_Operator_out4836_out1            : std_logic;
  SIGNAL Logical_Operator_out4837_out1            : std_logic;
  SIGNAL Logical_Operator_out4838_out1            : std_logic;
  SIGNAL Logical_Operator_out4839_out1            : std_logic;
  SIGNAL Logical_Operator_out4840_out1            : std_logic;
  SIGNAL Logical_Operator_out4841_out1            : std_logic;
  SIGNAL Logical_Operator_out4842_out1            : std_logic;
  SIGNAL Logical_Operator_out4843_out1            : std_logic;
  SIGNAL Logical_Operator_out4844_out1            : std_logic;
  SIGNAL Logical_Operator_out4845_out1            : std_logic;
  SIGNAL Logical_Operator_out4846_out1            : std_logic;
  SIGNAL Logical_Operator_out4847_out1            : std_logic;
  SIGNAL Logical_Operator_out4848_out1            : std_logic;
  SIGNAL Logical_Operator_out4849_out1            : std_logic;
  SIGNAL Logical_Operator_out4850_out1            : std_logic;
  SIGNAL Logical_Operator_out4851_out1            : std_logic;
  SIGNAL Logical_Operator_out4852_out1            : std_logic;
  SIGNAL Logical_Operator_out4853_out1            : std_logic;
  SIGNAL Logical_Operator_out4854_out1            : std_logic;
  SIGNAL Logical_Operator_out4855_out1            : std_logic;
  SIGNAL Logical_Operator_out4856_out1            : std_logic;
  SIGNAL Logical_Operator_out4857_out1            : std_logic;
  SIGNAL Logical_Operator_out4858_out1            : std_logic;
  SIGNAL Logical_Operator_out4859_out1            : std_logic;
  SIGNAL Logical_Operator_out4860_out1            : std_logic;
  SIGNAL Logical_Operator_out4861_out1            : std_logic;
  SIGNAL Logical_Operator_out4862_out1            : std_logic;
  SIGNAL Logical_Operator_out4863_out1            : std_logic;
  SIGNAL Logical_Operator_out4864_out1            : std_logic;
  SIGNAL Logical_Operator_out4865_out1            : std_logic;
  SIGNAL Logical_Operator_out4866_out1            : std_logic;
  SIGNAL Logical_Operator_out4867_out1            : std_logic;
  SIGNAL Logical_Operator_out4868_out1            : std_logic;
  SIGNAL Logical_Operator_out4869_out1            : std_logic;
  SIGNAL Logical_Operator_out4870_out1            : std_logic;
  SIGNAL Logical_Operator_out4871_out1            : std_logic;
  SIGNAL Logical_Operator_out4872_out1            : std_logic;
  SIGNAL Logical_Operator_out4873_out1            : std_logic;
  SIGNAL Logical_Operator_out4874_out1            : std_logic;
  SIGNAL Logical_Operator_out4875_out1            : std_logic;
  SIGNAL Logical_Operator_out4876_out1            : std_logic;
  SIGNAL Logical_Operator_out4877_out1            : std_logic;
  SIGNAL Logical_Operator_out4878_out1            : std_logic;
  SIGNAL Logical_Operator_out4879_out1            : std_logic;
  SIGNAL Logical_Operator_out4880_out1            : std_logic;
  SIGNAL Logical_Operator_out4881_out1            : std_logic;
  SIGNAL Logical_Operator_out4882_out1            : std_logic;
  SIGNAL Logical_Operator_out4883_out1            : std_logic;
  SIGNAL Logical_Operator_out4884_out1            : std_logic;
  SIGNAL Logical_Operator_out4885_out1            : std_logic;
  SIGNAL Logical_Operator_out4886_out1            : std_logic;
  SIGNAL Logical_Operator_out4887_out1            : std_logic;
  SIGNAL Logical_Operator_out4888_out1            : std_logic;
  SIGNAL Logical_Operator_out4889_out1            : std_logic;
  SIGNAL Logical_Operator_out4890_out1            : std_logic;
  SIGNAL Logical_Operator_out4891_out1            : std_logic;
  SIGNAL Logical_Operator_out4892_out1            : std_logic;
  SIGNAL Logical_Operator_out4893_out1            : std_logic;
  SIGNAL Logical_Operator_out4894_out1            : std_logic;
  SIGNAL Logical_Operator_out4895_out1            : std_logic;
  SIGNAL Logical_Operator_out4896_out1            : std_logic;
  SIGNAL Logical_Operator_out4897_out1            : std_logic;
  SIGNAL Logical_Operator_out4898_out1            : std_logic;
  SIGNAL Logical_Operator_out4899_out1            : std_logic;
  SIGNAL Logical_Operator_out4900_out1            : std_logic;
  SIGNAL Logical_Operator_out4901_out1            : std_logic;
  SIGNAL Logical_Operator_out4902_out1            : std_logic;
  SIGNAL Logical_Operator_out4903_out1            : std_logic;
  SIGNAL Logical_Operator_out4904_out1            : std_logic;
  SIGNAL Logical_Operator_out4905_out1            : std_logic;
  SIGNAL Logical_Operator_out4906_out1            : std_logic;
  SIGNAL Logical_Operator_out4907_out1            : std_logic;
  SIGNAL Logical_Operator_out4908_out1            : std_logic;
  SIGNAL Logical_Operator_out4909_out1            : std_logic;
  SIGNAL Logical_Operator_out4910_out1            : std_logic;
  SIGNAL Logical_Operator_out4911_out1            : std_logic;
  SIGNAL Logical_Operator_out4912_out1            : std_logic;
  SIGNAL Logical_Operator_out4913_out1            : std_logic;
  SIGNAL Logical_Operator_out4914_out1            : std_logic;
  SIGNAL Logical_Operator_out4915_out1            : std_logic;
  SIGNAL Logical_Operator_out4916_out1            : std_logic;
  SIGNAL Logical_Operator_out4917_out1            : std_logic;
  SIGNAL Logical_Operator_out4918_out1            : std_logic;
  SIGNAL Logical_Operator_out4919_out1            : std_logic;
  SIGNAL Logical_Operator_out4920_out1            : std_logic;
  SIGNAL Logical_Operator_out4921_out1            : std_logic;
  SIGNAL Logical_Operator_out4922_out1            : std_logic;
  SIGNAL Logical_Operator_out4923_out1            : std_logic;
  SIGNAL Logical_Operator_out4924_out1            : std_logic;
  SIGNAL Logical_Operator_out4925_out1            : std_logic;
  SIGNAL Logical_Operator_out4926_out1            : std_logic;
  SIGNAL Logical_Operator_out4927_out1            : std_logic;
  SIGNAL Logical_Operator_out4928_out1            : std_logic;
  SIGNAL Logical_Operator_out4929_out1            : std_logic;
  SIGNAL Logical_Operator_out4930_out1            : std_logic;
  SIGNAL Logical_Operator_out4931_out1            : std_logic;
  SIGNAL Logical_Operator_out4932_out1            : std_logic;
  SIGNAL Logical_Operator_out4933_out1            : std_logic;
  SIGNAL Logical_Operator_out4934_out1            : std_logic;
  SIGNAL Logical_Operator_out4935_out1            : std_logic;
  SIGNAL Logical_Operator_out4936_out1            : std_logic;
  SIGNAL Logical_Operator_out4937_out1            : std_logic;
  SIGNAL Logical_Operator_out4938_out1            : std_logic;
  SIGNAL Logical_Operator_out4939_out1            : std_logic;
  SIGNAL Logical_Operator_out4940_out1            : std_logic;
  SIGNAL Logical_Operator_out4941_out1            : std_logic;
  SIGNAL Logical_Operator_out4942_out1            : std_logic;
  SIGNAL Logical_Operator_out4943_out1            : std_logic;
  SIGNAL Logical_Operator_out4944_out1            : std_logic;
  SIGNAL Logical_Operator_out4945_out1            : std_logic;
  SIGNAL Logical_Operator_out4946_out1            : std_logic;
  SIGNAL Logical_Operator_out4947_out1            : std_logic;
  SIGNAL Logical_Operator_out4948_out1            : std_logic;
  SIGNAL Logical_Operator_out4949_out1            : std_logic;
  SIGNAL Logical_Operator_out4950_out1            : std_logic;
  SIGNAL Logical_Operator_out4951_out1            : std_logic;
  SIGNAL Logical_Operator_out4952_out1            : std_logic;
  SIGNAL Logical_Operator_out4953_out1            : std_logic;
  SIGNAL Logical_Operator_out4954_out1            : std_logic;
  SIGNAL Logical_Operator_out4955_out1            : std_logic;
  SIGNAL Logical_Operator_out4956_out1            : std_logic;
  SIGNAL Logical_Operator_out4957_out1            : std_logic;
  SIGNAL Logical_Operator_out4958_out1            : std_logic;
  SIGNAL Logical_Operator_out4959_out1            : std_logic;
  SIGNAL Logical_Operator_out4960_out1            : std_logic;
  SIGNAL Logical_Operator_out4961_out1            : std_logic;
  SIGNAL Logical_Operator_out4962_out1            : std_logic;
  SIGNAL Logical_Operator_out4963_out1            : std_logic;
  SIGNAL Logical_Operator_out4964_out1            : std_logic;
  SIGNAL Logical_Operator_out4965_out1            : std_logic;
  SIGNAL Logical_Operator_out4966_out1            : std_logic;
  SIGNAL Logical_Operator_out4967_out1            : std_logic;
  SIGNAL Logical_Operator_out4968_out1            : std_logic;
  SIGNAL Logical_Operator_out4969_out1            : std_logic;
  SIGNAL Logical_Operator_out4970_out1            : std_logic;
  SIGNAL Logical_Operator_out4971_out1            : std_logic;
  SIGNAL Logical_Operator_out4972_out1            : std_logic;
  SIGNAL Logical_Operator_out4973_out1            : std_logic;
  SIGNAL Logical_Operator_out4974_out1            : std_logic;
  SIGNAL Logical_Operator_out4975_out1            : std_logic;
  SIGNAL Logical_Operator_out4976_out1            : std_logic;
  SIGNAL Logical_Operator_out4977_out1            : std_logic;
  SIGNAL Logical_Operator_out4978_out1            : std_logic;
  SIGNAL Logical_Operator_out4979_out1            : std_logic;
  SIGNAL Logical_Operator_out4980_out1            : std_logic;
  SIGNAL Logical_Operator_out4981_out1            : std_logic;
  SIGNAL Logical_Operator_out4982_out1            : std_logic;
  SIGNAL Logical_Operator_out4983_out1            : std_logic;
  SIGNAL Logical_Operator_out4984_out1            : std_logic;
  SIGNAL Logical_Operator_out4985_out1            : std_logic;
  SIGNAL Logical_Operator_out4986_out1            : std_logic;
  SIGNAL Logical_Operator_out4987_out1            : std_logic;
  SIGNAL Logical_Operator_out4988_out1            : std_logic;
  SIGNAL Logical_Operator_out4989_out1            : std_logic;
  SIGNAL Logical_Operator_out4990_out1            : std_logic;
  SIGNAL Logical_Operator_out4991_out1            : std_logic;
  SIGNAL Logical_Operator_out4992_out1            : std_logic;
  SIGNAL Logical_Operator_out4993_out1            : std_logic;
  SIGNAL Logical_Operator_out4994_out1            : std_logic;
  SIGNAL Logical_Operator_out4995_out1            : std_logic;
  SIGNAL Logical_Operator_out4996_out1            : std_logic;
  SIGNAL Logical_Operator_out4997_out1            : std_logic;
  SIGNAL Logical_Operator_out4998_out1            : std_logic;
  SIGNAL Logical_Operator_out4999_out1            : std_logic;
  SIGNAL Logical_Operator_out5000_out1            : std_logic;
  SIGNAL Logical_Operator_out5001_out1            : std_logic;
  SIGNAL Logical_Operator_out5002_out1            : std_logic;
  SIGNAL Logical_Operator_out5003_out1            : std_logic;
  SIGNAL Logical_Operator_out5004_out1            : std_logic;
  SIGNAL Logical_Operator_out5005_out1            : std_logic;
  SIGNAL Logical_Operator_out5006_out1            : std_logic;
  SIGNAL Logical_Operator_out5007_out1            : std_logic;
  SIGNAL Logical_Operator_out5008_out1            : std_logic;
  SIGNAL Logical_Operator_out5009_out1            : std_logic;
  SIGNAL Logical_Operator_out5010_out1            : std_logic;
  SIGNAL Logical_Operator_out5011_out1            : std_logic;
  SIGNAL Logical_Operator_out5012_out1            : std_logic;
  SIGNAL Logical_Operator_out5013_out1            : std_logic;
  SIGNAL Logical_Operator_out5014_out1            : std_logic;
  SIGNAL Logical_Operator_out5015_out1            : std_logic;
  SIGNAL Logical_Operator_out5016_out1            : std_logic;
  SIGNAL Logical_Operator_out5017_out1            : std_logic;
  SIGNAL Logical_Operator_out5018_out1            : std_logic;
  SIGNAL Logical_Operator_out5019_out1            : std_logic;
  SIGNAL Logical_Operator_out5020_out1            : std_logic;
  SIGNAL Logical_Operator_out5021_out1            : std_logic;
  SIGNAL Logical_Operator_out5022_out1            : std_logic;
  SIGNAL Logical_Operator_out5023_out1            : std_logic;
  SIGNAL Logical_Operator_out5024_out1            : std_logic;
  SIGNAL Logical_Operator_out5025_out1            : std_logic;
  SIGNAL Logical_Operator_out5026_out1            : std_logic;
  SIGNAL Logical_Operator_out5027_out1            : std_logic;
  SIGNAL Logical_Operator_out5028_out1            : std_logic;
  SIGNAL Logical_Operator_out5029_out1            : std_logic;
  SIGNAL Logical_Operator_out5030_out1            : std_logic;
  SIGNAL Logical_Operator_out5031_out1            : std_logic;
  SIGNAL Logical_Operator_out5032_out1            : std_logic;
  SIGNAL Logical_Operator_out5033_out1            : std_logic;
  SIGNAL Logical_Operator_out5034_out1            : std_logic;
  SIGNAL Logical_Operator_out5035_out1            : std_logic;
  SIGNAL Logical_Operator_out5036_out1            : std_logic;
  SIGNAL Logical_Operator_out5037_out1            : std_logic;
  SIGNAL Logical_Operator_out5038_out1            : std_logic;
  SIGNAL Logical_Operator_out5039_out1            : std_logic;
  SIGNAL Logical_Operator_out5040_out1            : std_logic;
  SIGNAL Logical_Operator_out5041_out1            : std_logic;
  SIGNAL Logical_Operator_out5042_out1            : std_logic;
  SIGNAL Logical_Operator_out5043_out1            : std_logic;
  SIGNAL Logical_Operator_out5044_out1            : std_logic;
  SIGNAL Logical_Operator_out5045_out1            : std_logic;
  SIGNAL Logical_Operator_out5046_out1            : std_logic;
  SIGNAL Logical_Operator_out5047_out1            : std_logic;
  SIGNAL Logical_Operator_out5048_out1            : std_logic;
  SIGNAL Logical_Operator_out5049_out1            : std_logic;
  SIGNAL Logical_Operator_out5050_out1            : std_logic;
  SIGNAL Logical_Operator_out5051_out1            : std_logic;
  SIGNAL Logical_Operator_out5052_out1            : std_logic;
  SIGNAL Logical_Operator_out5053_out1            : std_logic;
  SIGNAL Logical_Operator_out5054_out1            : std_logic;
  SIGNAL Logical_Operator_out5055_out1            : std_logic;
  SIGNAL Logical_Operator_out5056_out1            : std_logic;
  SIGNAL Logical_Operator_out5057_out1            : std_logic;
  SIGNAL Logical_Operator_out5058_out1            : std_logic;
  SIGNAL Logical_Operator_out5059_out1            : std_logic;
  SIGNAL Logical_Operator_out5060_out1            : std_logic;
  SIGNAL Logical_Operator_out5061_out1            : std_logic;
  SIGNAL Logical_Operator_out5062_out1            : std_logic;
  SIGNAL Logical_Operator_out5063_out1            : std_logic;
  SIGNAL Logical_Operator_out5064_out1            : std_logic;
  SIGNAL Logical_Operator_out5065_out1            : std_logic;
  SIGNAL Logical_Operator_out5066_out1            : std_logic;
  SIGNAL Logical_Operator_out5067_out1            : std_logic;
  SIGNAL Logical_Operator_out5068_out1            : std_logic;
  SIGNAL Logical_Operator_out5069_out1            : std_logic;
  SIGNAL Logical_Operator_out5070_out1            : std_logic;
  SIGNAL Logical_Operator_out5071_out1            : std_logic;
  SIGNAL Logical_Operator_out5072_out1            : std_logic;
  SIGNAL Logical_Operator_out5073_out1            : std_logic;
  SIGNAL Logical_Operator_out5074_out1            : std_logic;
  SIGNAL Logical_Operator_out5075_out1            : std_logic;
  SIGNAL Logical_Operator_out5076_out1            : std_logic;
  SIGNAL Logical_Operator_out5077_out1            : std_logic;
  SIGNAL Logical_Operator_out5078_out1            : std_logic;
  SIGNAL Logical_Operator_out5079_out1            : std_logic;
  SIGNAL Logical_Operator_out5080_out1            : std_logic;
  SIGNAL Logical_Operator_out5081_out1            : std_logic;
  SIGNAL Logical_Operator_out5082_out1            : std_logic;
  SIGNAL Logical_Operator_out5083_out1            : std_logic;
  SIGNAL Logical_Operator_out5084_out1            : std_logic;
  SIGNAL Logical_Operator_out5085_out1            : std_logic;
  SIGNAL Logical_Operator_out5086_out1            : std_logic;
  SIGNAL Logical_Operator_out5087_out1            : std_logic;
  SIGNAL Logical_Operator_out5088_out1            : std_logic;
  SIGNAL Logical_Operator_out5089_out1            : std_logic;
  SIGNAL Logical_Operator_out5090_out1            : std_logic;
  SIGNAL Logical_Operator_out5091_out1            : std_logic;
  SIGNAL Logical_Operator_out5092_out1            : std_logic;
  SIGNAL Logical_Operator_out5093_out1            : std_logic;
  SIGNAL Logical_Operator_out5094_out1            : std_logic;
  SIGNAL Logical_Operator_out5095_out1            : std_logic;
  SIGNAL Logical_Operator_out5096_out1            : std_logic;
  SIGNAL Logical_Operator_out5097_out1            : std_logic;
  SIGNAL Logical_Operator_out5098_out1            : std_logic;
  SIGNAL Logical_Operator_out5099_out1            : std_logic;
  SIGNAL Logical_Operator_out5100_out1            : std_logic;
  SIGNAL Logical_Operator_out5101_out1            : std_logic;
  SIGNAL Logical_Operator_out5102_out1            : std_logic;
  SIGNAL Logical_Operator_out5103_out1            : std_logic;
  SIGNAL Logical_Operator_out5104_out1            : std_logic;
  SIGNAL Logical_Operator_out5105_out1            : std_logic;
  SIGNAL Logical_Operator_out5106_out1            : std_logic;
  SIGNAL Logical_Operator_out5107_out1            : std_logic;
  SIGNAL Logical_Operator_out5108_out1            : std_logic;
  SIGNAL Logical_Operator_out5109_out1            : std_logic;
  SIGNAL Logical_Operator_out5110_out1            : std_logic;
  SIGNAL Logical_Operator_out5111_out1            : std_logic;
  SIGNAL Logical_Operator_out5112_out1            : std_logic;
  SIGNAL Logical_Operator_out5113_out1            : std_logic;
  SIGNAL Logical_Operator_out5114_out1            : std_logic;
  SIGNAL Logical_Operator_out5115_out1            : std_logic;
  SIGNAL Logical_Operator_out5116_out1            : std_logic;
  SIGNAL Logical_Operator_out5117_out1            : std_logic;
  SIGNAL Logical_Operator_out5118_out1            : std_logic;
  SIGNAL Logical_Operator_out5119_out1            : std_logic;
  SIGNAL Logical_Operator_out5120_out1            : std_logic;
  SIGNAL Logical_Operator_out5121_out1            : std_logic;
  SIGNAL Logical_Operator_out5122_out1            : std_logic;
  SIGNAL Logical_Operator_out5123_out1            : std_logic;
  SIGNAL Logical_Operator_out5124_out1            : std_logic;
  SIGNAL Logical_Operator_out5125_out1            : std_logic;
  SIGNAL Logical_Operator_out5126_out1            : std_logic;
  SIGNAL Logical_Operator_out5127_out1            : std_logic;
  SIGNAL Logical_Operator_out5128_out1            : std_logic;
  SIGNAL Logical_Operator_out5129_out1            : std_logic;
  SIGNAL Logical_Operator_out5130_out1            : std_logic;
  SIGNAL Logical_Operator_out5131_out1            : std_logic;
  SIGNAL Logical_Operator_out5132_out1            : std_logic;
  SIGNAL Logical_Operator_out5133_out1            : std_logic;
  SIGNAL Logical_Operator_out5134_out1            : std_logic;
  SIGNAL Logical_Operator_out5135_out1            : std_logic;
  SIGNAL Logical_Operator_out5136_out1            : std_logic;
  SIGNAL Logical_Operator_out5137_out1            : std_logic;
  SIGNAL Logical_Operator_out5138_out1            : std_logic;
  SIGNAL Logical_Operator_out5139_out1            : std_logic;
  SIGNAL Logical_Operator_out5140_out1            : std_logic;
  SIGNAL Logical_Operator_out5141_out1            : std_logic;
  SIGNAL Logical_Operator_out5142_out1            : std_logic;
  SIGNAL Logical_Operator_out5143_out1            : std_logic;
  SIGNAL Logical_Operator_out5144_out1            : std_logic;
  SIGNAL Logical_Operator_out5145_out1            : std_logic;
  SIGNAL Logical_Operator_out5146_out1            : std_logic;
  SIGNAL Logical_Operator_out5147_out1            : std_logic;
  SIGNAL Logical_Operator_out5148_out1            : std_logic;
  SIGNAL Logical_Operator_out5149_out1            : std_logic;
  SIGNAL Logical_Operator_out5150_out1            : std_logic;
  SIGNAL Logical_Operator_out5151_out1            : std_logic;
  SIGNAL Logical_Operator_out5152_out1            : std_logic;
  SIGNAL Logical_Operator_out5153_out1            : std_logic;
  SIGNAL Logical_Operator_out5154_out1            : std_logic;
  SIGNAL Logical_Operator_out5155_out1            : std_logic;
  SIGNAL Logical_Operator_out5156_out1            : std_logic;
  SIGNAL Logical_Operator_out5157_out1            : std_logic;
  SIGNAL Logical_Operator_out5158_out1            : std_logic;
  SIGNAL Logical_Operator_out5159_out1            : std_logic;
  SIGNAL Logical_Operator_out5160_out1            : std_logic;
  SIGNAL Logical_Operator_out5161_out1            : std_logic;
  SIGNAL Logical_Operator_out5162_out1            : std_logic;
  SIGNAL Logical_Operator_out5163_out1            : std_logic;
  SIGNAL Logical_Operator_out5164_out1            : std_logic;
  SIGNAL Logical_Operator_out5165_out1            : std_logic;
  SIGNAL Logical_Operator_out5166_out1            : std_logic;
  SIGNAL Logical_Operator_out5167_out1            : std_logic;
  SIGNAL Logical_Operator_out5168_out1            : std_logic;
  SIGNAL Logical_Operator_out5169_out1            : std_logic;
  SIGNAL Logical_Operator_out5170_out1            : std_logic;
  SIGNAL Logical_Operator_out5171_out1            : std_logic;
  SIGNAL Logical_Operator_out5172_out1            : std_logic;
  SIGNAL Logical_Operator_out5173_out1            : std_logic;
  SIGNAL Logical_Operator_out5174_out1            : std_logic;
  SIGNAL Logical_Operator_out5175_out1            : std_logic;
  SIGNAL Logical_Operator_out5176_out1            : std_logic;
  SIGNAL Logical_Operator_out5177_out1            : std_logic;
  SIGNAL Logical_Operator_out5178_out1            : std_logic;
  SIGNAL Logical_Operator_out5179_out1            : std_logic;
  SIGNAL Logical_Operator_out5180_out1            : std_logic;
  SIGNAL Logical_Operator_out5181_out1            : std_logic;
  SIGNAL Logical_Operator_out5182_out1            : std_logic;
  SIGNAL Logical_Operator_out5183_out1            : std_logic;
  SIGNAL Logical_Operator_out5184_out1            : std_logic;
  SIGNAL Logical_Operator_out5185_out1            : std_logic;
  SIGNAL Logical_Operator_out5186_out1            : std_logic;
  SIGNAL Logical_Operator_out5187_out1            : std_logic;
  SIGNAL Logical_Operator_out5188_out1            : std_logic;
  SIGNAL Logical_Operator_out5189_out1            : std_logic;
  SIGNAL Logical_Operator_out5190_out1            : std_logic;
  SIGNAL Logical_Operator_out5191_out1            : std_logic;
  SIGNAL Logical_Operator_out5192_out1            : std_logic;
  SIGNAL Logical_Operator_out5193_out1            : std_logic;
  SIGNAL Logical_Operator_out5194_out1            : std_logic;
  SIGNAL Logical_Operator_out5195_out1            : std_logic;
  SIGNAL Logical_Operator_out5196_out1            : std_logic;
  SIGNAL Logical_Operator_out5197_out1            : std_logic;
  SIGNAL Logical_Operator_out5198_out1            : std_logic;
  SIGNAL Logical_Operator_out5199_out1            : std_logic;
  SIGNAL Logical_Operator_out5200_out1            : std_logic;
  SIGNAL Logical_Operator_out5201_out1            : std_logic;
  SIGNAL Logical_Operator_out5202_out1            : std_logic;
  SIGNAL Logical_Operator_out5203_out1            : std_logic;
  SIGNAL Logical_Operator_out5204_out1            : std_logic;
  SIGNAL Logical_Operator_out5205_out1            : std_logic;
  SIGNAL Logical_Operator_out5206_out1            : std_logic;
  SIGNAL Logical_Operator_out5207_out1            : std_logic;
  SIGNAL Logical_Operator_out5208_out1            : std_logic;
  SIGNAL Logical_Operator_out5209_out1            : std_logic;
  SIGNAL Logical_Operator_out5210_out1            : std_logic;
  SIGNAL Logical_Operator_out5211_out1            : std_logic;
  SIGNAL Logical_Operator_out5212_out1            : std_logic;
  SIGNAL Logical_Operator_out5213_out1            : std_logic;
  SIGNAL Logical_Operator_out5214_out1            : std_logic;
  SIGNAL Logical_Operator_out5215_out1            : std_logic;
  SIGNAL Logical_Operator_out5216_out1            : std_logic;
  SIGNAL Logical_Operator_out5217_out1            : std_logic;
  SIGNAL Logical_Operator_out5218_out1            : std_logic;
  SIGNAL Logical_Operator_out5219_out1            : std_logic;
  SIGNAL Logical_Operator_out5220_out1            : std_logic;
  SIGNAL Logical_Operator_out5221_out1            : std_logic;
  SIGNAL Logical_Operator_out5222_out1            : std_logic;
  SIGNAL Logical_Operator_out5223_out1            : std_logic;
  SIGNAL Logical_Operator_out5224_out1            : std_logic;
  SIGNAL Logical_Operator_out5225_out1            : std_logic;
  SIGNAL Logical_Operator_out5226_out1            : std_logic;
  SIGNAL Logical_Operator_out5227_out1            : std_logic;
  SIGNAL Logical_Operator_out5228_out1            : std_logic;
  SIGNAL Logical_Operator_out5229_out1            : std_logic;
  SIGNAL Logical_Operator_out5230_out1            : std_logic;
  SIGNAL Logical_Operator_out5231_out1            : std_logic;
  SIGNAL Logical_Operator_out5232_out1            : std_logic;
  SIGNAL Logical_Operator_out5233_out1            : std_logic;
  SIGNAL Logical_Operator_out5234_out1            : std_logic;
  SIGNAL Logical_Operator_out5235_out1            : std_logic;
  SIGNAL Logical_Operator_out5236_out1            : std_logic;
  SIGNAL Logical_Operator_out5237_out1            : std_logic;
  SIGNAL Logical_Operator_out5238_out1            : std_logic;
  SIGNAL Logical_Operator_out5239_out1            : std_logic;
  SIGNAL Logical_Operator_out5240_out1            : std_logic;
  SIGNAL Logical_Operator_out5241_out1            : std_logic;
  SIGNAL Logical_Operator_out5242_out1            : std_logic;
  SIGNAL Logical_Operator_out5243_out1            : std_logic;
  SIGNAL Logical_Operator_out5244_out1            : std_logic;
  SIGNAL Logical_Operator_out5245_out1            : std_logic;
  SIGNAL Logical_Operator_out5246_out1            : std_logic;
  SIGNAL Logical_Operator_out5247_out1            : std_logic;
  SIGNAL Logical_Operator_out5248_out1            : std_logic;
  SIGNAL Logical_Operator_out5249_out1            : std_logic;
  SIGNAL Logical_Operator_out5250_out1            : std_logic;
  SIGNAL Logical_Operator_out5251_out1            : std_logic;
  SIGNAL Logical_Operator_out5252_out1            : std_logic;
  SIGNAL Logical_Operator_out5253_out1            : std_logic;
  SIGNAL Logical_Operator_out5254_out1            : std_logic;
  SIGNAL Logical_Operator_out5255_out1            : std_logic;
  SIGNAL Logical_Operator_out5256_out1            : std_logic;
  SIGNAL Logical_Operator_out5257_out1            : std_logic;
  SIGNAL Logical_Operator_out5258_out1            : std_logic;
  SIGNAL Logical_Operator_out5259_out1            : std_logic;
  SIGNAL Logical_Operator_out5260_out1            : std_logic;
  SIGNAL Logical_Operator_out5261_out1            : std_logic;
  SIGNAL Logical_Operator_out5262_out1            : std_logic;
  SIGNAL Logical_Operator_out5263_out1            : std_logic;
  SIGNAL Logical_Operator_out5264_out1            : std_logic;
  SIGNAL Logical_Operator_out5265_out1            : std_logic;
  SIGNAL Logical_Operator_out5266_out1            : std_logic;
  SIGNAL Logical_Operator_out5267_out1            : std_logic;
  SIGNAL Logical_Operator_out5268_out1            : std_logic;
  SIGNAL Logical_Operator_out5269_out1            : std_logic;
  SIGNAL Logical_Operator_out5270_out1            : std_logic;
  SIGNAL Logical_Operator_out5271_out1            : std_logic;
  SIGNAL Logical_Operator_out5272_out1            : std_logic;
  SIGNAL Logical_Operator_out5273_out1            : std_logic;
  SIGNAL Logical_Operator_out5274_out1            : std_logic;
  SIGNAL Logical_Operator_out5275_out1            : std_logic;
  SIGNAL Logical_Operator_out5276_out1            : std_logic;
  SIGNAL Logical_Operator_out5277_out1            : std_logic;
  SIGNAL Logical_Operator_out5278_out1            : std_logic;
  SIGNAL Logical_Operator_out5279_out1            : std_logic;
  SIGNAL Logical_Operator_out5280_out1            : std_logic;
  SIGNAL Logical_Operator_out5281_out1            : std_logic;
  SIGNAL Logical_Operator_out5282_out1            : std_logic;
  SIGNAL Logical_Operator_out5283_out1            : std_logic;
  SIGNAL Logical_Operator_out5284_out1            : std_logic;
  SIGNAL Logical_Operator_out5285_out1            : std_logic;
  SIGNAL Logical_Operator_out5286_out1            : std_logic;
  SIGNAL Logical_Operator_out5287_out1            : std_logic;
  SIGNAL Logical_Operator_out5288_out1            : std_logic;
  SIGNAL Logical_Operator_out5289_out1            : std_logic;
  SIGNAL Logical_Operator_out5290_out1            : std_logic;
  SIGNAL Logical_Operator_out5291_out1            : std_logic;
  SIGNAL Logical_Operator_out5292_out1            : std_logic;
  SIGNAL Logical_Operator_out5293_out1            : std_logic;
  SIGNAL Logical_Operator_out5294_out1            : std_logic;
  SIGNAL Logical_Operator_out5295_out1            : std_logic;
  SIGNAL Logical_Operator_out5296_out1            : std_logic;
  SIGNAL Logical_Operator_out5297_out1            : std_logic;
  SIGNAL Logical_Operator_out5298_out1            : std_logic;
  SIGNAL Logical_Operator_out5299_out1            : std_logic;
  SIGNAL Logical_Operator_out5300_out1            : std_logic;
  SIGNAL Logical_Operator_out5301_out1            : std_logic;
  SIGNAL Logical_Operator_out5302_out1            : std_logic;
  SIGNAL Logical_Operator_out5303_out1            : std_logic;
  SIGNAL Logical_Operator_out5304_out1            : std_logic;
  SIGNAL Logical_Operator_out5305_out1            : std_logic;
  SIGNAL Logical_Operator_out5306_out1            : std_logic;
  SIGNAL Logical_Operator_out5307_out1            : std_logic;
  SIGNAL Logical_Operator_out5308_out1            : std_logic;
  SIGNAL Logical_Operator_out5309_out1            : std_logic;
  SIGNAL Logical_Operator_out5310_out1            : std_logic;
  SIGNAL Logical_Operator_out5311_out1            : std_logic;
  SIGNAL Logical_Operator_out5312_out1            : std_logic;
  SIGNAL Logical_Operator_out5313_out1            : std_logic;
  SIGNAL Logical_Operator_out5314_out1            : std_logic;
  SIGNAL Logical_Operator_out5315_out1            : std_logic;
  SIGNAL Logical_Operator_out5316_out1            : std_logic;
  SIGNAL Logical_Operator_out5317_out1            : std_logic;
  SIGNAL Logical_Operator_out5318_out1            : std_logic;
  SIGNAL Logical_Operator_out5319_out1            : std_logic;
  SIGNAL Logical_Operator_out5320_out1            : std_logic;
  SIGNAL Logical_Operator_out5321_out1            : std_logic;
  SIGNAL Logical_Operator_out5322_out1            : std_logic;
  SIGNAL Logical_Operator_out5323_out1            : std_logic;
  SIGNAL Logical_Operator_out5324_out1            : std_logic;
  SIGNAL Logical_Operator_out5325_out1            : std_logic;
  SIGNAL Logical_Operator_out5326_out1            : std_logic;
  SIGNAL Logical_Operator_out5327_out1            : std_logic;
  SIGNAL Logical_Operator_out5328_out1            : std_logic;
  SIGNAL Logical_Operator_out5329_out1            : std_logic;
  SIGNAL Logical_Operator_out5330_out1            : std_logic;
  SIGNAL Logical_Operator_out5331_out1            : std_logic;
  SIGNAL Logical_Operator_out5332_out1            : std_logic;
  SIGNAL Logical_Operator_out5333_out1            : std_logic;
  SIGNAL Logical_Operator_out5334_out1            : std_logic;
  SIGNAL Logical_Operator_out5335_out1            : std_logic;
  SIGNAL Logical_Operator_out5336_out1            : std_logic;
  SIGNAL Logical_Operator_out5337_out1            : std_logic;
  SIGNAL Logical_Operator_out5338_out1            : std_logic;
  SIGNAL Logical_Operator_out5339_out1            : std_logic;
  SIGNAL Logical_Operator_out5340_out1            : std_logic;
  SIGNAL Logical_Operator_out5341_out1            : std_logic;
  SIGNAL Logical_Operator_out5342_out1            : std_logic;
  SIGNAL Logical_Operator_out5343_out1            : std_logic;
  SIGNAL Logical_Operator_out5344_out1            : std_logic;
  SIGNAL Logical_Operator_out5345_out1            : std_logic;
  SIGNAL Logical_Operator_out5346_out1            : std_logic;
  SIGNAL Logical_Operator_out5347_out1            : std_logic;
  SIGNAL Logical_Operator_out5348_out1            : std_logic;
  SIGNAL Logical_Operator_out5349_out1            : std_logic;
  SIGNAL Logical_Operator_out5350_out1            : std_logic;
  SIGNAL Logical_Operator_out5351_out1            : std_logic;
  SIGNAL Logical_Operator_out5352_out1            : std_logic;
  SIGNAL Logical_Operator_out5353_out1            : std_logic;
  SIGNAL Logical_Operator_out5354_out1            : std_logic;
  SIGNAL Logical_Operator_out5355_out1            : std_logic;
  SIGNAL Logical_Operator_out5356_out1            : std_logic;
  SIGNAL Logical_Operator_out5357_out1            : std_logic;
  SIGNAL Logical_Operator_out5358_out1            : std_logic;
  SIGNAL Logical_Operator_out5359_out1            : std_logic;
  SIGNAL Logical_Operator_out5360_out1            : std_logic;
  SIGNAL Logical_Operator_out5361_out1            : std_logic;
  SIGNAL Logical_Operator_out5362_out1            : std_logic;
  SIGNAL Logical_Operator_out5363_out1            : std_logic;
  SIGNAL Logical_Operator_out5364_out1            : std_logic;
  SIGNAL Logical_Operator_out5365_out1            : std_logic;
  SIGNAL Logical_Operator_out5366_out1            : std_logic;
  SIGNAL Logical_Operator_out5367_out1            : std_logic;
  SIGNAL Logical_Operator_out5368_out1            : std_logic;
  SIGNAL Logical_Operator_out5369_out1            : std_logic;
  SIGNAL Logical_Operator_out5370_out1            : std_logic;
  SIGNAL Logical_Operator_out5371_out1            : std_logic;
  SIGNAL Logical_Operator_out5372_out1            : std_logic;
  SIGNAL Logical_Operator_out5373_out1            : std_logic;
  SIGNAL Logical_Operator_out5374_out1            : std_logic;
  SIGNAL Logical_Operator_out5375_out1            : std_logic;
  SIGNAL Logical_Operator_out5376_out1            : std_logic;
  SIGNAL Logical_Operator_out5377_out1            : std_logic;
  SIGNAL Logical_Operator_out5378_out1            : std_logic;
  SIGNAL Logical_Operator_out5379_out1            : std_logic;
  SIGNAL Logical_Operator_out5380_out1            : std_logic;
  SIGNAL Logical_Operator_out5381_out1            : std_logic;
  SIGNAL Logical_Operator_out5382_out1            : std_logic;
  SIGNAL Logical_Operator_out5383_out1            : std_logic;
  SIGNAL Logical_Operator_out5384_out1            : std_logic;
  SIGNAL Logical_Operator_out5385_out1            : std_logic;
  SIGNAL Logical_Operator_out5386_out1            : std_logic;
  SIGNAL Logical_Operator_out5387_out1            : std_logic;
  SIGNAL Logical_Operator_out5388_out1            : std_logic;
  SIGNAL Logical_Operator_out5389_out1            : std_logic;
  SIGNAL Logical_Operator_out5390_out1            : std_logic;
  SIGNAL Logical_Operator_out5391_out1            : std_logic;
  SIGNAL Logical_Operator_out5392_out1            : std_logic;
  SIGNAL Logical_Operator_out5393_out1            : std_logic;
  SIGNAL Logical_Operator_out5394_out1            : std_logic;
  SIGNAL Logical_Operator_out5395_out1            : std_logic;
  SIGNAL Logical_Operator_out5396_out1            : std_logic;
  SIGNAL Logical_Operator_out5397_out1            : std_logic;
  SIGNAL Logical_Operator_out5398_out1            : std_logic;
  SIGNAL Logical_Operator_out5399_out1            : std_logic;
  SIGNAL Logical_Operator_out5400_out1            : std_logic;
  SIGNAL Logical_Operator_out5401_out1            : std_logic;
  SIGNAL Logical_Operator_out5402_out1            : std_logic;
  SIGNAL Logical_Operator_out5403_out1            : std_logic;
  SIGNAL Logical_Operator_out5404_out1            : std_logic;
  SIGNAL Logical_Operator_out5405_out1            : std_logic;
  SIGNAL Logical_Operator_out5406_out1            : std_logic;
  SIGNAL Logical_Operator_out5407_out1            : std_logic;
  SIGNAL Logical_Operator_out5408_out1            : std_logic;
  SIGNAL Logical_Operator_out5409_out1            : std_logic;
  SIGNAL Logical_Operator_out5410_out1            : std_logic;
  SIGNAL Logical_Operator_out5411_out1            : std_logic;
  SIGNAL Logical_Operator_out5412_out1            : std_logic;
  SIGNAL Logical_Operator_out5413_out1            : std_logic;
  SIGNAL Logical_Operator_out5414_out1            : std_logic;
  SIGNAL Logical_Operator_out5415_out1            : std_logic;
  SIGNAL Logical_Operator_out5416_out1            : std_logic;
  SIGNAL Logical_Operator_out5417_out1            : std_logic;
  SIGNAL Logical_Operator_out5418_out1            : std_logic;
  SIGNAL Logical_Operator_out5419_out1            : std_logic;
  SIGNAL Logical_Operator_out5420_out1            : std_logic;
  SIGNAL Logical_Operator_out5421_out1            : std_logic;
  SIGNAL Logical_Operator_out5422_out1            : std_logic;
  SIGNAL Logical_Operator_out5423_out1            : std_logic;
  SIGNAL Logical_Operator_out5424_out1            : std_logic;
  SIGNAL Logical_Operator_out5425_out1            : std_logic;
  SIGNAL Logical_Operator_out5426_out1            : std_logic;
  SIGNAL Logical_Operator_out5427_out1            : std_logic;
  SIGNAL Logical_Operator_out5428_out1            : std_logic;
  SIGNAL Logical_Operator_out5429_out1            : std_logic;
  SIGNAL Logical_Operator_out5430_out1            : std_logic;
  SIGNAL Logical_Operator_out5431_out1            : std_logic;
  SIGNAL Logical_Operator_out5432_out1            : std_logic;
  SIGNAL Logical_Operator_out5433_out1            : std_logic;
  SIGNAL Logical_Operator_out5434_out1            : std_logic;
  SIGNAL Logical_Operator_out5435_out1            : std_logic;
  SIGNAL Logical_Operator_out5436_out1            : std_logic;
  SIGNAL Logical_Operator_out5437_out1            : std_logic;
  SIGNAL Logical_Operator_out5438_out1            : std_logic;
  SIGNAL Logical_Operator_out5439_out1            : std_logic;
  SIGNAL Logical_Operator_out5440_out1            : std_logic;
  SIGNAL Logical_Operator_out5441_out1            : std_logic;
  SIGNAL Logical_Operator_out5442_out1            : std_logic;
  SIGNAL Logical_Operator_out5443_out1            : std_logic;
  SIGNAL Logical_Operator_out5444_out1            : std_logic;
  SIGNAL Logical_Operator_out5445_out1            : std_logic;
  SIGNAL Logical_Operator_out5446_out1            : std_logic;
  SIGNAL Logical_Operator_out5447_out1            : std_logic;
  SIGNAL Logical_Operator_out5448_out1            : std_logic;
  SIGNAL Logical_Operator_out5449_out1            : std_logic;
  SIGNAL Logical_Operator_out5450_out1            : std_logic;
  SIGNAL Logical_Operator_out5451_out1            : std_logic;
  SIGNAL Logical_Operator_out5452_out1            : std_logic;
  SIGNAL Logical_Operator_out5453_out1            : std_logic;
  SIGNAL Logical_Operator_out5454_out1            : std_logic;
  SIGNAL Logical_Operator_out5455_out1            : std_logic;
  SIGNAL Logical_Operator_out5456_out1            : std_logic;
  SIGNAL Logical_Operator_out5457_out1            : std_logic;
  SIGNAL Logical_Operator_out5458_out1            : std_logic;
  SIGNAL Logical_Operator_out5459_out1            : std_logic;
  SIGNAL Logical_Operator_out5460_out1            : std_logic;
  SIGNAL Logical_Operator_out5461_out1            : std_logic;
  SIGNAL Logical_Operator_out5462_out1            : std_logic;
  SIGNAL Logical_Operator_out5463_out1            : std_logic;
  SIGNAL Logical_Operator_out5464_out1            : std_logic;
  SIGNAL Logical_Operator_out5465_out1            : std_logic;
  SIGNAL Logical_Operator_out5466_out1            : std_logic;
  SIGNAL Logical_Operator_out5467_out1            : std_logic;
  SIGNAL Logical_Operator_out5468_out1            : std_logic;
  SIGNAL Logical_Operator_out5469_out1            : std_logic;
  SIGNAL Logical_Operator_out5470_out1            : std_logic;
  SIGNAL Logical_Operator_out5471_out1            : std_logic;
  SIGNAL Logical_Operator_out5472_out1            : std_logic;
  SIGNAL Logical_Operator_out5473_out1            : std_logic;
  SIGNAL Logical_Operator_out5474_out1            : std_logic;
  SIGNAL Logical_Operator_out5475_out1            : std_logic;
  SIGNAL Logical_Operator_out5476_out1            : std_logic;
  SIGNAL Logical_Operator_out5477_out1            : std_logic;
  SIGNAL Logical_Operator_out5478_out1            : std_logic;
  SIGNAL Logical_Operator_out5479_out1            : std_logic;
  SIGNAL Logical_Operator_out5480_out1            : std_logic;
  SIGNAL Logical_Operator_out5481_out1            : std_logic;
  SIGNAL Logical_Operator_out5482_out1            : std_logic;
  SIGNAL Logical_Operator_out5483_out1            : std_logic;
  SIGNAL Logical_Operator_out5484_out1            : std_logic;
  SIGNAL Logical_Operator_out5485_out1            : std_logic;
  SIGNAL Logical_Operator_out5486_out1            : std_logic;
  SIGNAL Logical_Operator_out5487_out1            : std_logic;
  SIGNAL Logical_Operator_out5488_out1            : std_logic;
  SIGNAL Logical_Operator_out5489_out1            : std_logic;
  SIGNAL Logical_Operator_out5490_out1            : std_logic;
  SIGNAL Logical_Operator_out5491_out1            : std_logic;
  SIGNAL Logical_Operator_out5492_out1            : std_logic;
  SIGNAL Logical_Operator_out5493_out1            : std_logic;
  SIGNAL Logical_Operator_out5494_out1            : std_logic;
  SIGNAL Logical_Operator_out5495_out1            : std_logic;
  SIGNAL Logical_Operator_out5496_out1            : std_logic;
  SIGNAL Logical_Operator_out5497_out1            : std_logic;
  SIGNAL Logical_Operator_out5498_out1            : std_logic;
  SIGNAL Logical_Operator_out5499_out1            : std_logic;
  SIGNAL Logical_Operator_out5500_out1            : std_logic;
  SIGNAL Logical_Operator_out5501_out1            : std_logic;
  SIGNAL Logical_Operator_out5502_out1            : std_logic;
  SIGNAL Logical_Operator_out5503_out1            : std_logic;
  SIGNAL Logical_Operator_out5504_out1            : std_logic;
  SIGNAL Logical_Operator_out5505_out1            : std_logic;
  SIGNAL Logical_Operator_out5506_out1            : std_logic;
  SIGNAL Logical_Operator_out5507_out1            : std_logic;
  SIGNAL Logical_Operator_out5508_out1            : std_logic;
  SIGNAL Logical_Operator_out5509_out1            : std_logic;
  SIGNAL Logical_Operator_out5510_out1            : std_logic;
  SIGNAL Logical_Operator_out5511_out1            : std_logic;
  SIGNAL Logical_Operator_out5512_out1            : std_logic;
  SIGNAL Logical_Operator_out5513_out1            : std_logic;
  SIGNAL Logical_Operator_out5514_out1            : std_logic;
  SIGNAL Logical_Operator_out5515_out1            : std_logic;
  SIGNAL Logical_Operator_out5516_out1            : std_logic;
  SIGNAL Logical_Operator_out5517_out1            : std_logic;
  SIGNAL Logical_Operator_out5518_out1            : std_logic;
  SIGNAL Logical_Operator_out5519_out1            : std_logic;
  SIGNAL Logical_Operator_out5520_out1            : std_logic;
  SIGNAL Logical_Operator_out5521_out1            : std_logic;
  SIGNAL Logical_Operator_out5522_out1            : std_logic;
  SIGNAL Logical_Operator_out5523_out1            : std_logic;
  SIGNAL Logical_Operator_out5524_out1            : std_logic;
  SIGNAL Logical_Operator_out5525_out1            : std_logic;
  SIGNAL Logical_Operator_out5526_out1            : std_logic;
  SIGNAL Logical_Operator_out5527_out1            : std_logic;
  SIGNAL Logical_Operator_out5528_out1            : std_logic;
  SIGNAL Logical_Operator_out5529_out1            : std_logic;
  SIGNAL Logical_Operator_out5530_out1            : std_logic;
  SIGNAL Logical_Operator_out5531_out1            : std_logic;
  SIGNAL Logical_Operator_out5532_out1            : std_logic;
  SIGNAL Logical_Operator_out5533_out1            : std_logic;
  SIGNAL Logical_Operator_out5534_out1            : std_logic;
  SIGNAL Logical_Operator_out5535_out1            : std_logic;
  SIGNAL Logical_Operator_out5536_out1            : std_logic;
  SIGNAL Logical_Operator_out5537_out1            : std_logic;
  SIGNAL Logical_Operator_out5538_out1            : std_logic;
  SIGNAL Logical_Operator_out5539_out1            : std_logic;
  SIGNAL Logical_Operator_out5540_out1            : std_logic;
  SIGNAL Logical_Operator_out5541_out1            : std_logic;
  SIGNAL Logical_Operator_out5542_out1            : std_logic;
  SIGNAL Logical_Operator_out5543_out1            : std_logic;
  SIGNAL Logical_Operator_out5544_out1            : std_logic;
  SIGNAL Logical_Operator_out5545_out1            : std_logic;
  SIGNAL Logical_Operator_out5546_out1            : std_logic;
  SIGNAL Logical_Operator_out5547_out1            : std_logic;
  SIGNAL Logical_Operator_out5548_out1            : std_logic;
  SIGNAL Logical_Operator_out5549_out1            : std_logic;
  SIGNAL Logical_Operator_out5550_out1            : std_logic;
  SIGNAL Logical_Operator_out5551_out1            : std_logic;
  SIGNAL Logical_Operator_out5552_out1            : std_logic;
  SIGNAL Logical_Operator_out5553_out1            : std_logic;
  SIGNAL Logical_Operator_out5554_out1            : std_logic;
  SIGNAL Logical_Operator_out5555_out1            : std_logic;
  SIGNAL Logical_Operator_out5556_out1            : std_logic;
  SIGNAL Logical_Operator_out5557_out1            : std_logic;
  SIGNAL Logical_Operator_out5558_out1            : std_logic;
  SIGNAL Logical_Operator_out5559_out1            : std_logic;
  SIGNAL Logical_Operator_out5560_out1            : std_logic;
  SIGNAL Logical_Operator_out5561_out1            : std_logic;
  SIGNAL Logical_Operator_out5562_out1            : std_logic;
  SIGNAL Logical_Operator_out5563_out1            : std_logic;
  SIGNAL Logical_Operator_out5564_out1            : std_logic;
  SIGNAL Logical_Operator_out5565_out1            : std_logic;
  SIGNAL Logical_Operator_out5566_out1            : std_logic;
  SIGNAL Logical_Operator_out5567_out1            : std_logic;
  SIGNAL Logical_Operator_out5568_out1            : std_logic;
  SIGNAL Logical_Operator_out5569_out1            : std_logic;
  SIGNAL Logical_Operator_out5570_out1            : std_logic;
  SIGNAL Logical_Operator_out5571_out1            : std_logic;
  SIGNAL Logical_Operator_out5572_out1            : std_logic;
  SIGNAL Logical_Operator_out5573_out1            : std_logic;
  SIGNAL Logical_Operator_out5574_out1            : std_logic;
  SIGNAL Logical_Operator_out5575_out1            : std_logic;
  SIGNAL Logical_Operator_out5576_out1            : std_logic;
  SIGNAL Logical_Operator_out5577_out1            : std_logic;
  SIGNAL Logical_Operator_out5578_out1            : std_logic;
  SIGNAL Logical_Operator_out5579_out1            : std_logic;
  SIGNAL Logical_Operator_out5580_out1            : std_logic;
  SIGNAL Logical_Operator_out5581_out1            : std_logic;
  SIGNAL Logical_Operator_out5582_out1            : std_logic;
  SIGNAL Logical_Operator_out5583_out1            : std_logic;
  SIGNAL Logical_Operator_out5584_out1            : std_logic;
  SIGNAL Logical_Operator_out5585_out1            : std_logic;
  SIGNAL Logical_Operator_out5586_out1            : std_logic;
  SIGNAL Logical_Operator_out5587_out1            : std_logic;
  SIGNAL Logical_Operator_out5588_out1            : std_logic;
  SIGNAL Logical_Operator_out5589_out1            : std_logic;
  SIGNAL Logical_Operator_out5590_out1            : std_logic;
  SIGNAL Logical_Operator_out5591_out1            : std_logic;
  SIGNAL Logical_Operator_out5592_out1            : std_logic;
  SIGNAL Logical_Operator_out5593_out1            : std_logic;
  SIGNAL Logical_Operator_out5594_out1            : std_logic;
  SIGNAL Logical_Operator_out5595_out1            : std_logic;
  SIGNAL Logical_Operator_out5596_out1            : std_logic;
  SIGNAL Logical_Operator_out5597_out1            : std_logic;
  SIGNAL Logical_Operator_out5598_out1            : std_logic;
  SIGNAL Logical_Operator_out5599_out1            : std_logic;
  SIGNAL Logical_Operator_out5600_out1            : std_logic;
  SIGNAL Logical_Operator_out5601_out1            : std_logic;
  SIGNAL Logical_Operator_out5602_out1            : std_logic;
  SIGNAL Logical_Operator_out5603_out1            : std_logic;
  SIGNAL Logical_Operator_out5604_out1            : std_logic;
  SIGNAL Logical_Operator_out5605_out1            : std_logic;
  SIGNAL Logical_Operator_out5606_out1            : std_logic;
  SIGNAL Logical_Operator_out5607_out1            : std_logic;
  SIGNAL Logical_Operator_out5608_out1            : std_logic;
  SIGNAL Logical_Operator_out5609_out1            : std_logic;
  SIGNAL Logical_Operator_out5610_out1            : std_logic;
  SIGNAL Logical_Operator_out5611_out1            : std_logic;
  SIGNAL Logical_Operator_out5612_out1            : std_logic;
  SIGNAL Logical_Operator_out5613_out1            : std_logic;
  SIGNAL Logical_Operator_out5614_out1            : std_logic;
  SIGNAL Logical_Operator_out5615_out1            : std_logic;
  SIGNAL Logical_Operator_out5616_out1            : std_logic;
  SIGNAL Logical_Operator_out5617_out1            : std_logic;
  SIGNAL Logical_Operator_out5618_out1            : std_logic;
  SIGNAL Logical_Operator_out5619_out1            : std_logic;
  SIGNAL Logical_Operator_out5620_out1            : std_logic;
  SIGNAL Logical_Operator_out5621_out1            : std_logic;
  SIGNAL Logical_Operator_out5622_out1            : std_logic;
  SIGNAL Logical_Operator_out5623_out1            : std_logic;
  SIGNAL Logical_Operator_out5624_out1            : std_logic;
  SIGNAL Logical_Operator_out5625_out1            : std_logic;
  SIGNAL Logical_Operator_out5626_out1            : std_logic;
  SIGNAL Logical_Operator_out5627_out1            : std_logic;
  SIGNAL Logical_Operator_out5628_out1            : std_logic;
  SIGNAL Logical_Operator_out5629_out1            : std_logic;
  SIGNAL Logical_Operator_out5630_out1            : std_logic;
  SIGNAL Logical_Operator_out5631_out1            : std_logic;
  SIGNAL Logical_Operator_out5632_out1            : std_logic;
  SIGNAL Logical_Operator_out5633_out1            : std_logic;
  SIGNAL Logical_Operator_out5634_out1            : std_logic;
  SIGNAL Logical_Operator_out5635_out1            : std_logic;
  SIGNAL Logical_Operator_out5636_out1            : std_logic;
  SIGNAL Logical_Operator_out5637_out1            : std_logic;
  SIGNAL Logical_Operator_out5638_out1            : std_logic;
  SIGNAL Logical_Operator_out5639_out1            : std_logic;
  SIGNAL Logical_Operator_out5640_out1            : std_logic;
  SIGNAL Logical_Operator_out5641_out1            : std_logic;
  SIGNAL Logical_Operator_out5642_out1            : std_logic;
  SIGNAL Logical_Operator_out5643_out1            : std_logic;
  SIGNAL Logical_Operator_out5644_out1            : std_logic;
  SIGNAL Logical_Operator_out5645_out1            : std_logic;
  SIGNAL Logical_Operator_out5646_out1            : std_logic;
  SIGNAL Logical_Operator_out5647_out1            : std_logic;
  SIGNAL Logical_Operator_out5648_out1            : std_logic;
  SIGNAL Logical_Operator_out5649_out1            : std_logic;
  SIGNAL Logical_Operator_out5650_out1            : std_logic;
  SIGNAL Logical_Operator_out5651_out1            : std_logic;
  SIGNAL Logical_Operator_out5652_out1            : std_logic;
  SIGNAL Logical_Operator_out5653_out1            : std_logic;
  SIGNAL Logical_Operator_out5654_out1            : std_logic;
  SIGNAL Logical_Operator_out5655_out1            : std_logic;
  SIGNAL Logical_Operator_out5656_out1            : std_logic;
  SIGNAL Logical_Operator_out5657_out1            : std_logic;
  SIGNAL Logical_Operator_out5658_out1            : std_logic;
  SIGNAL Logical_Operator_out5659_out1            : std_logic;
  SIGNAL Logical_Operator_out5660_out1            : std_logic;
  SIGNAL Logical_Operator_out5661_out1            : std_logic;
  SIGNAL Logical_Operator_out5662_out1            : std_logic;
  SIGNAL Logical_Operator_out5663_out1            : std_logic;
  SIGNAL Logical_Operator_out5664_out1            : std_logic;
  SIGNAL Logical_Operator_out5665_out1            : std_logic;
  SIGNAL Logical_Operator_out5666_out1            : std_logic;
  SIGNAL Logical_Operator_out5667_out1            : std_logic;
  SIGNAL Logical_Operator_out5668_out1            : std_logic;
  SIGNAL Logical_Operator_out5669_out1            : std_logic;
  SIGNAL Logical_Operator_out5670_out1            : std_logic;
  SIGNAL Logical_Operator_out5671_out1            : std_logic;
  SIGNAL Logical_Operator_out5672_out1            : std_logic;
  SIGNAL Logical_Operator_out5673_out1            : std_logic;
  SIGNAL Logical_Operator_out5674_out1            : std_logic;
  SIGNAL Logical_Operator_out5675_out1            : std_logic;
  SIGNAL Logical_Operator_out5676_out1            : std_logic;
  SIGNAL Logical_Operator_out5677_out1            : std_logic;
  SIGNAL Logical_Operator_out5678_out1            : std_logic;
  SIGNAL Logical_Operator_out5679_out1            : std_logic;
  SIGNAL Logical_Operator_out5680_out1            : std_logic;
  SIGNAL Logical_Operator_out5681_out1            : std_logic;
  SIGNAL Logical_Operator_out5682_out1            : std_logic;
  SIGNAL Logical_Operator_out5683_out1            : std_logic;
  SIGNAL Logical_Operator_out5684_out1            : std_logic;
  SIGNAL Logical_Operator_out5685_out1            : std_logic;
  SIGNAL Logical_Operator_out5686_out1            : std_logic;
  SIGNAL Logical_Operator_out5687_out1            : std_logic;
  SIGNAL Logical_Operator_out5688_out1            : std_logic;
  SIGNAL Logical_Operator_out5689_out1            : std_logic;
  SIGNAL Logical_Operator_out5690_out1            : std_logic;
  SIGNAL Logical_Operator_out5691_out1            : std_logic;
  SIGNAL Logical_Operator_out5692_out1            : std_logic;
  SIGNAL Logical_Operator_out5693_out1            : std_logic;
  SIGNAL Logical_Operator_out5694_out1            : std_logic;
  SIGNAL Logical_Operator_out5695_out1            : std_logic;
  SIGNAL Logical_Operator_out5696_out1            : std_logic;
  SIGNAL Logical_Operator_out5697_out1            : std_logic;
  SIGNAL Logical_Operator_out5698_out1            : std_logic;
  SIGNAL Logical_Operator_out5699_out1            : std_logic;
  SIGNAL Logical_Operator_out5700_out1            : std_logic;
  SIGNAL Logical_Operator_out5701_out1            : std_logic;
  SIGNAL Logical_Operator_out5702_out1            : std_logic;
  SIGNAL Logical_Operator_out5703_out1            : std_logic;
  SIGNAL Logical_Operator_out5704_out1            : std_logic;
  SIGNAL Logical_Operator_out5705_out1            : std_logic;
  SIGNAL Logical_Operator_out5706_out1            : std_logic;
  SIGNAL Logical_Operator_out5707_out1            : std_logic;
  SIGNAL Logical_Operator_out5708_out1            : std_logic;
  SIGNAL Logical_Operator_out5709_out1            : std_logic;
  SIGNAL Logical_Operator_out5710_out1            : std_logic;
  SIGNAL Logical_Operator_out5711_out1            : std_logic;
  SIGNAL Logical_Operator_out5712_out1            : std_logic;
  SIGNAL Logical_Operator_out5713_out1            : std_logic;
  SIGNAL Logical_Operator_out5714_out1            : std_logic;
  SIGNAL Logical_Operator_out5715_out1            : std_logic;
  SIGNAL Logical_Operator_out5716_out1            : std_logic;
  SIGNAL Logical_Operator_out5717_out1            : std_logic;
  SIGNAL Logical_Operator_out5718_out1            : std_logic;
  SIGNAL Logical_Operator_out5719_out1            : std_logic;
  SIGNAL Logical_Operator_out5720_out1            : std_logic;
  SIGNAL Logical_Operator_out5721_out1            : std_logic;
  SIGNAL Logical_Operator_out5722_out1            : std_logic;
  SIGNAL Logical_Operator_out5723_out1            : std_logic;
  SIGNAL Logical_Operator_out5724_out1            : std_logic;
  SIGNAL Logical_Operator_out5725_out1            : std_logic;
  SIGNAL Logical_Operator_out5726_out1            : std_logic;
  SIGNAL Logical_Operator_out5727_out1            : std_logic;
  SIGNAL Logical_Operator_out5728_out1            : std_logic;
  SIGNAL Logical_Operator_out5729_out1            : std_logic;
  SIGNAL Logical_Operator_out5730_out1            : std_logic;
  SIGNAL Logical_Operator_out5731_out1            : std_logic;
  SIGNAL Logical_Operator_out5732_out1            : std_logic;
  SIGNAL Logical_Operator_out5733_out1            : std_logic;
  SIGNAL Logical_Operator_out5734_out1            : std_logic;
  SIGNAL Logical_Operator_out5735_out1            : std_logic;
  SIGNAL Logical_Operator_out5736_out1            : std_logic;
  SIGNAL Logical_Operator_out5737_out1            : std_logic;
  SIGNAL Logical_Operator_out5738_out1            : std_logic;
  SIGNAL Logical_Operator_out5739_out1            : std_logic;
  SIGNAL Logical_Operator_out5740_out1            : std_logic;
  SIGNAL Logical_Operator_out5741_out1            : std_logic;
  SIGNAL Logical_Operator_out5742_out1            : std_logic;
  SIGNAL Logical_Operator_out5743_out1            : std_logic;
  SIGNAL Logical_Operator_out5744_out1            : std_logic;
  SIGNAL Logical_Operator_out5745_out1            : std_logic;
  SIGNAL Logical_Operator_out5746_out1            : std_logic;
  SIGNAL Logical_Operator_out5747_out1            : std_logic;
  SIGNAL Logical_Operator_out5748_out1            : std_logic;
  SIGNAL Logical_Operator_out5749_out1            : std_logic;
  SIGNAL Logical_Operator_out5750_out1            : std_logic;
  SIGNAL Logical_Operator_out5751_out1            : std_logic;
  SIGNAL Logical_Operator_out5752_out1            : std_logic;
  SIGNAL Logical_Operator_out5753_out1            : std_logic;
  SIGNAL Logical_Operator_out5754_out1            : std_logic;
  SIGNAL Logical_Operator_out5755_out1            : std_logic;
  SIGNAL Logical_Operator_out5756_out1            : std_logic;
  SIGNAL Logical_Operator_out5757_out1            : std_logic;
  SIGNAL Logical_Operator_out5758_out1            : std_logic;
  SIGNAL Logical_Operator_out5759_out1            : std_logic;
  SIGNAL Logical_Operator_out5760_out1            : std_logic;
  SIGNAL Logical_Operator_out5761_out1            : std_logic;
  SIGNAL Logical_Operator_out5762_out1            : std_logic;
  SIGNAL Logical_Operator_out5763_out1            : std_logic;
  SIGNAL Logical_Operator_out5764_out1            : std_logic;
  SIGNAL Logical_Operator_out5765_out1            : std_logic;
  SIGNAL Logical_Operator_out5766_out1            : std_logic;
  SIGNAL Logical_Operator_out5767_out1            : std_logic;
  SIGNAL Logical_Operator_out5768_out1            : std_logic;
  SIGNAL Logical_Operator_out5769_out1            : std_logic;
  SIGNAL Logical_Operator_out5770_out1            : std_logic;
  SIGNAL Logical_Operator_out5771_out1            : std_logic;
  SIGNAL Logical_Operator_out5772_out1            : std_logic;
  SIGNAL Logical_Operator_out5773_out1            : std_logic;
  SIGNAL Logical_Operator_out5774_out1            : std_logic;
  SIGNAL Logical_Operator_out5775_out1            : std_logic;
  SIGNAL Logical_Operator_out5776_out1            : std_logic;
  SIGNAL Logical_Operator_out5777_out1            : std_logic;
  SIGNAL Logical_Operator_out5778_out1            : std_logic;
  SIGNAL Logical_Operator_out5779_out1            : std_logic;
  SIGNAL Logical_Operator_out5780_out1            : std_logic;
  SIGNAL Logical_Operator_out5781_out1            : std_logic;
  SIGNAL Logical_Operator_out5782_out1            : std_logic;
  SIGNAL Logical_Operator_out5783_out1            : std_logic;
  SIGNAL Logical_Operator_out5784_out1            : std_logic;
  SIGNAL Logical_Operator_out5785_out1            : std_logic;
  SIGNAL Logical_Operator_out5786_out1            : std_logic;
  SIGNAL Logical_Operator_out5787_out1            : std_logic;
  SIGNAL Logical_Operator_out5788_out1            : std_logic;
  SIGNAL Logical_Operator_out5789_out1            : std_logic;
  SIGNAL Logical_Operator_out5790_out1            : std_logic;
  SIGNAL Logical_Operator_out5791_out1            : std_logic;
  SIGNAL Logical_Operator_out5792_out1            : std_logic;
  SIGNAL Logical_Operator_out5793_out1            : std_logic;
  SIGNAL Logical_Operator_out5794_out1            : std_logic;
  SIGNAL Logical_Operator_out5795_out1            : std_logic;
  SIGNAL Logical_Operator_out5796_out1            : std_logic;
  SIGNAL Logical_Operator_out5797_out1            : std_logic;
  SIGNAL Logical_Operator_out5798_out1            : std_logic;
  SIGNAL Logical_Operator_out5799_out1            : std_logic;
  SIGNAL Logical_Operator_out5800_out1            : std_logic;
  SIGNAL Logical_Operator_out5801_out1            : std_logic;
  SIGNAL Logical_Operator_out5802_out1            : std_logic;
  SIGNAL Logical_Operator_out5803_out1            : std_logic;
  SIGNAL Logical_Operator_out5804_out1            : std_logic;
  SIGNAL Logical_Operator_out5805_out1            : std_logic;
  SIGNAL Logical_Operator_out5806_out1            : std_logic;
  SIGNAL Logical_Operator_out5807_out1            : std_logic;
  SIGNAL Logical_Operator_out5808_out1            : std_logic;
  SIGNAL Logical_Operator_out5809_out1            : std_logic;
  SIGNAL Logical_Operator_out5810_out1            : std_logic;
  SIGNAL Logical_Operator_out5811_out1            : std_logic;
  SIGNAL Logical_Operator_out5812_out1            : std_logic;
  SIGNAL Logical_Operator_out5813_out1            : std_logic;
  SIGNAL Logical_Operator_out5814_out1            : std_logic;
  SIGNAL Logical_Operator_out5815_out1            : std_logic;
  SIGNAL Logical_Operator_out5816_out1            : std_logic;
  SIGNAL Logical_Operator_out5817_out1            : std_logic;
  SIGNAL Logical_Operator_out5818_out1            : std_logic;
  SIGNAL Logical_Operator_out5819_out1            : std_logic;
  SIGNAL Logical_Operator_out5820_out1            : std_logic;
  SIGNAL Logical_Operator_out5821_out1            : std_logic;
  SIGNAL Logical_Operator_out5822_out1            : std_logic;
  SIGNAL Logical_Operator_out5823_out1            : std_logic;
  SIGNAL Logical_Operator_out5824_out1            : std_logic;
  SIGNAL Logical_Operator_out5825_out1            : std_logic;
  SIGNAL Logical_Operator_out5826_out1            : std_logic;
  SIGNAL Logical_Operator_out5827_out1            : std_logic;
  SIGNAL Logical_Operator_out5828_out1            : std_logic;
  SIGNAL Logical_Operator_out5829_out1            : std_logic;
  SIGNAL Logical_Operator_out5830_out1            : std_logic;
  SIGNAL Logical_Operator_out5831_out1            : std_logic;
  SIGNAL Logical_Operator_out5832_out1            : std_logic;
  SIGNAL Logical_Operator_out5833_out1            : std_logic;
  SIGNAL Logical_Operator_out5834_out1            : std_logic;
  SIGNAL Logical_Operator_out5835_out1            : std_logic;
  SIGNAL Logical_Operator_out5836_out1            : std_logic;
  SIGNAL Logical_Operator_out5837_out1            : std_logic;
  SIGNAL Logical_Operator_out5838_out1            : std_logic;
  SIGNAL Logical_Operator_out5839_out1            : std_logic;
  SIGNAL Logical_Operator_out5840_out1            : std_logic;
  SIGNAL Logical_Operator_out5841_out1            : std_logic;
  SIGNAL Logical_Operator_out5842_out1            : std_logic;
  SIGNAL Logical_Operator_out5843_out1            : std_logic;
  SIGNAL Logical_Operator_out5844_out1            : std_logic;
  SIGNAL Logical_Operator_out5845_out1            : std_logic;
  SIGNAL Logical_Operator_out5846_out1            : std_logic;
  SIGNAL Logical_Operator_out5847_out1            : std_logic;
  SIGNAL Logical_Operator_out5848_out1            : std_logic;
  SIGNAL Logical_Operator_out5849_out1            : std_logic;
  SIGNAL Logical_Operator_out5850_out1            : std_logic;
  SIGNAL Logical_Operator_out5851_out1            : std_logic;
  SIGNAL Logical_Operator_out5852_out1            : std_logic;
  SIGNAL Logical_Operator_out5853_out1            : std_logic;
  SIGNAL Logical_Operator_out5854_out1            : std_logic;
  SIGNAL Logical_Operator_out5855_out1            : std_logic;
  SIGNAL Logical_Operator_out5856_out1            : std_logic;
  SIGNAL Logical_Operator_out5857_out1            : std_logic;
  SIGNAL Logical_Operator_out5858_out1            : std_logic;
  SIGNAL Logical_Operator_out5859_out1            : std_logic;
  SIGNAL Logical_Operator_out5860_out1            : std_logic;
  SIGNAL Logical_Operator_out5861_out1            : std_logic;
  SIGNAL Logical_Operator_out5862_out1            : std_logic;
  SIGNAL Logical_Operator_out5863_out1            : std_logic;
  SIGNAL Logical_Operator_out5864_out1            : std_logic;
  SIGNAL Logical_Operator_out5865_out1            : std_logic;
  SIGNAL Logical_Operator_out5866_out1            : std_logic;
  SIGNAL Logical_Operator_out5867_out1            : std_logic;
  SIGNAL Logical_Operator_out5868_out1            : std_logic;
  SIGNAL Logical_Operator_out5869_out1            : std_logic;
  SIGNAL Logical_Operator_out5870_out1            : std_logic;
  SIGNAL Logical_Operator_out5871_out1            : std_logic;
  SIGNAL Logical_Operator_out5872_out1            : std_logic;
  SIGNAL Logical_Operator_out5873_out1            : std_logic;
  SIGNAL Logical_Operator_out5874_out1            : std_logic;
  SIGNAL Logical_Operator_out5875_out1            : std_logic;
  SIGNAL Logical_Operator_out5876_out1            : std_logic;
  SIGNAL Logical_Operator_out5877_out1            : std_logic;
  SIGNAL Logical_Operator_out5878_out1            : std_logic;
  SIGNAL Logical_Operator_out5879_out1            : std_logic;
  SIGNAL Logical_Operator_out5880_out1            : std_logic;
  SIGNAL Logical_Operator_out5881_out1            : std_logic;
  SIGNAL Logical_Operator_out5882_out1            : std_logic;
  SIGNAL Logical_Operator_out5883_out1            : std_logic;
  SIGNAL Logical_Operator_out5884_out1            : std_logic;
  SIGNAL Logical_Operator_out5885_out1            : std_logic;
  SIGNAL Logical_Operator_out5886_out1            : std_logic;
  SIGNAL Logical_Operator_out5887_out1            : std_logic;
  SIGNAL Logical_Operator_out5888_out1            : std_logic;
  SIGNAL Logical_Operator_out5889_out1            : std_logic;
  SIGNAL Logical_Operator_out5890_out1            : std_logic;
  SIGNAL Logical_Operator_out5891_out1            : std_logic;
  SIGNAL Logical_Operator_out5892_out1            : std_logic;
  SIGNAL Logical_Operator_out5893_out1            : std_logic;
  SIGNAL Logical_Operator_out5894_out1            : std_logic;
  SIGNAL Logical_Operator_out5895_out1            : std_logic;
  SIGNAL Logical_Operator_out5896_out1            : std_logic;
  SIGNAL Logical_Operator_out5897_out1            : std_logic;
  SIGNAL Logical_Operator_out5898_out1            : std_logic;
  SIGNAL Logical_Operator_out5899_out1            : std_logic;
  SIGNAL Logical_Operator_out5900_out1            : std_logic;
  SIGNAL Logical_Operator_out5901_out1            : std_logic;
  SIGNAL Logical_Operator_out5902_out1            : std_logic;
  SIGNAL Logical_Operator_out5903_out1            : std_logic;
  SIGNAL Logical_Operator_out5904_out1            : std_logic;
  SIGNAL Logical_Operator_out5905_out1            : std_logic;
  SIGNAL Logical_Operator_out5906_out1            : std_logic;
  SIGNAL Logical_Operator_out5907_out1            : std_logic;
  SIGNAL Logical_Operator_out5908_out1            : std_logic;
  SIGNAL Logical_Operator_out5909_out1            : std_logic;
  SIGNAL Logical_Operator_out5910_out1            : std_logic;
  SIGNAL Logical_Operator_out5911_out1            : std_logic;
  SIGNAL Logical_Operator_out5912_out1            : std_logic;
  SIGNAL Logical_Operator_out5913_out1            : std_logic;
  SIGNAL Logical_Operator_out5914_out1            : std_logic;
  SIGNAL Logical_Operator_out5915_out1            : std_logic;
  SIGNAL Logical_Operator_out5916_out1            : std_logic;
  SIGNAL Logical_Operator_out5917_out1            : std_logic;
  SIGNAL Logical_Operator_out5918_out1            : std_logic;
  SIGNAL Logical_Operator_out5919_out1            : std_logic;
  SIGNAL Logical_Operator_out5920_out1            : std_logic;
  SIGNAL Logical_Operator_out5921_out1            : std_logic;
  SIGNAL Logical_Operator_out5922_out1            : std_logic;
  SIGNAL Logical_Operator_out5923_out1            : std_logic;
  SIGNAL Logical_Operator_out5924_out1            : std_logic;
  SIGNAL Logical_Operator_out5925_out1            : std_logic;
  SIGNAL Logical_Operator_out5926_out1            : std_logic;
  SIGNAL Logical_Operator_out5927_out1            : std_logic;
  SIGNAL Logical_Operator_out5928_out1            : std_logic;
  SIGNAL Logical_Operator_out5929_out1            : std_logic;
  SIGNAL Logical_Operator_out5930_out1            : std_logic;
  SIGNAL Logical_Operator_out5931_out1            : std_logic;
  SIGNAL Logical_Operator_out5932_out1            : std_logic;
  SIGNAL Logical_Operator_out5933_out1            : std_logic;
  SIGNAL Logical_Operator_out5934_out1            : std_logic;
  SIGNAL Logical_Operator_out5935_out1            : std_logic;
  SIGNAL Logical_Operator_out5936_out1            : std_logic;
  SIGNAL Logical_Operator_out5937_out1            : std_logic;
  SIGNAL Logical_Operator_out5938_out1            : std_logic;
  SIGNAL Logical_Operator_out5939_out1            : std_logic;
  SIGNAL Logical_Operator_out5940_out1            : std_logic;
  SIGNAL Logical_Operator_out5941_out1            : std_logic;
  SIGNAL Logical_Operator_out5942_out1            : std_logic;
  SIGNAL Logical_Operator_out5943_out1            : std_logic;
  SIGNAL Logical_Operator_out5944_out1            : std_logic;
  SIGNAL Logical_Operator_out5945_out1            : std_logic;
  SIGNAL Logical_Operator_out5946_out1            : std_logic;
  SIGNAL Logical_Operator_out5947_out1            : std_logic;
  SIGNAL Logical_Operator_out5948_out1            : std_logic;
  SIGNAL Logical_Operator_out5949_out1            : std_logic;
  SIGNAL Logical_Operator_out5950_out1            : std_logic;
  SIGNAL Logical_Operator_out5951_out1            : std_logic;
  SIGNAL Logical_Operator_out5952_out1            : std_logic;
  SIGNAL Logical_Operator_out5953_out1            : std_logic;
  SIGNAL Logical_Operator_out5954_out1            : std_logic;
  SIGNAL Logical_Operator_out5955_out1            : std_logic;
  SIGNAL Logical_Operator_out5956_out1            : std_logic;
  SIGNAL Logical_Operator_out5957_out1            : std_logic;
  SIGNAL Logical_Operator_out5958_out1            : std_logic;
  SIGNAL Logical_Operator_out5959_out1            : std_logic;
  SIGNAL Logical_Operator_out5960_out1            : std_logic;
  SIGNAL Logical_Operator_out5961_out1            : std_logic;
  SIGNAL Logical_Operator_out5962_out1            : std_logic;
  SIGNAL Logical_Operator_out5963_out1            : std_logic;
  SIGNAL Logical_Operator_out5964_out1            : std_logic;
  SIGNAL Logical_Operator_out5965_out1            : std_logic;
  SIGNAL Logical_Operator_out5966_out1            : std_logic;
  SIGNAL Logical_Operator_out5967_out1            : std_logic;
  SIGNAL Logical_Operator_out5968_out1            : std_logic;
  SIGNAL Logical_Operator_out5969_out1            : std_logic;
  SIGNAL Logical_Operator_out5970_out1            : std_logic;
  SIGNAL Logical_Operator_out5971_out1            : std_logic;
  SIGNAL Logical_Operator_out5972_out1            : std_logic;
  SIGNAL Logical_Operator_out5973_out1            : std_logic;
  SIGNAL Logical_Operator_out5974_out1            : std_logic;
  SIGNAL Logical_Operator_out5975_out1            : std_logic;
  SIGNAL Logical_Operator_out5976_out1            : std_logic;
  SIGNAL Logical_Operator_out5977_out1            : std_logic;
  SIGNAL Logical_Operator_out5978_out1            : std_logic;
  SIGNAL Logical_Operator_out5979_out1            : std_logic;
  SIGNAL Logical_Operator_out5980_out1            : std_logic;
  SIGNAL Logical_Operator_out5981_out1            : std_logic;
  SIGNAL Logical_Operator_out5982_out1            : std_logic;
  SIGNAL Logical_Operator_out5983_out1            : std_logic;
  SIGNAL Logical_Operator_out5984_out1            : std_logic;
  SIGNAL Logical_Operator_out5985_out1            : std_logic;
  SIGNAL Logical_Operator_out5986_out1            : std_logic;
  SIGNAL Logical_Operator_out5987_out1            : std_logic;
  SIGNAL Logical_Operator_out5988_out1            : std_logic;
  SIGNAL Logical_Operator_out5989_out1            : std_logic;
  SIGNAL Logical_Operator_out5990_out1            : std_logic;
  SIGNAL Logical_Operator_out5991_out1            : std_logic;
  SIGNAL Logical_Operator_out5992_out1            : std_logic;
  SIGNAL Logical_Operator_out5993_out1            : std_logic;
  SIGNAL Logical_Operator_out5994_out1            : std_logic;
  SIGNAL Logical_Operator_out5995_out1            : std_logic;
  SIGNAL Logical_Operator_out5996_out1            : std_logic;
  SIGNAL Logical_Operator_out5997_out1            : std_logic;
  SIGNAL Logical_Operator_out5998_out1            : std_logic;
  SIGNAL Logical_Operator_out5999_out1            : std_logic;
  SIGNAL Logical_Operator_out6000_out1            : std_logic;
  SIGNAL Logical_Operator_out6001_out1            : std_logic;
  SIGNAL Logical_Operator_out6002_out1            : std_logic;
  SIGNAL Logical_Operator_out6003_out1            : std_logic;
  SIGNAL Logical_Operator_out6004_out1            : std_logic;
  SIGNAL Logical_Operator_out6005_out1            : std_logic;
  SIGNAL Logical_Operator_out6006_out1            : std_logic;
  SIGNAL Logical_Operator_out6007_out1            : std_logic;
  SIGNAL Logical_Operator_out6008_out1            : std_logic;
  SIGNAL Logical_Operator_out6009_out1            : std_logic;
  SIGNAL Logical_Operator_out6010_out1            : std_logic;
  SIGNAL Logical_Operator_out6011_out1            : std_logic;
  SIGNAL Logical_Operator_out6012_out1            : std_logic;
  SIGNAL Logical_Operator_out6013_out1            : std_logic;
  SIGNAL Logical_Operator_out6014_out1            : std_logic;
  SIGNAL Logical_Operator_out6015_out1            : std_logic;
  SIGNAL Logical_Operator_out6016_out1            : std_logic;
  SIGNAL Logical_Operator_out6017_out1            : std_logic;
  SIGNAL Logical_Operator_out6018_out1            : std_logic;
  SIGNAL Logical_Operator_out6019_out1            : std_logic;
  SIGNAL Logical_Operator_out6020_out1            : std_logic;
  SIGNAL Logical_Operator_out6021_out1            : std_logic;
  SIGNAL Logical_Operator_out6022_out1            : std_logic;
  SIGNAL Logical_Operator_out6023_out1            : std_logic;
  SIGNAL Logical_Operator_out6024_out1            : std_logic;
  SIGNAL Logical_Operator_out6025_out1            : std_logic;
  SIGNAL Logical_Operator_out6026_out1            : std_logic;
  SIGNAL Logical_Operator_out6027_out1            : std_logic;
  SIGNAL Logical_Operator_out6028_out1            : std_logic;
  SIGNAL Logical_Operator_out6029_out1            : std_logic;
  SIGNAL Logical_Operator_out6030_out1            : std_logic;
  SIGNAL Logical_Operator_out6031_out1            : std_logic;
  SIGNAL Logical_Operator_out6032_out1            : std_logic;
  SIGNAL Logical_Operator_out6033_out1            : std_logic;
  SIGNAL Logical_Operator_out6034_out1            : std_logic;
  SIGNAL Logical_Operator_out6035_out1            : std_logic;
  SIGNAL Logical_Operator_out6036_out1            : std_logic;
  SIGNAL Logical_Operator_out6037_out1            : std_logic;
  SIGNAL Logical_Operator_out6038_out1            : std_logic;
  SIGNAL Logical_Operator_out6039_out1            : std_logic;
  SIGNAL Logical_Operator_out6040_out1            : std_logic;
  SIGNAL Logical_Operator_out6041_out1            : std_logic;
  SIGNAL Logical_Operator_out6042_out1            : std_logic;
  SIGNAL Logical_Operator_out6043_out1            : std_logic;
  SIGNAL Logical_Operator_out6044_out1            : std_logic;
  SIGNAL Logical_Operator_out6045_out1            : std_logic;
  SIGNAL Logical_Operator_out6046_out1            : std_logic;
  SIGNAL Logical_Operator_out6047_out1            : std_logic;
  SIGNAL Logical_Operator_out6048_out1            : std_logic;
  SIGNAL Logical_Operator_out6049_out1            : std_logic;
  SIGNAL Logical_Operator_out6050_out1            : std_logic;
  SIGNAL Logical_Operator_out6051_out1            : std_logic;
  SIGNAL Logical_Operator_out6052_out1            : std_logic;
  SIGNAL Logical_Operator_out6053_out1            : std_logic;
  SIGNAL Logical_Operator_out6054_out1            : std_logic;
  SIGNAL Logical_Operator_out6055_out1            : std_logic;
  SIGNAL Logical_Operator_out6056_out1            : std_logic;
  SIGNAL Logical_Operator_out6057_out1            : std_logic;
  SIGNAL Logical_Operator_out6058_out1            : std_logic;
  SIGNAL Logical_Operator_out6059_out1            : std_logic;
  SIGNAL Logical_Operator_out6060_out1            : std_logic;
  SIGNAL Logical_Operator_out6061_out1            : std_logic;
  SIGNAL Logical_Operator_out6062_out1            : std_logic;
  SIGNAL Logical_Operator_out6063_out1            : std_logic;
  SIGNAL Logical_Operator_out6064_out1            : std_logic;
  SIGNAL Logical_Operator_out6065_out1            : std_logic;
  SIGNAL Logical_Operator_out6066_out1            : std_logic;
  SIGNAL Logical_Operator_out6067_out1            : std_logic;
  SIGNAL Logical_Operator_out6068_out1            : std_logic;
  SIGNAL Logical_Operator_out6069_out1            : std_logic;
  SIGNAL Logical_Operator_out6070_out1            : std_logic;
  SIGNAL Logical_Operator_out6071_out1            : std_logic;
  SIGNAL Logical_Operator_out6072_out1            : std_logic;
  SIGNAL Logical_Operator_out6073_out1            : std_logic;
  SIGNAL Logical_Operator_out6074_out1            : std_logic;
  SIGNAL Logical_Operator_out6075_out1            : std_logic;
  SIGNAL Logical_Operator_out6076_out1            : std_logic;
  SIGNAL Logical_Operator_out6077_out1            : std_logic;
  SIGNAL Logical_Operator_out6078_out1            : std_logic;
  SIGNAL Logical_Operator_out6079_out1            : std_logic;
  SIGNAL Logical_Operator_out6080_out1            : std_logic;
  SIGNAL Logical_Operator_out6081_out1            : std_logic;
  SIGNAL Logical_Operator_out6082_out1            : std_logic;
  SIGNAL Logical_Operator_out6083_out1            : std_logic;
  SIGNAL Logical_Operator_out6084_out1            : std_logic;
  SIGNAL Logical_Operator_out6085_out1            : std_logic;
  SIGNAL Logical_Operator_out6086_out1            : std_logic;
  SIGNAL Logical_Operator_out6087_out1            : std_logic;
  SIGNAL Logical_Operator_out6088_out1            : std_logic;
  SIGNAL Logical_Operator_out6089_out1            : std_logic;
  SIGNAL Logical_Operator_out6090_out1            : std_logic;
  SIGNAL Logical_Operator_out6091_out1            : std_logic;
  SIGNAL Logical_Operator_out6092_out1            : std_logic;
  SIGNAL Logical_Operator_out6093_out1            : std_logic;
  SIGNAL Logical_Operator_out6094_out1            : std_logic;
  SIGNAL Logical_Operator_out6095_out1            : std_logic;
  SIGNAL Logical_Operator_out6096_out1            : std_logic;
  SIGNAL Logical_Operator_out6097_out1            : std_logic;
  SIGNAL Logical_Operator_out6098_out1            : std_logic;
  SIGNAL Logical_Operator_out6099_out1            : std_logic;
  SIGNAL Logical_Operator_out6100_out1            : std_logic;
  SIGNAL Logical_Operator_out6101_out1            : std_logic;
  SIGNAL Logical_Operator_out6102_out1            : std_logic;
  SIGNAL Logical_Operator_out6103_out1            : std_logic;
  SIGNAL Logical_Operator_out6104_out1            : std_logic;
  SIGNAL Logical_Operator_out6105_out1            : std_logic;
  SIGNAL Logical_Operator_out6106_out1            : std_logic;
  SIGNAL Logical_Operator_out6107_out1            : std_logic;
  SIGNAL Logical_Operator_out6108_out1            : std_logic;
  SIGNAL Logical_Operator_out6109_out1            : std_logic;
  SIGNAL Logical_Operator_out6110_out1            : std_logic;
  SIGNAL Logical_Operator_out6111_out1            : std_logic;
  SIGNAL Logical_Operator_out6112_out1            : std_logic;
  SIGNAL Logical_Operator_out6113_out1            : std_logic;
  SIGNAL Logical_Operator_out6114_out1            : std_logic;
  SIGNAL Logical_Operator_out6115_out1            : std_logic;
  SIGNAL Logical_Operator_out6116_out1            : std_logic;
  SIGNAL Logical_Operator_out6117_out1            : std_logic;
  SIGNAL Logical_Operator_out6118_out1            : std_logic;
  SIGNAL Logical_Operator_out6119_out1            : std_logic;
  SIGNAL Logical_Operator_out6120_out1            : std_logic;
  SIGNAL Logical_Operator_out6121_out1            : std_logic;
  SIGNAL Logical_Operator_out6122_out1            : std_logic;
  SIGNAL Logical_Operator_out6123_out1            : std_logic;
  SIGNAL Logical_Operator_out6124_out1            : std_logic;
  SIGNAL Logical_Operator_out6125_out1            : std_logic;
  SIGNAL Logical_Operator_out6126_out1            : std_logic;
  SIGNAL Logical_Operator_out6127_out1            : std_logic;
  SIGNAL Logical_Operator_out6128_out1            : std_logic;
  SIGNAL Logical_Operator_out6129_out1            : std_logic;
  SIGNAL Logical_Operator_out6130_out1            : std_logic;
  SIGNAL Logical_Operator_out6131_out1            : std_logic;
  SIGNAL Logical_Operator_out6132_out1            : std_logic;
  SIGNAL Logical_Operator_out6133_out1            : std_logic;
  SIGNAL Logical_Operator_out6134_out1            : std_logic;
  SIGNAL Logical_Operator_out6135_out1            : std_logic;
  SIGNAL Logical_Operator_out6136_out1            : std_logic;
  SIGNAL Logical_Operator_out6137_out1            : std_logic;
  SIGNAL Logical_Operator_out6138_out1            : std_logic;
  SIGNAL Logical_Operator_out6139_out1            : std_logic;
  SIGNAL Logical_Operator_out6140_out1            : std_logic;
  SIGNAL Logical_Operator_out6141_out1            : std_logic;
  SIGNAL Logical_Operator_out6142_out1            : std_logic;
  SIGNAL Logical_Operator_out6143_out1            : std_logic;
  SIGNAL Logical_Operator_out6144_out1            : std_logic;
  SIGNAL Logical_Operator_out6145_out1            : std_logic;
  SIGNAL Logical_Operator_out6146_out1            : std_logic;
  SIGNAL Logical_Operator_out6147_out1            : std_logic;
  SIGNAL Logical_Operator_out6148_out1            : std_logic;
  SIGNAL Logical_Operator_out6149_out1            : std_logic;
  SIGNAL Logical_Operator_out6150_out1            : std_logic;
  SIGNAL Logical_Operator_out6151_out1            : std_logic;
  SIGNAL Logical_Operator_out6152_out1            : std_logic;
  SIGNAL Logical_Operator_out6153_out1            : std_logic;
  SIGNAL Logical_Operator_out6154_out1            : std_logic;
  SIGNAL Logical_Operator_out6155_out1            : std_logic;
  SIGNAL Logical_Operator_out6156_out1            : std_logic;
  SIGNAL Logical_Operator_out6157_out1            : std_logic;
  SIGNAL Logical_Operator_out6158_out1            : std_logic;
  SIGNAL Logical_Operator_out6159_out1            : std_logic;
  SIGNAL Logical_Operator_out6160_out1            : std_logic;
  SIGNAL Logical_Operator_out6161_out1            : std_logic;
  SIGNAL Logical_Operator_out6162_out1            : std_logic;
  SIGNAL Logical_Operator_out6163_out1            : std_logic;
  SIGNAL Logical_Operator_out6164_out1            : std_logic;
  SIGNAL Logical_Operator_out6165_out1            : std_logic;
  SIGNAL Logical_Operator_out6166_out1            : std_logic;
  SIGNAL Logical_Operator_out6167_out1            : std_logic;
  SIGNAL Logical_Operator_out6168_out1            : std_logic;
  SIGNAL Logical_Operator_out6169_out1            : std_logic;
  SIGNAL Logical_Operator_out6170_out1            : std_logic;
  SIGNAL Logical_Operator_out6171_out1            : std_logic;
  SIGNAL Logical_Operator_out6172_out1            : std_logic;
  SIGNAL Logical_Operator_out6173_out1            : std_logic;
  SIGNAL Logical_Operator_out6174_out1            : std_logic;
  SIGNAL Logical_Operator_out6175_out1            : std_logic;
  SIGNAL Logical_Operator_out6176_out1            : std_logic;
  SIGNAL Logical_Operator_out6177_out1            : std_logic;
  SIGNAL Logical_Operator_out6178_out1            : std_logic;
  SIGNAL Logical_Operator_out6179_out1            : std_logic;
  SIGNAL Logical_Operator_out6180_out1            : std_logic;
  SIGNAL Logical_Operator_out6181_out1            : std_logic;
  SIGNAL Logical_Operator_out6182_out1            : std_logic;
  SIGNAL Logical_Operator_out6183_out1            : std_logic;
  SIGNAL Logical_Operator_out6184_out1            : std_logic;
  SIGNAL Logical_Operator_out6185_out1            : std_logic;
  SIGNAL Logical_Operator_out6186_out1            : std_logic;
  SIGNAL Logical_Operator_out6187_out1            : std_logic;
  SIGNAL Logical_Operator_out6188_out1            : std_logic;
  SIGNAL Logical_Operator_out6189_out1            : std_logic;
  SIGNAL Logical_Operator_out6190_out1            : std_logic;
  SIGNAL Logical_Operator_out6191_out1            : std_logic;
  SIGNAL Logical_Operator_out6192_out1            : std_logic;
  SIGNAL Logical_Operator_out6193_out1            : std_logic;
  SIGNAL Logical_Operator_out6194_out1            : std_logic;
  SIGNAL Logical_Operator_out6195_out1            : std_logic;
  SIGNAL Logical_Operator_out6196_out1            : std_logic;
  SIGNAL Logical_Operator_out6197_out1            : std_logic;
  SIGNAL Logical_Operator_out6198_out1            : std_logic;
  SIGNAL Logical_Operator_out6199_out1            : std_logic;
  SIGNAL Logical_Operator_out6200_out1            : std_logic;
  SIGNAL Logical_Operator_out6201_out1            : std_logic;
  SIGNAL Logical_Operator_out6202_out1            : std_logic;
  SIGNAL Logical_Operator_out6203_out1            : std_logic;
  SIGNAL Logical_Operator_out6204_out1            : std_logic;
  SIGNAL Logical_Operator_out6205_out1            : std_logic;
  SIGNAL Logical_Operator_out6206_out1            : std_logic;
  SIGNAL Logical_Operator_out6207_out1            : std_logic;
  SIGNAL Logical_Operator_out6208_out1            : std_logic;
  SIGNAL Logical_Operator_out6209_out1            : std_logic;
  SIGNAL Logical_Operator_out6210_out1            : std_logic;
  SIGNAL Logical_Operator_out6211_out1            : std_logic;
  SIGNAL Logical_Operator_out6212_out1            : std_logic;
  SIGNAL Logical_Operator_out6213_out1            : std_logic;
  SIGNAL Logical_Operator_out6214_out1            : std_logic;
  SIGNAL Logical_Operator_out6215_out1            : std_logic;
  SIGNAL Logical_Operator_out6216_out1            : std_logic;
  SIGNAL Logical_Operator_out6217_out1            : std_logic;
  SIGNAL Logical_Operator_out6218_out1            : std_logic;
  SIGNAL Logical_Operator_out6219_out1            : std_logic;
  SIGNAL Logical_Operator_out6220_out1            : std_logic;
  SIGNAL Logical_Operator_out6221_out1            : std_logic;
  SIGNAL Logical_Operator_out6222_out1            : std_logic;
  SIGNAL Logical_Operator_out6223_out1            : std_logic;
  SIGNAL Logical_Operator_out6224_out1            : std_logic;
  SIGNAL Logical_Operator_out6225_out1            : std_logic;
  SIGNAL Logical_Operator_out6226_out1            : std_logic;
  SIGNAL Logical_Operator_out6227_out1            : std_logic;
  SIGNAL Logical_Operator_out6228_out1            : std_logic;
  SIGNAL Logical_Operator_out6229_out1            : std_logic;
  SIGNAL Logical_Operator_out6230_out1            : std_logic;
  SIGNAL Logical_Operator_out6231_out1            : std_logic;
  SIGNAL Logical_Operator_out6232_out1            : std_logic;
  SIGNAL Logical_Operator_out6233_out1            : std_logic;
  SIGNAL Logical_Operator_out6234_out1            : std_logic;
  SIGNAL Logical_Operator_out6235_out1            : std_logic;
  SIGNAL Logical_Operator_out6236_out1            : std_logic;
  SIGNAL Logical_Operator_out6237_out1            : std_logic;
  SIGNAL Logical_Operator_out6238_out1            : std_logic;
  SIGNAL Logical_Operator_out6239_out1            : std_logic;
  SIGNAL Logical_Operator_out6240_out1            : std_logic;
  SIGNAL Logical_Operator_out6241_out1            : std_logic;
  SIGNAL Logical_Operator_out6242_out1            : std_logic;
  SIGNAL Logical_Operator_out6243_out1            : std_logic;
  SIGNAL Logical_Operator_out6244_out1            : std_logic;
  SIGNAL Logical_Operator_out6245_out1            : std_logic;
  SIGNAL Logical_Operator_out6246_out1            : std_logic;
  SIGNAL Logical_Operator_out6247_out1            : std_logic;
  SIGNAL Logical_Operator_out6248_out1            : std_logic;
  SIGNAL Logical_Operator_out6249_out1            : std_logic;
  SIGNAL Logical_Operator_out6250_out1            : std_logic;
  SIGNAL Logical_Operator_out6251_out1            : std_logic;
  SIGNAL Logical_Operator_out6252_out1            : std_logic;
  SIGNAL Logical_Operator_out6253_out1            : std_logic;
  SIGNAL Logical_Operator_out6254_out1            : std_logic;
  SIGNAL Logical_Operator_out6255_out1            : std_logic;
  SIGNAL Logical_Operator_out6256_out1            : std_logic;
  SIGNAL Logical_Operator_out6257_out1            : std_logic;
  SIGNAL Logical_Operator_out6258_out1            : std_logic;
  SIGNAL Logical_Operator_out6259_out1            : std_logic;
  SIGNAL Logical_Operator_out6260_out1            : std_logic;
  SIGNAL Logical_Operator_out6261_out1            : std_logic;
  SIGNAL Logical_Operator_out6262_out1            : std_logic;
  SIGNAL Logical_Operator_out6263_out1            : std_logic;
  SIGNAL Logical_Operator_out6264_out1            : std_logic;
  SIGNAL Logical_Operator_out6265_out1            : std_logic;
  SIGNAL Logical_Operator_out6266_out1            : std_logic;
  SIGNAL Logical_Operator_out6267_out1            : std_logic;
  SIGNAL Logical_Operator_out6268_out1            : std_logic;
  SIGNAL Logical_Operator_out6269_out1            : std_logic;
  SIGNAL Logical_Operator_out6270_out1            : std_logic;
  SIGNAL Logical_Operator_out6271_out1            : std_logic;
  SIGNAL Logical_Operator_out6272_out1            : std_logic;
  SIGNAL Logical_Operator_out6273_out1            : std_logic;
  SIGNAL Logical_Operator_out6274_out1            : std_logic;
  SIGNAL Logical_Operator_out6275_out1            : std_logic;
  SIGNAL Logical_Operator_out6276_out1            : std_logic;
  SIGNAL Logical_Operator_out6277_out1            : std_logic;
  SIGNAL Logical_Operator_out6278_out1            : std_logic;
  SIGNAL Logical_Operator_out6279_out1            : std_logic;
  SIGNAL Logical_Operator_out6280_out1            : std_logic;
  SIGNAL Logical_Operator_out6281_out1            : std_logic;
  SIGNAL Logical_Operator_out6282_out1            : std_logic;
  SIGNAL Logical_Operator_out6283_out1            : std_logic;
  SIGNAL Logical_Operator_out6284_out1            : std_logic;
  SIGNAL Logical_Operator_out6285_out1            : std_logic;
  SIGNAL Logical_Operator_out6286_out1            : std_logic;
  SIGNAL Logical_Operator_out6287_out1            : std_logic;
  SIGNAL Logical_Operator_out6288_out1            : std_logic;
  SIGNAL Logical_Operator_out6289_out1            : std_logic;
  SIGNAL Logical_Operator_out6290_out1            : std_logic;
  SIGNAL Logical_Operator_out6291_out1            : std_logic;
  SIGNAL Logical_Operator_out6292_out1            : std_logic;
  SIGNAL Logical_Operator_out6293_out1            : std_logic;
  SIGNAL Logical_Operator_out6294_out1            : std_logic;
  SIGNAL Logical_Operator_out6295_out1            : std_logic;
  SIGNAL Logical_Operator_out6296_out1            : std_logic;
  SIGNAL Logical_Operator_out6297_out1            : std_logic;
  SIGNAL Logical_Operator_out6298_out1            : std_logic;
  SIGNAL Logical_Operator_out6299_out1            : std_logic;
  SIGNAL Logical_Operator_out6300_out1            : std_logic;
  SIGNAL Logical_Operator_out6301_out1            : std_logic;
  SIGNAL Logical_Operator_out6302_out1            : std_logic;
  SIGNAL Logical_Operator_out6303_out1            : std_logic;
  SIGNAL Logical_Operator_out6304_out1            : std_logic;
  SIGNAL Logical_Operator_out6305_out1            : std_logic;
  SIGNAL Logical_Operator_out6306_out1            : std_logic;
  SIGNAL Logical_Operator_out6307_out1            : std_logic;
  SIGNAL Logical_Operator_out6308_out1            : std_logic;
  SIGNAL Logical_Operator_out6309_out1            : std_logic;
  SIGNAL Logical_Operator_out6310_out1            : std_logic;
  SIGNAL Logical_Operator_out6311_out1            : std_logic;
  SIGNAL Logical_Operator_out6312_out1            : std_logic;
  SIGNAL Logical_Operator_out6313_out1            : std_logic;
  SIGNAL Logical_Operator_out6314_out1            : std_logic;
  SIGNAL Logical_Operator_out6315_out1            : std_logic;
  SIGNAL Logical_Operator_out6316_out1            : std_logic;
  SIGNAL Logical_Operator_out6317_out1            : std_logic;
  SIGNAL Logical_Operator_out6318_out1            : std_logic;
  SIGNAL Logical_Operator_out6319_out1            : std_logic;
  SIGNAL Logical_Operator_out6320_out1            : std_logic;
  SIGNAL Logical_Operator_out6321_out1            : std_logic;
  SIGNAL Logical_Operator_out6322_out1            : std_logic;
  SIGNAL Logical_Operator_out6323_out1            : std_logic;
  SIGNAL Logical_Operator_out6324_out1            : std_logic;
  SIGNAL Logical_Operator_out6325_out1            : std_logic;
  SIGNAL Logical_Operator_out6326_out1            : std_logic;
  SIGNAL Logical_Operator_out6327_out1            : std_logic;
  SIGNAL Logical_Operator_out6328_out1            : std_logic;
  SIGNAL Logical_Operator_out6329_out1            : std_logic;
  SIGNAL Logical_Operator_out6330_out1            : std_logic;
  SIGNAL Logical_Operator_out6331_out1            : std_logic;
  SIGNAL Logical_Operator_out6332_out1            : std_logic;
  SIGNAL Logical_Operator_out6333_out1            : std_logic;
  SIGNAL Logical_Operator_out6334_out1            : std_logic;
  SIGNAL Logical_Operator_out6335_out1            : std_logic;
  SIGNAL Logical_Operator_out6336_out1            : std_logic;
  SIGNAL Logical_Operator_out6337_out1            : std_logic;
  SIGNAL Logical_Operator_out6338_out1            : std_logic;
  SIGNAL Logical_Operator_out6339_out1            : std_logic;
  SIGNAL Logical_Operator_out6340_out1            : std_logic;
  SIGNAL Logical_Operator_out6341_out1            : std_logic;
  SIGNAL Logical_Operator_out6342_out1            : std_logic;
  SIGNAL Logical_Operator_out6343_out1            : std_logic;
  SIGNAL Logical_Operator_out6344_out1            : std_logic;
  SIGNAL Logical_Operator_out6345_out1            : std_logic;
  SIGNAL Logical_Operator_out6346_out1            : std_logic;
  SIGNAL Logical_Operator_out6347_out1            : std_logic;
  SIGNAL Logical_Operator_out6348_out1            : std_logic;
  SIGNAL Logical_Operator_out6349_out1            : std_logic;
  SIGNAL Logical_Operator_out6350_out1            : std_logic;
  SIGNAL Logical_Operator_out6351_out1            : std_logic;
  SIGNAL Logical_Operator_out6352_out1            : std_logic;
  SIGNAL Logical_Operator_out6353_out1            : std_logic;
  SIGNAL Logical_Operator_out6354_out1            : std_logic;
  SIGNAL Logical_Operator_out6355_out1            : std_logic;
  SIGNAL Logical_Operator_out6356_out1            : std_logic;
  SIGNAL Logical_Operator_out6357_out1            : std_logic;
  SIGNAL Logical_Operator_out6358_out1            : std_logic;
  SIGNAL Logical_Operator_out6359_out1            : std_logic;
  SIGNAL Logical_Operator_out6360_out1            : std_logic;
  SIGNAL Logical_Operator_out6361_out1            : std_logic;
  SIGNAL Logical_Operator_out6362_out1            : std_logic;
  SIGNAL Logical_Operator_out6363_out1            : std_logic;
  SIGNAL Logical_Operator_out6364_out1            : std_logic;
  SIGNAL Logical_Operator_out6365_out1            : std_logic;
  SIGNAL Logical_Operator_out6366_out1            : std_logic;
  SIGNAL Logical_Operator_out6367_out1            : std_logic;
  SIGNAL Logical_Operator_out6368_out1            : std_logic;
  SIGNAL Logical_Operator_out6369_out1            : std_logic;
  SIGNAL Logical_Operator_out6370_out1            : std_logic;
  SIGNAL Logical_Operator_out6371_out1            : std_logic;
  SIGNAL Logical_Operator_out6372_out1            : std_logic;
  SIGNAL Logical_Operator_out6373_out1            : std_logic;
  SIGNAL Logical_Operator_out6374_out1            : std_logic;
  SIGNAL Logical_Operator_out6375_out1            : std_logic;
  SIGNAL Logical_Operator_out6376_out1            : std_logic;
  SIGNAL Logical_Operator_out6377_out1            : std_logic;
  SIGNAL Logical_Operator_out6378_out1            : std_logic;
  SIGNAL Logical_Operator_out6379_out1            : std_logic;
  SIGNAL Logical_Operator_out6380_out1            : std_logic;
  SIGNAL Logical_Operator_out6381_out1            : std_logic;
  SIGNAL Logical_Operator_out6382_out1            : std_logic;
  SIGNAL Logical_Operator_out6383_out1            : std_logic;
  SIGNAL Logical_Operator_out6384_out1            : std_logic;
  SIGNAL Logical_Operator_out6385_out1            : std_logic;
  SIGNAL Logical_Operator_out6386_out1            : std_logic;
  SIGNAL Logical_Operator_out6387_out1            : std_logic;
  SIGNAL Logical_Operator_out6388_out1            : std_logic;
  SIGNAL Logical_Operator_out6389_out1            : std_logic;
  SIGNAL Logical_Operator_out6390_out1            : std_logic;
  SIGNAL Logical_Operator_out6391_out1            : std_logic;
  SIGNAL Logical_Operator_out6392_out1            : std_logic;
  SIGNAL Logical_Operator_out6393_out1            : std_logic;
  SIGNAL Logical_Operator_out6394_out1            : std_logic;
  SIGNAL Logical_Operator_out6395_out1            : std_logic;
  SIGNAL Logical_Operator_out6396_out1            : std_logic;
  SIGNAL Logical_Operator_out6397_out1            : std_logic;
  SIGNAL Logical_Operator_out6398_out1            : std_logic;
  SIGNAL Logical_Operator_out6399_out1            : std_logic;
  SIGNAL Logical_Operator_out6400_out1            : std_logic;
  SIGNAL Logical_Operator_out6401_out1            : std_logic;
  SIGNAL Logical_Operator_out6402_out1            : std_logic;
  SIGNAL Logical_Operator_out6403_out1            : std_logic;
  SIGNAL Logical_Operator_out6404_out1            : std_logic;
  SIGNAL Logical_Operator_out6405_out1            : std_logic;
  SIGNAL Logical_Operator_out6406_out1            : std_logic;
  SIGNAL Logical_Operator_out6407_out1            : std_logic;
  SIGNAL Logical_Operator_out6408_out1            : std_logic;
  SIGNAL Logical_Operator_out6409_out1            : std_logic;
  SIGNAL Logical_Operator_out6410_out1            : std_logic;
  SIGNAL Logical_Operator_out6411_out1            : std_logic;
  SIGNAL Logical_Operator_out6412_out1            : std_logic;
  SIGNAL Logical_Operator_out6413_out1            : std_logic;
  SIGNAL Logical_Operator_out6414_out1            : std_logic;
  SIGNAL Logical_Operator_out6415_out1            : std_logic;
  SIGNAL Logical_Operator_out6416_out1            : std_logic;
  SIGNAL Logical_Operator_out6417_out1            : std_logic;
  SIGNAL Logical_Operator_out6418_out1            : std_logic;
  SIGNAL Logical_Operator_out6419_out1            : std_logic;
  SIGNAL Logical_Operator_out6420_out1            : std_logic;
  SIGNAL Logical_Operator_out6421_out1            : std_logic;
  SIGNAL Logical_Operator_out6422_out1            : std_logic;
  SIGNAL Logical_Operator_out6423_out1            : std_logic;
  SIGNAL Logical_Operator_out6424_out1            : std_logic;
  SIGNAL Logical_Operator_out6425_out1            : std_logic;
  SIGNAL Logical_Operator_out6426_out1            : std_logic;
  SIGNAL Logical_Operator_out6427_out1            : std_logic;
  SIGNAL Logical_Operator_out6428_out1            : std_logic;
  SIGNAL Logical_Operator_out6429_out1            : std_logic;
  SIGNAL Logical_Operator_out6430_out1            : std_logic;
  SIGNAL Logical_Operator_out6431_out1            : std_logic;
  SIGNAL Logical_Operator_out6432_out1            : std_logic;
  SIGNAL Logical_Operator_out6433_out1            : std_logic;
  SIGNAL Logical_Operator_out6434_out1            : std_logic;
  SIGNAL Logical_Operator_out6435_out1            : std_logic;
  SIGNAL Logical_Operator_out6436_out1            : std_logic;
  SIGNAL Logical_Operator_out6437_out1            : std_logic;
  SIGNAL Logical_Operator_out6438_out1            : std_logic;
  SIGNAL Logical_Operator_out6439_out1            : std_logic;
  SIGNAL Logical_Operator_out6440_out1            : std_logic;
  SIGNAL Logical_Operator_out6441_out1            : std_logic;
  SIGNAL Logical_Operator_out6442_out1            : std_logic;
  SIGNAL Logical_Operator_out6443_out1            : std_logic;
  SIGNAL Logical_Operator_out6444_out1            : std_logic;
  SIGNAL Logical_Operator_out6445_out1            : std_logic;
  SIGNAL Logical_Operator_out6446_out1            : std_logic;
  SIGNAL Logical_Operator_out6447_out1            : std_logic;
  SIGNAL Logical_Operator_out6448_out1            : std_logic;
  SIGNAL Logical_Operator_out6449_out1            : std_logic;
  SIGNAL Logical_Operator_out6450_out1            : std_logic;
  SIGNAL Logical_Operator_out6451_out1            : std_logic;
  SIGNAL Logical_Operator_out6452_out1            : std_logic;
  SIGNAL Logical_Operator_out6453_out1            : std_logic;
  SIGNAL Logical_Operator_out6454_out1            : std_logic;
  SIGNAL Logical_Operator_out6455_out1            : std_logic;
  SIGNAL Logical_Operator_out6456_out1            : std_logic;
  SIGNAL Logical_Operator_out6457_out1            : std_logic;
  SIGNAL Logical_Operator_out6458_out1            : std_logic;
  SIGNAL Logical_Operator_out6459_out1            : std_logic;
  SIGNAL Logical_Operator_out6460_out1            : std_logic;
  SIGNAL Logical_Operator_out6461_out1            : std_logic;
  SIGNAL Logical_Operator_out6462_out1            : std_logic;
  SIGNAL Logical_Operator_out6463_out1            : std_logic;
  SIGNAL Logical_Operator_out6464_out1            : std_logic;
  SIGNAL Logical_Operator_out6465_out1            : std_logic;
  SIGNAL Logical_Operator_out6466_out1            : std_logic;
  SIGNAL Logical_Operator_out6467_out1            : std_logic;
  SIGNAL Logical_Operator_out6468_out1            : std_logic;
  SIGNAL Logical_Operator_out6469_out1            : std_logic;
  SIGNAL Logical_Operator_out6470_out1            : std_logic;
  SIGNAL Logical_Operator_out6471_out1            : std_logic;
  SIGNAL Logical_Operator_out6472_out1            : std_logic;
  SIGNAL Logical_Operator_out6473_out1            : std_logic;
  SIGNAL Logical_Operator_out6474_out1            : std_logic;
  SIGNAL Logical_Operator_out6475_out1            : std_logic;
  SIGNAL Logical_Operator_out6476_out1            : std_logic;
  SIGNAL Logical_Operator_out6477_out1            : std_logic;
  SIGNAL Logical_Operator_out6478_out1            : std_logic;
  SIGNAL Logical_Operator_out6479_out1            : std_logic;
  SIGNAL Logical_Operator_out6480_out1            : std_logic;
  SIGNAL Logical_Operator_out6481_out1            : std_logic;
  SIGNAL Logical_Operator_out6482_out1            : std_logic;
  SIGNAL Logical_Operator_out6483_out1            : std_logic;
  SIGNAL Logical_Operator_out6484_out1            : std_logic;
  SIGNAL Logical_Operator_out6485_out1            : std_logic;
  SIGNAL Logical_Operator_out6486_out1            : std_logic;
  SIGNAL Logical_Operator_out6487_out1            : std_logic;
  SIGNAL Logical_Operator_out6488_out1            : std_logic;
  SIGNAL Logical_Operator_out6489_out1            : std_logic;
  SIGNAL Logical_Operator_out6490_out1            : std_logic;
  SIGNAL Logical_Operator_out6491_out1            : std_logic;
  SIGNAL Logical_Operator_out6492_out1            : std_logic;
  SIGNAL Logical_Operator_out6493_out1            : std_logic;
  SIGNAL Logical_Operator_out6494_out1            : std_logic;
  SIGNAL Logical_Operator_out6495_out1            : std_logic;
  SIGNAL Logical_Operator_out6496_out1            : std_logic;
  SIGNAL Logical_Operator_out6497_out1            : std_logic;
  SIGNAL Logical_Operator_out6498_out1            : std_logic;
  SIGNAL Logical_Operator_out6499_out1            : std_logic;
  SIGNAL Logical_Operator_out6500_out1            : std_logic;
  SIGNAL Logical_Operator_out6501_out1            : std_logic;
  SIGNAL Logical_Operator_out6502_out1            : std_logic;
  SIGNAL Logical_Operator_out6503_out1            : std_logic;
  SIGNAL Logical_Operator_out6504_out1            : std_logic;
  SIGNAL Logical_Operator_out6505_out1            : std_logic;
  SIGNAL Logical_Operator_out6506_out1            : std_logic;
  SIGNAL Logical_Operator_out6507_out1            : std_logic;
  SIGNAL Logical_Operator_out6508_out1            : std_logic;
  SIGNAL Logical_Operator_out6509_out1            : std_logic;
  SIGNAL Logical_Operator_out6510_out1            : std_logic;
  SIGNAL Logical_Operator_out6511_out1            : std_logic;
  SIGNAL Logical_Operator_out6512_out1            : std_logic;
  SIGNAL Logical_Operator_out6513_out1            : std_logic;
  SIGNAL Logical_Operator_out6514_out1            : std_logic;
  SIGNAL Logical_Operator_out6515_out1            : std_logic;
  SIGNAL Logical_Operator_out6516_out1            : std_logic;
  SIGNAL Logical_Operator_out6517_out1            : std_logic;
  SIGNAL Logical_Operator_out6518_out1            : std_logic;
  SIGNAL Logical_Operator_out6519_out1            : std_logic;
  SIGNAL Logical_Operator_out6520_out1            : std_logic;
  SIGNAL Logical_Operator_out6521_out1            : std_logic;
  SIGNAL Logical_Operator_out6522_out1            : std_logic;
  SIGNAL Logical_Operator_out6523_out1            : std_logic;
  SIGNAL Logical_Operator_out6524_out1            : std_logic;
  SIGNAL Logical_Operator_out6525_out1            : std_logic;
  SIGNAL Logical_Operator_out6526_out1            : std_logic;
  SIGNAL Logical_Operator_out6527_out1            : std_logic;
  SIGNAL Logical_Operator_out6528_out1            : std_logic;
  SIGNAL Logical_Operator_out6529_out1            : std_logic;
  SIGNAL Logical_Operator_out6530_out1            : std_logic;
  SIGNAL Logical_Operator_out6531_out1            : std_logic;
  SIGNAL Logical_Operator_out6532_out1            : std_logic;
  SIGNAL Logical_Operator_out6533_out1            : std_logic;
  SIGNAL Logical_Operator_out6534_out1            : std_logic;
  SIGNAL Logical_Operator_out6535_out1            : std_logic;
  SIGNAL Logical_Operator_out6536_out1            : std_logic;
  SIGNAL Logical_Operator_out6537_out1            : std_logic;
  SIGNAL Logical_Operator_out6538_out1            : std_logic;
  SIGNAL Logical_Operator_out6539_out1            : std_logic;
  SIGNAL Logical_Operator_out6540_out1            : std_logic;
  SIGNAL Logical_Operator_out6541_out1            : std_logic;
  SIGNAL Logical_Operator_out6542_out1            : std_logic;
  SIGNAL Logical_Operator_out6543_out1            : std_logic;
  SIGNAL Logical_Operator_out6544_out1            : std_logic;
  SIGNAL Logical_Operator_out6545_out1            : std_logic;
  SIGNAL Logical_Operator_out6546_out1            : std_logic;
  SIGNAL Logical_Operator_out6547_out1            : std_logic;
  SIGNAL Logical_Operator_out6548_out1            : std_logic;
  SIGNAL Logical_Operator_out6549_out1            : std_logic;
  SIGNAL Logical_Operator_out6550_out1            : std_logic;
  SIGNAL Logical_Operator_out6551_out1            : std_logic;
  SIGNAL Logical_Operator_out6552_out1            : std_logic;
  SIGNAL Logical_Operator_out6553_out1            : std_logic;
  SIGNAL Logical_Operator_out6554_out1            : std_logic;
  SIGNAL Logical_Operator_out6555_out1            : std_logic;
  SIGNAL Logical_Operator_out6556_out1            : std_logic;
  SIGNAL Logical_Operator_out6557_out1            : std_logic;
  SIGNAL Logical_Operator_out6558_out1            : std_logic;
  SIGNAL Logical_Operator_out6559_out1            : std_logic;
  SIGNAL Logical_Operator_out6560_out1            : std_logic;
  SIGNAL Logical_Operator_out6561_out1            : std_logic;
  SIGNAL Logical_Operator_out6562_out1            : std_logic;
  SIGNAL Logical_Operator_out6563_out1            : std_logic;
  SIGNAL Logical_Operator_out6564_out1            : std_logic;
  SIGNAL Logical_Operator_out6565_out1            : std_logic;
  SIGNAL Logical_Operator_out6566_out1            : std_logic;
  SIGNAL Logical_Operator_out6567_out1            : std_logic;
  SIGNAL Logical_Operator_out6568_out1            : std_logic;
  SIGNAL Logical_Operator_out6569_out1            : std_logic;
  SIGNAL Logical_Operator_out6570_out1            : std_logic;
  SIGNAL Logical_Operator_out6571_out1            : std_logic;
  SIGNAL Logical_Operator_out6572_out1            : std_logic;
  SIGNAL Logical_Operator_out6573_out1            : std_logic;
  SIGNAL Logical_Operator_out6574_out1            : std_logic;
  SIGNAL Logical_Operator_out6575_out1            : std_logic;
  SIGNAL Logical_Operator_out6576_out1            : std_logic;
  SIGNAL Logical_Operator_out6577_out1            : std_logic;
  SIGNAL Logical_Operator_out6578_out1            : std_logic;
  SIGNAL Logical_Operator_out6579_out1            : std_logic;
  SIGNAL Logical_Operator_out6580_out1            : std_logic;
  SIGNAL Logical_Operator_out6581_out1            : std_logic;
  SIGNAL Logical_Operator_out6582_out1            : std_logic;
  SIGNAL Logical_Operator_out6583_out1            : std_logic;
  SIGNAL Logical_Operator_out6584_out1            : std_logic;
  SIGNAL Logical_Operator_out6585_out1            : std_logic;
  SIGNAL Logical_Operator_out6586_out1            : std_logic;
  SIGNAL Logical_Operator_out6587_out1            : std_logic;
  SIGNAL Logical_Operator_out6588_out1            : std_logic;
  SIGNAL Logical_Operator_out6589_out1            : std_logic;
  SIGNAL Logical_Operator_out6590_out1            : std_logic;
  SIGNAL Logical_Operator_out6591_out1            : std_logic;
  SIGNAL Logical_Operator_out6592_out1            : std_logic;
  SIGNAL Logical_Operator_out6593_out1            : std_logic;
  SIGNAL Logical_Operator_out6594_out1            : std_logic;
  SIGNAL Logical_Operator_out6595_out1            : std_logic;
  SIGNAL Logical_Operator_out6596_out1            : std_logic;
  SIGNAL Logical_Operator_out6597_out1            : std_logic;
  SIGNAL Logical_Operator_out6598_out1            : std_logic;
  SIGNAL Logical_Operator_out6599_out1            : std_logic;
  SIGNAL Logical_Operator_out6600_out1            : std_logic;
  SIGNAL Logical_Operator_out6601_out1            : std_logic;
  SIGNAL Logical_Operator_out6602_out1            : std_logic;
  SIGNAL Logical_Operator_out6603_out1            : std_logic;
  SIGNAL Logical_Operator_out6604_out1            : std_logic;
  SIGNAL Logical_Operator_out6605_out1            : std_logic;
  SIGNAL Logical_Operator_out6606_out1            : std_logic;
  SIGNAL Logical_Operator_out6607_out1            : std_logic;
  SIGNAL Logical_Operator_out6608_out1            : std_logic;
  SIGNAL Logical_Operator_out6609_out1            : std_logic;
  SIGNAL Logical_Operator_out6610_out1            : std_logic;
  SIGNAL Logical_Operator_out6611_out1            : std_logic;
  SIGNAL Logical_Operator_out6612_out1            : std_logic;
  SIGNAL Logical_Operator_out6613_out1            : std_logic;
  SIGNAL Logical_Operator_out6614_out1            : std_logic;
  SIGNAL Logical_Operator_out6615_out1            : std_logic;
  SIGNAL Logical_Operator_out6616_out1            : std_logic;
  SIGNAL Logical_Operator_out6617_out1            : std_logic;
  SIGNAL Logical_Operator_out6618_out1            : std_logic;
  SIGNAL Logical_Operator_out6619_out1            : std_logic;
  SIGNAL Logical_Operator_out6620_out1            : std_logic;
  SIGNAL Logical_Operator_out6621_out1            : std_logic;
  SIGNAL Logical_Operator_out6622_out1            : std_logic;
  SIGNAL Logical_Operator_out6623_out1            : std_logic;
  SIGNAL Logical_Operator_out6624_out1            : std_logic;
  SIGNAL Logical_Operator_out6625_out1            : std_logic;
  SIGNAL Logical_Operator_out6626_out1            : std_logic;
  SIGNAL Logical_Operator_out6627_out1            : std_logic;
  SIGNAL Logical_Operator_out6628_out1            : std_logic;
  SIGNAL Logical_Operator_out6629_out1            : std_logic;
  SIGNAL Logical_Operator_out6630_out1            : std_logic;
  SIGNAL Logical_Operator_out6631_out1            : std_logic;
  SIGNAL Logical_Operator_out6632_out1            : std_logic;
  SIGNAL Logical_Operator_out6633_out1            : std_logic;
  SIGNAL Logical_Operator_out6634_out1            : std_logic;
  SIGNAL Logical_Operator_out6635_out1            : std_logic;
  SIGNAL Logical_Operator_out6636_out1            : std_logic;
  SIGNAL Logical_Operator_out6637_out1            : std_logic;
  SIGNAL Logical_Operator_out6638_out1            : std_logic;
  SIGNAL Logical_Operator_out6639_out1            : std_logic;
  SIGNAL Logical_Operator_out6640_out1            : std_logic;
  SIGNAL Logical_Operator_out6641_out1            : std_logic;
  SIGNAL Logical_Operator_out6642_out1            : std_logic;
  SIGNAL Logical_Operator_out6643_out1            : std_logic;
  SIGNAL Logical_Operator_out6644_out1            : std_logic;
  SIGNAL Logical_Operator_out6645_out1            : std_logic;
  SIGNAL Logical_Operator_out6646_out1            : std_logic;
  SIGNAL Logical_Operator_out6647_out1            : std_logic;
  SIGNAL Logical_Operator_out6648_out1            : std_logic;
  SIGNAL Logical_Operator_out6649_out1            : std_logic;
  SIGNAL Logical_Operator_out6650_out1            : std_logic;
  SIGNAL Logical_Operator_out6651_out1            : std_logic;
  SIGNAL Logical_Operator_out6652_out1            : std_logic;
  SIGNAL Logical_Operator_out6653_out1            : std_logic;
  SIGNAL Logical_Operator_out6654_out1            : std_logic;
  SIGNAL Logical_Operator_out6655_out1            : std_logic;
  SIGNAL Logical_Operator_out6656_out1            : std_logic;
  SIGNAL Logical_Operator_out6657_out1            : std_logic;
  SIGNAL Logical_Operator_out6658_out1            : std_logic;
  SIGNAL Logical_Operator_out6659_out1            : std_logic;
  SIGNAL Logical_Operator_out6660_out1            : std_logic;
  SIGNAL Logical_Operator_out6661_out1            : std_logic;
  SIGNAL Logical_Operator_out6662_out1            : std_logic;
  SIGNAL Logical_Operator_out6663_out1            : std_logic;
  SIGNAL Logical_Operator_out6664_out1            : std_logic;
  SIGNAL Logical_Operator_out6665_out1            : std_logic;
  SIGNAL Logical_Operator_out6666_out1            : std_logic;
  SIGNAL Logical_Operator_out6667_out1            : std_logic;
  SIGNAL Logical_Operator_out6668_out1            : std_logic;
  SIGNAL Logical_Operator_out6669_out1            : std_logic;
  SIGNAL Logical_Operator_out6670_out1            : std_logic;
  SIGNAL Logical_Operator_out6671_out1            : std_logic;
  SIGNAL Logical_Operator_out6672_out1            : std_logic;
  SIGNAL Logical_Operator_out6673_out1            : std_logic;
  SIGNAL Logical_Operator_out6674_out1            : std_logic;
  SIGNAL Logical_Operator_out6675_out1            : std_logic;
  SIGNAL Logical_Operator_out6676_out1            : std_logic;
  SIGNAL Logical_Operator_out6677_out1            : std_logic;
  SIGNAL Logical_Operator_out6678_out1            : std_logic;
  SIGNAL Logical_Operator_out6679_out1            : std_logic;
  SIGNAL Logical_Operator_out6680_out1            : std_logic;
  SIGNAL Logical_Operator_out6681_out1            : std_logic;
  SIGNAL Logical_Operator_out6682_out1            : std_logic;
  SIGNAL Logical_Operator_out6683_out1            : std_logic;
  SIGNAL Logical_Operator_out6684_out1            : std_logic;
  SIGNAL Logical_Operator_out6685_out1            : std_logic;
  SIGNAL Logical_Operator_out6686_out1            : std_logic;
  SIGNAL Logical_Operator_out6687_out1            : std_logic;
  SIGNAL Logical_Operator_out6688_out1            : std_logic;
  SIGNAL Logical_Operator_out6689_out1            : std_logic;
  SIGNAL Logical_Operator_out6690_out1            : std_logic;
  SIGNAL Logical_Operator_out6691_out1            : std_logic;
  SIGNAL Logical_Operator_out6692_out1            : std_logic;
  SIGNAL Logical_Operator_out6693_out1            : std_logic;
  SIGNAL Logical_Operator_out6694_out1            : std_logic;
  SIGNAL Logical_Operator_out6695_out1            : std_logic;
  SIGNAL Logical_Operator_out6696_out1            : std_logic;
  SIGNAL Logical_Operator_out6697_out1            : std_logic;
  SIGNAL Logical_Operator_out6698_out1            : std_logic;
  SIGNAL Logical_Operator_out6699_out1            : std_logic;
  SIGNAL Logical_Operator_out6700_out1            : std_logic;
  SIGNAL Logical_Operator_out6701_out1            : std_logic;
  SIGNAL Logical_Operator_out6702_out1            : std_logic;
  SIGNAL Logical_Operator_out6703_out1            : std_logic;
  SIGNAL Logical_Operator_out6704_out1            : std_logic;
  SIGNAL Logical_Operator_out6705_out1            : std_logic;
  SIGNAL Logical_Operator_out6706_out1            : std_logic;
  SIGNAL Logical_Operator_out6707_out1            : std_logic;
  SIGNAL Logical_Operator_out6708_out1            : std_logic;
  SIGNAL Logical_Operator_out6709_out1            : std_logic;
  SIGNAL Logical_Operator_out6710_out1            : std_logic;
  SIGNAL Logical_Operator_out6711_out1            : std_logic;
  SIGNAL Logical_Operator_out6712_out1            : std_logic;
  SIGNAL Logical_Operator_out6713_out1            : std_logic;
  SIGNAL Logical_Operator_out6714_out1            : std_logic;
  SIGNAL Logical_Operator_out6715_out1            : std_logic;
  SIGNAL Logical_Operator_out6716_out1            : std_logic;
  SIGNAL Logical_Operator_out6717_out1            : std_logic;
  SIGNAL Logical_Operator_out6718_out1            : std_logic;
  SIGNAL Logical_Operator_out6719_out1            : std_logic;
  SIGNAL Logical_Operator_out6720_out1            : std_logic;
  SIGNAL Logical_Operator_out6721_out1            : std_logic;
  SIGNAL Logical_Operator_out6722_out1            : std_logic;
  SIGNAL Logical_Operator_out6723_out1            : std_logic;
  SIGNAL Logical_Operator_out6724_out1            : std_logic;
  SIGNAL Logical_Operator_out6725_out1            : std_logic;
  SIGNAL Logical_Operator_out6726_out1            : std_logic;
  SIGNAL Logical_Operator_out6727_out1            : std_logic;
  SIGNAL Logical_Operator_out6728_out1            : std_logic;
  SIGNAL Logical_Operator_out6729_out1            : std_logic;
  SIGNAL Logical_Operator_out6730_out1            : std_logic;
  SIGNAL Logical_Operator_out6731_out1            : std_logic;
  SIGNAL Logical_Operator_out6732_out1            : std_logic;
  SIGNAL Logical_Operator_out6733_out1            : std_logic;
  SIGNAL Logical_Operator_out6734_out1            : std_logic;
  SIGNAL Logical_Operator_out6735_out1            : std_logic;
  SIGNAL Logical_Operator_out6736_out1            : std_logic;
  SIGNAL Logical_Operator_out6737_out1            : std_logic;
  SIGNAL Logical_Operator_out6738_out1            : std_logic;
  SIGNAL Logical_Operator_out6739_out1            : std_logic;
  SIGNAL Logical_Operator_out6740_out1            : std_logic;
  SIGNAL Logical_Operator_out6741_out1            : std_logic;
  SIGNAL Logical_Operator_out6742_out1            : std_logic;
  SIGNAL Logical_Operator_out6743_out1            : std_logic;
  SIGNAL Logical_Operator_out6744_out1            : std_logic;
  SIGNAL Logical_Operator_out6745_out1            : std_logic;
  SIGNAL Logical_Operator_out6746_out1            : std_logic;
  SIGNAL Logical_Operator_out6747_out1            : std_logic;
  SIGNAL Logical_Operator_out6748_out1            : std_logic;
  SIGNAL Logical_Operator_out6749_out1            : std_logic;
  SIGNAL Logical_Operator_out6750_out1            : std_logic;
  SIGNAL Logical_Operator_out6751_out1            : std_logic;
  SIGNAL Logical_Operator_out6752_out1            : std_logic;
  SIGNAL Logical_Operator_out6753_out1            : std_logic;
  SIGNAL Logical_Operator_out6754_out1            : std_logic;
  SIGNAL Logical_Operator_out6755_out1            : std_logic;
  SIGNAL Logical_Operator_out6756_out1            : std_logic;
  SIGNAL Logical_Operator_out6757_out1            : std_logic;
  SIGNAL Logical_Operator_out6758_out1            : std_logic;
  SIGNAL Logical_Operator_out6759_out1            : std_logic;
  SIGNAL Logical_Operator_out6760_out1            : std_logic;
  SIGNAL Logical_Operator_out6761_out1            : std_logic;
  SIGNAL Logical_Operator_out6762_out1            : std_logic;
  SIGNAL Logical_Operator_out6763_out1            : std_logic;
  SIGNAL Logical_Operator_out6764_out1            : std_logic;
  SIGNAL Logical_Operator_out6765_out1            : std_logic;
  SIGNAL Logical_Operator_out6766_out1            : std_logic;
  SIGNAL Logical_Operator_out6767_out1            : std_logic;
  SIGNAL Logical_Operator_out6768_out1            : std_logic;
  SIGNAL Logical_Operator_out6769_out1            : std_logic;
  SIGNAL Logical_Operator_out6770_out1            : std_logic;
  SIGNAL Logical_Operator_out6771_out1            : std_logic;
  SIGNAL Logical_Operator_out6772_out1            : std_logic;
  SIGNAL Logical_Operator_out6773_out1            : std_logic;
  SIGNAL Logical_Operator_out6774_out1            : std_logic;
  SIGNAL Logical_Operator_out6775_out1            : std_logic;
  SIGNAL Logical_Operator_out6776_out1            : std_logic;
  SIGNAL Logical_Operator_out6777_out1            : std_logic;
  SIGNAL Logical_Operator_out6778_out1            : std_logic;
  SIGNAL Logical_Operator_out6779_out1            : std_logic;
  SIGNAL Logical_Operator_out6780_out1            : std_logic;
  SIGNAL Logical_Operator_out6781_out1            : std_logic;
  SIGNAL Logical_Operator_out6782_out1            : std_logic;
  SIGNAL Logical_Operator_out6783_out1            : std_logic;
  SIGNAL Logical_Operator_out6784_out1            : std_logic;
  SIGNAL Logical_Operator_out6785_out1            : std_logic;
  SIGNAL Logical_Operator_out6786_out1            : std_logic;
  SIGNAL Logical_Operator_out6787_out1            : std_logic;
  SIGNAL Logical_Operator_out6788_out1            : std_logic;
  SIGNAL Logical_Operator_out6789_out1            : std_logic;
  SIGNAL Logical_Operator_out6790_out1            : std_logic;
  SIGNAL Logical_Operator_out6791_out1            : std_logic;
  SIGNAL Logical_Operator_out6792_out1            : std_logic;
  SIGNAL Logical_Operator_out6793_out1            : std_logic;
  SIGNAL Logical_Operator_out6794_out1            : std_logic;
  SIGNAL Logical_Operator_out6795_out1            : std_logic;
  SIGNAL Logical_Operator_out6796_out1            : std_logic;
  SIGNAL Logical_Operator_out6797_out1            : std_logic;
  SIGNAL Logical_Operator_out6798_out1            : std_logic;
  SIGNAL Logical_Operator_out6799_out1            : std_logic;
  SIGNAL Logical_Operator_out6800_out1            : std_logic;
  SIGNAL Logical_Operator_out6801_out1            : std_logic;
  SIGNAL Logical_Operator_out6802_out1            : std_logic;
  SIGNAL Logical_Operator_out6803_out1            : std_logic;
  SIGNAL Logical_Operator_out6804_out1            : std_logic;
  SIGNAL Logical_Operator_out6805_out1            : std_logic;
  SIGNAL Logical_Operator_out6806_out1            : std_logic;
  SIGNAL Logical_Operator_out6807_out1            : std_logic;
  SIGNAL Logical_Operator_out6808_out1            : std_logic;
  SIGNAL Logical_Operator_out6809_out1            : std_logic;
  SIGNAL Logical_Operator_out6810_out1            : std_logic;
  SIGNAL Logical_Operator_out6811_out1            : std_logic;
  SIGNAL Logical_Operator_out6812_out1            : std_logic;
  SIGNAL Logical_Operator_out6813_out1            : std_logic;
  SIGNAL Logical_Operator_out6814_out1            : std_logic;
  SIGNAL Logical_Operator_out6815_out1            : std_logic;
  SIGNAL Logical_Operator_out6816_out1            : std_logic;
  SIGNAL Logical_Operator_out6817_out1            : std_logic;
  SIGNAL Logical_Operator_out6818_out1            : std_logic;
  SIGNAL Logical_Operator_out6819_out1            : std_logic;
  SIGNAL Logical_Operator_out6820_out1            : std_logic;
  SIGNAL Logical_Operator_out6821_out1            : std_logic;
  SIGNAL Logical_Operator_out6822_out1            : std_logic;
  SIGNAL Logical_Operator_out6823_out1            : std_logic;
  SIGNAL Logical_Operator_out6824_out1            : std_logic;
  SIGNAL Logical_Operator_out6825_out1            : std_logic;
  SIGNAL Logical_Operator_out6826_out1            : std_logic;
  SIGNAL Logical_Operator_out6827_out1            : std_logic;
  SIGNAL Logical_Operator_out6828_out1            : std_logic;
  SIGNAL Logical_Operator_out6829_out1            : std_logic;
  SIGNAL Logical_Operator_out6830_out1            : std_logic;
  SIGNAL Logical_Operator_out6831_out1            : std_logic;
  SIGNAL Logical_Operator_out6832_out1            : std_logic;
  SIGNAL Logical_Operator_out6833_out1            : std_logic;
  SIGNAL Logical_Operator_out6834_out1            : std_logic;
  SIGNAL Logical_Operator_out6835_out1            : std_logic;
  SIGNAL Logical_Operator_out6836_out1            : std_logic;
  SIGNAL Logical_Operator_out6837_out1            : std_logic;
  SIGNAL Logical_Operator_out6838_out1            : std_logic;
  SIGNAL Logical_Operator_out6839_out1            : std_logic;
  SIGNAL Logical_Operator_out6840_out1            : std_logic;
  SIGNAL Logical_Operator_out6841_out1            : std_logic;
  SIGNAL Logical_Operator_out6842_out1            : std_logic;
  SIGNAL Logical_Operator_out6843_out1            : std_logic;
  SIGNAL Logical_Operator_out6844_out1            : std_logic;
  SIGNAL Logical_Operator_out6845_out1            : std_logic;
  SIGNAL Logical_Operator_out6846_out1            : std_logic;
  SIGNAL Logical_Operator_out6847_out1            : std_logic;
  SIGNAL Logical_Operator_out6848_out1            : std_logic;
  SIGNAL Logical_Operator_out6849_out1            : std_logic;
  SIGNAL Logical_Operator_out6850_out1            : std_logic;
  SIGNAL Logical_Operator_out6851_out1            : std_logic;
  SIGNAL Logical_Operator_out6852_out1            : std_logic;
  SIGNAL Logical_Operator_out6853_out1            : std_logic;
  SIGNAL Logical_Operator_out6854_out1            : std_logic;
  SIGNAL Logical_Operator_out6855_out1            : std_logic;
  SIGNAL Logical_Operator_out6856_out1            : std_logic;
  SIGNAL Logical_Operator_out6857_out1            : std_logic;
  SIGNAL Logical_Operator_out6858_out1            : std_logic;
  SIGNAL Logical_Operator_out6859_out1            : std_logic;
  SIGNAL Logical_Operator_out6860_out1            : std_logic;
  SIGNAL Logical_Operator_out6861_out1            : std_logic;
  SIGNAL Logical_Operator_out6862_out1            : std_logic;
  SIGNAL Logical_Operator_out6863_out1            : std_logic;
  SIGNAL Logical_Operator_out6864_out1            : std_logic;
  SIGNAL Logical_Operator_out6865_out1            : std_logic;
  SIGNAL Logical_Operator_out6866_out1            : std_logic;
  SIGNAL Logical_Operator_out6867_out1            : std_logic;
  SIGNAL Logical_Operator_out6868_out1            : std_logic;
  SIGNAL Logical_Operator_out6869_out1            : std_logic;
  SIGNAL Logical_Operator_out6870_out1            : std_logic;
  SIGNAL Logical_Operator_out6871_out1            : std_logic;
  SIGNAL Logical_Operator_out6872_out1            : std_logic;
  SIGNAL Logical_Operator_out6873_out1            : std_logic;
  SIGNAL Logical_Operator_out6874_out1            : std_logic;
  SIGNAL Logical_Operator_out6875_out1            : std_logic;
  SIGNAL Logical_Operator_out6876_out1            : std_logic;
  SIGNAL Logical_Operator_out6877_out1            : std_logic;
  SIGNAL Logical_Operator_out6878_out1            : std_logic;
  SIGNAL Logical_Operator_out6879_out1            : std_logic;
  SIGNAL Logical_Operator_out6880_out1            : std_logic;
  SIGNAL Logical_Operator_out6881_out1            : std_logic;
  SIGNAL Logical_Operator_out6882_out1            : std_logic;
  SIGNAL Logical_Operator_out6883_out1            : std_logic;
  SIGNAL Logical_Operator_out6884_out1            : std_logic;
  SIGNAL Logical_Operator_out6885_out1            : std_logic;
  SIGNAL Logical_Operator_out6886_out1            : std_logic;
  SIGNAL Logical_Operator_out6887_out1            : std_logic;
  SIGNAL Logical_Operator_out6888_out1            : std_logic;
  SIGNAL Logical_Operator_out6889_out1            : std_logic;
  SIGNAL Logical_Operator_out6890_out1            : std_logic;
  SIGNAL Logical_Operator_out6891_out1            : std_logic;
  SIGNAL Logical_Operator_out6892_out1            : std_logic;
  SIGNAL Logical_Operator_out6893_out1            : std_logic;
  SIGNAL Logical_Operator_out6894_out1            : std_logic;
  SIGNAL Logical_Operator_out6895_out1            : std_logic;
  SIGNAL Logical_Operator_out6896_out1            : std_logic;
  SIGNAL Logical_Operator_out6897_out1            : std_logic;
  SIGNAL Logical_Operator_out6898_out1            : std_logic;
  SIGNAL Logical_Operator_out6899_out1            : std_logic;
  SIGNAL Logical_Operator_out6900_out1            : std_logic;
  SIGNAL Logical_Operator_out6901_out1            : std_logic;
  SIGNAL Logical_Operator_out6902_out1            : std_logic;
  SIGNAL Logical_Operator_out6903_out1            : std_logic;
  SIGNAL Logical_Operator_out6904_out1            : std_logic;
  SIGNAL Logical_Operator_out6905_out1            : std_logic;
  SIGNAL Logical_Operator_out6906_out1            : std_logic;
  SIGNAL Logical_Operator_out6907_out1            : std_logic;
  SIGNAL Logical_Operator_out6908_out1            : std_logic;
  SIGNAL Logical_Operator_out6909_out1            : std_logic;
  SIGNAL Logical_Operator_out6910_out1            : std_logic;
  SIGNAL Logical_Operator_out6911_out1            : std_logic;
  SIGNAL Logical_Operator_out6912_out1            : std_logic;
  SIGNAL Logical_Operator_out6913_out1            : std_logic;
  SIGNAL Logical_Operator_out6914_out1            : std_logic;
  SIGNAL Logical_Operator_out6915_out1            : std_logic;
  SIGNAL Logical_Operator_out6916_out1            : std_logic;
  SIGNAL Logical_Operator_out6917_out1            : std_logic;
  SIGNAL Logical_Operator_out6918_out1            : std_logic;
  SIGNAL Logical_Operator_out6919_out1            : std_logic;
  SIGNAL Logical_Operator_out6920_out1            : std_logic;
  SIGNAL Logical_Operator_out6921_out1            : std_logic;
  SIGNAL Logical_Operator_out6922_out1            : std_logic;
  SIGNAL Logical_Operator_out6923_out1            : std_logic;
  SIGNAL Logical_Operator_out6924_out1            : std_logic;
  SIGNAL Logical_Operator_out6925_out1            : std_logic;
  SIGNAL Logical_Operator_out6926_out1            : std_logic;
  SIGNAL Logical_Operator_out6927_out1            : std_logic;
  SIGNAL Logical_Operator_out6928_out1            : std_logic;
  SIGNAL Logical_Operator_out6929_out1            : std_logic;
  SIGNAL Logical_Operator_out6930_out1            : std_logic;
  SIGNAL Logical_Operator_out6931_out1            : std_logic;
  SIGNAL Logical_Operator_out6932_out1            : std_logic;
  SIGNAL Logical_Operator_out6933_out1            : std_logic;
  SIGNAL Logical_Operator_out6934_out1            : std_logic;
  SIGNAL Logical_Operator_out6935_out1            : std_logic;
  SIGNAL Logical_Operator_out6936_out1            : std_logic;
  SIGNAL Logical_Operator_out6937_out1            : std_logic;
  SIGNAL Logical_Operator_out6938_out1            : std_logic;
  SIGNAL Logical_Operator_out6939_out1            : std_logic;
  SIGNAL Logical_Operator_out6940_out1            : std_logic;
  SIGNAL Logical_Operator_out6941_out1            : std_logic;
  SIGNAL Logical_Operator_out6942_out1            : std_logic;
  SIGNAL Logical_Operator_out6943_out1            : std_logic;
  SIGNAL Logical_Operator_out6944_out1            : std_logic;
  SIGNAL Logical_Operator_out6945_out1            : std_logic;
  SIGNAL Logical_Operator_out6946_out1            : std_logic;
  SIGNAL Logical_Operator_out6947_out1            : std_logic;
  SIGNAL Logical_Operator_out6948_out1            : std_logic;
  SIGNAL Logical_Operator_out6949_out1            : std_logic;
  SIGNAL Logical_Operator_out6950_out1            : std_logic;
  SIGNAL Logical_Operator_out6951_out1            : std_logic;
  SIGNAL Logical_Operator_out6952_out1            : std_logic;
  SIGNAL Logical_Operator_out6953_out1            : std_logic;
  SIGNAL Logical_Operator_out6954_out1            : std_logic;
  SIGNAL Logical_Operator_out6955_out1            : std_logic;
  SIGNAL Logical_Operator_out6956_out1            : std_logic;
  SIGNAL Logical_Operator_out6957_out1            : std_logic;
  SIGNAL Logical_Operator_out6958_out1            : std_logic;
  SIGNAL Logical_Operator_out6959_out1            : std_logic;
  SIGNAL Logical_Operator_out6960_out1            : std_logic;
  SIGNAL Logical_Operator_out6961_out1            : std_logic;
  SIGNAL Logical_Operator_out6962_out1            : std_logic;
  SIGNAL Logical_Operator_out6963_out1            : std_logic;
  SIGNAL Logical_Operator_out6964_out1            : std_logic;
  SIGNAL Logical_Operator_out6965_out1            : std_logic;
  SIGNAL Logical_Operator_out6966_out1            : std_logic;
  SIGNAL Logical_Operator_out6967_out1            : std_logic;
  SIGNAL Logical_Operator_out6968_out1            : std_logic;
  SIGNAL Logical_Operator_out6969_out1            : std_logic;
  SIGNAL Logical_Operator_out6970_out1            : std_logic;
  SIGNAL Logical_Operator_out6971_out1            : std_logic;
  SIGNAL Logical_Operator_out6972_out1            : std_logic;
  SIGNAL Logical_Operator_out6973_out1            : std_logic;
  SIGNAL Logical_Operator_out6974_out1            : std_logic;
  SIGNAL Logical_Operator_out6975_out1            : std_logic;
  SIGNAL Logical_Operator_out6976_out1            : std_logic;
  SIGNAL Logical_Operator_out6977_out1            : std_logic;
  SIGNAL Logical_Operator_out6978_out1            : std_logic;
  SIGNAL Logical_Operator_out6979_out1            : std_logic;
  SIGNAL Logical_Operator_out6980_out1            : std_logic;
  SIGNAL Logical_Operator_out6981_out1            : std_logic;
  SIGNAL Logical_Operator_out6982_out1            : std_logic;
  SIGNAL Logical_Operator_out6983_out1            : std_logic;
  SIGNAL Logical_Operator_out6984_out1            : std_logic;
  SIGNAL Logical_Operator_out6985_out1            : std_logic;
  SIGNAL Logical_Operator_out6986_out1            : std_logic;
  SIGNAL Logical_Operator_out6987_out1            : std_logic;
  SIGNAL Logical_Operator_out6988_out1            : std_logic;
  SIGNAL Logical_Operator_out6989_out1            : std_logic;
  SIGNAL Logical_Operator_out6990_out1            : std_logic;
  SIGNAL Logical_Operator_out6991_out1            : std_logic;
  SIGNAL Logical_Operator_out6992_out1            : std_logic;
  SIGNAL Logical_Operator_out6993_out1            : std_logic;
  SIGNAL Logical_Operator_out6994_out1            : std_logic;
  SIGNAL Logical_Operator_out6995_out1            : std_logic;
  SIGNAL Logical_Operator_out6996_out1            : std_logic;
  SIGNAL Logical_Operator_out6997_out1            : std_logic;
  SIGNAL Logical_Operator_out6998_out1            : std_logic;
  SIGNAL Logical_Operator_out6999_out1            : std_logic;
  SIGNAL Logical_Operator_out7000_out1            : std_logic;
  SIGNAL Logical_Operator_out7001_out1            : std_logic;
  SIGNAL Logical_Operator_out7002_out1            : std_logic;
  SIGNAL Logical_Operator_out7003_out1            : std_logic;
  SIGNAL Logical_Operator_out7004_out1            : std_logic;
  SIGNAL Logical_Operator_out7005_out1            : std_logic;
  SIGNAL Logical_Operator_out7006_out1            : std_logic;
  SIGNAL Logical_Operator_out7007_out1            : std_logic;
  SIGNAL Logical_Operator_out7008_out1            : std_logic;
  SIGNAL Logical_Operator_out7009_out1            : std_logic;
  SIGNAL Logical_Operator_out7010_out1            : std_logic;
  SIGNAL Logical_Operator_out7011_out1            : std_logic;
  SIGNAL Logical_Operator_out7012_out1            : std_logic;
  SIGNAL Logical_Operator_out7013_out1            : std_logic;
  SIGNAL Logical_Operator_out7014_out1            : std_logic;
  SIGNAL Logical_Operator_out7015_out1            : std_logic;
  SIGNAL Logical_Operator_out7016_out1            : std_logic;
  SIGNAL Logical_Operator_out7017_out1            : std_logic;
  SIGNAL Logical_Operator_out7018_out1            : std_logic;
  SIGNAL Logical_Operator_out7019_out1            : std_logic;
  SIGNAL Logical_Operator_out7020_out1            : std_logic;
  SIGNAL Logical_Operator_out7021_out1            : std_logic;
  SIGNAL Logical_Operator_out7022_out1            : std_logic;
  SIGNAL Logical_Operator_out7023_out1            : std_logic;
  SIGNAL Logical_Operator_out7024_out1            : std_logic;
  SIGNAL Logical_Operator_out7025_out1            : std_logic;
  SIGNAL Logical_Operator_out7026_out1            : std_logic;
  SIGNAL Logical_Operator_out7027_out1            : std_logic;
  SIGNAL Logical_Operator_out7028_out1            : std_logic;
  SIGNAL Logical_Operator_out7029_out1            : std_logic;
  SIGNAL Logical_Operator_out7030_out1            : std_logic;
  SIGNAL Logical_Operator_out7031_out1            : std_logic;
  SIGNAL Logical_Operator_out7032_out1            : std_logic;
  SIGNAL Logical_Operator_out7033_out1            : std_logic;
  SIGNAL Logical_Operator_out7034_out1            : std_logic;
  SIGNAL Logical_Operator_out7035_out1            : std_logic;
  SIGNAL Logical_Operator_out7036_out1            : std_logic;
  SIGNAL Logical_Operator_out7037_out1            : std_logic;
  SIGNAL Logical_Operator_out7038_out1            : std_logic;
  SIGNAL Logical_Operator_out7039_out1            : std_logic;
  SIGNAL Logical_Operator_out7040_out1            : std_logic;
  SIGNAL Logical_Operator_out7041_out1            : std_logic;
  SIGNAL Logical_Operator_out7042_out1            : std_logic;
  SIGNAL Logical_Operator_out7043_out1            : std_logic;
  SIGNAL Logical_Operator_out7044_out1            : std_logic;
  SIGNAL Logical_Operator_out7045_out1            : std_logic;
  SIGNAL Logical_Operator_out7046_out1            : std_logic;
  SIGNAL Logical_Operator_out7047_out1            : std_logic;
  SIGNAL Logical_Operator_out7048_out1            : std_logic;
  SIGNAL Logical_Operator_out7049_out1            : std_logic;
  SIGNAL Logical_Operator_out7050_out1            : std_logic;
  SIGNAL Logical_Operator_out7051_out1            : std_logic;
  SIGNAL Logical_Operator_out7052_out1            : std_logic;
  SIGNAL Logical_Operator_out7053_out1            : std_logic;
  SIGNAL Logical_Operator_out7054_out1            : std_logic;
  SIGNAL Logical_Operator_out7055_out1            : std_logic;
  SIGNAL Logical_Operator_out7056_out1            : std_logic;
  SIGNAL Logical_Operator_out7057_out1            : std_logic;
  SIGNAL Logical_Operator_out7058_out1            : std_logic;
  SIGNAL Logical_Operator_out7059_out1            : std_logic;
  SIGNAL Logical_Operator_out7060_out1            : std_logic;
  SIGNAL Logical_Operator_out7061_out1            : std_logic;
  SIGNAL Logical_Operator_out7062_out1            : std_logic;
  SIGNAL Logical_Operator_out7063_out1            : std_logic;
  SIGNAL Logical_Operator_out7064_out1            : std_logic;
  SIGNAL Logical_Operator_out7065_out1            : std_logic;
  SIGNAL Logical_Operator_out7066_out1            : std_logic;
  SIGNAL Logical_Operator_out7067_out1            : std_logic;
  SIGNAL Logical_Operator_out7068_out1            : std_logic;
  SIGNAL Logical_Operator_out7069_out1            : std_logic;
  SIGNAL Logical_Operator_out7070_out1            : std_logic;
  SIGNAL Logical_Operator_out7071_out1            : std_logic;
  SIGNAL Logical_Operator_out7072_out1            : std_logic;
  SIGNAL Logical_Operator_out7073_out1            : std_logic;
  SIGNAL Logical_Operator_out7074_out1            : std_logic;
  SIGNAL Logical_Operator_out7075_out1            : std_logic;
  SIGNAL Logical_Operator_out7076_out1            : std_logic;
  SIGNAL Logical_Operator_out7077_out1            : std_logic;
  SIGNAL Logical_Operator_out7078_out1            : std_logic;
  SIGNAL Logical_Operator_out7079_out1            : std_logic;
  SIGNAL Logical_Operator_out7080_out1            : std_logic;
  SIGNAL Logical_Operator_out7081_out1            : std_logic;
  SIGNAL Logical_Operator_out7082_out1            : std_logic;
  SIGNAL Logical_Operator_out7083_out1            : std_logic;
  SIGNAL Logical_Operator_out7084_out1            : std_logic;
  SIGNAL Logical_Operator_out7085_out1            : std_logic;
  SIGNAL Logical_Operator_out7086_out1            : std_logic;
  SIGNAL Logical_Operator_out7087_out1            : std_logic;
  SIGNAL Logical_Operator_out7088_out1            : std_logic;
  SIGNAL Logical_Operator_out7089_out1            : std_logic;
  SIGNAL Logical_Operator_out7090_out1            : std_logic;
  SIGNAL Logical_Operator_out7091_out1            : std_logic;
  SIGNAL Logical_Operator_out7092_out1            : std_logic;
  SIGNAL Logical_Operator_out7093_out1            : std_logic;
  SIGNAL Logical_Operator_out7094_out1            : std_logic;
  SIGNAL Logical_Operator_out7095_out1            : std_logic;
  SIGNAL Logical_Operator_out7096_out1            : std_logic;
  SIGNAL Logical_Operator_out7097_out1            : std_logic;
  SIGNAL Logical_Operator_out7098_out1            : std_logic;
  SIGNAL Logical_Operator_out7099_out1            : std_logic;
  SIGNAL Logical_Operator_out7100_out1            : std_logic;
  SIGNAL Logical_Operator_out7101_out1            : std_logic;
  SIGNAL Logical_Operator_out7102_out1            : std_logic;
  SIGNAL Logical_Operator_out7103_out1            : std_logic;
  SIGNAL Logical_Operator_out7104_out1            : std_logic;
  SIGNAL Logical_Operator_out7105_out1            : std_logic;
  SIGNAL Logical_Operator_out7106_out1            : std_logic;
  SIGNAL Logical_Operator_out7107_out1            : std_logic;
  SIGNAL Logical_Operator_out7108_out1            : std_logic;
  SIGNAL Logical_Operator_out7109_out1            : std_logic;
  SIGNAL Logical_Operator_out7110_out1            : std_logic;
  SIGNAL Logical_Operator_out7111_out1            : std_logic;
  SIGNAL Logical_Operator_out7112_out1            : std_logic;
  SIGNAL Logical_Operator_out7113_out1            : std_logic;
  SIGNAL Logical_Operator_out7114_out1            : std_logic;
  SIGNAL Logical_Operator_out7115_out1            : std_logic;
  SIGNAL Logical_Operator_out7116_out1            : std_logic;
  SIGNAL Logical_Operator_out7117_out1            : std_logic;
  SIGNAL Logical_Operator_out7118_out1            : std_logic;
  SIGNAL Logical_Operator_out7119_out1            : std_logic;
  SIGNAL Logical_Operator_out7120_out1            : std_logic;
  SIGNAL Logical_Operator_out7121_out1            : std_logic;
  SIGNAL Logical_Operator_out7122_out1            : std_logic;
  SIGNAL Logical_Operator_out7123_out1            : std_logic;
  SIGNAL Logical_Operator_out7124_out1            : std_logic;
  SIGNAL Logical_Operator_out7125_out1            : std_logic;
  SIGNAL Logical_Operator_out7126_out1            : std_logic;
  SIGNAL Logical_Operator_out7127_out1            : std_logic;
  SIGNAL Logical_Operator_out7128_out1            : std_logic;
  SIGNAL Logical_Operator_out7129_out1            : std_logic;
  SIGNAL Logical_Operator_out7130_out1            : std_logic;
  SIGNAL Logical_Operator_out7131_out1            : std_logic;
  SIGNAL Logical_Operator_out7132_out1            : std_logic;
  SIGNAL Logical_Operator_out7133_out1            : std_logic;
  SIGNAL Logical_Operator_out7134_out1            : std_logic;
  SIGNAL Logical_Operator_out7135_out1            : std_logic;
  SIGNAL Logical_Operator_out7136_out1            : std_logic;
  SIGNAL Logical_Operator_out7137_out1            : std_logic;
  SIGNAL Logical_Operator_out7138_out1            : std_logic;
  SIGNAL Logical_Operator_out7139_out1            : std_logic;
  SIGNAL Logical_Operator_out7140_out1            : std_logic;
  SIGNAL Logical_Operator_out7141_out1            : std_logic;
  SIGNAL Logical_Operator_out7142_out1            : std_logic;
  SIGNAL Logical_Operator_out7143_out1            : std_logic;
  SIGNAL Logical_Operator_out7144_out1            : std_logic;
  SIGNAL Logical_Operator_out7145_out1            : std_logic;
  SIGNAL Logical_Operator_out7146_out1            : std_logic;
  SIGNAL Logical_Operator_out7147_out1            : std_logic;
  SIGNAL Logical_Operator_out7148_out1            : std_logic;
  SIGNAL Logical_Operator_out7149_out1            : std_logic;
  SIGNAL Logical_Operator_out7150_out1            : std_logic;
  SIGNAL Logical_Operator_out7151_out1            : std_logic;
  SIGNAL Logical_Operator_out7152_out1            : std_logic;
  SIGNAL Logical_Operator_out7153_out1            : std_logic;
  SIGNAL Logical_Operator_out7154_out1            : std_logic;
  SIGNAL Logical_Operator_out7155_out1            : std_logic;
  SIGNAL Logical_Operator_out7156_out1            : std_logic;
  SIGNAL Logical_Operator_out7157_out1            : std_logic;
  SIGNAL Logical_Operator_out7158_out1            : std_logic;
  SIGNAL Logical_Operator_out7159_out1            : std_logic;
  SIGNAL Logical_Operator_out7160_out1            : std_logic;
  SIGNAL Logical_Operator_out7161_out1            : std_logic;
  SIGNAL Logical_Operator_out7162_out1            : std_logic;
  SIGNAL Logical_Operator_out7163_out1            : std_logic;
  SIGNAL Logical_Operator_out7164_out1            : std_logic;
  SIGNAL Logical_Operator_out7165_out1            : std_logic;
  SIGNAL Logical_Operator_out7166_out1            : std_logic;
  SIGNAL Logical_Operator_out7167_out1            : std_logic;
  SIGNAL Logical_Operator_out7168_out1            : std_logic;
  SIGNAL Logical_Operator_out7169_out1            : std_logic;
  SIGNAL Logical_Operator_out7170_out1            : std_logic;
  SIGNAL Logical_Operator_out7171_out1            : std_logic;
  SIGNAL Logical_Operator_out7172_out1            : std_logic;
  SIGNAL Logical_Operator_out7173_out1            : std_logic;
  SIGNAL Logical_Operator_out7174_out1            : std_logic;
  SIGNAL Logical_Operator_out7175_out1            : std_logic;
  SIGNAL Logical_Operator_out7176_out1            : std_logic;
  SIGNAL Logical_Operator_out7177_out1            : std_logic;
  SIGNAL Logical_Operator_out7178_out1            : std_logic;
  SIGNAL Logical_Operator_out7179_out1            : std_logic;
  SIGNAL Logical_Operator_out7180_out1            : std_logic;
  SIGNAL Logical_Operator_out7181_out1            : std_logic;
  SIGNAL Logical_Operator_out7182_out1            : std_logic;
  SIGNAL Logical_Operator_out7183_out1            : std_logic;
  SIGNAL Logical_Operator_out7184_out1            : std_logic;
  SIGNAL Logical_Operator_out7185_out1            : std_logic;
  SIGNAL Logical_Operator_out7186_out1            : std_logic;
  SIGNAL Logical_Operator_out7187_out1            : std_logic;
  SIGNAL Logical_Operator_out7188_out1            : std_logic;
  SIGNAL Logical_Operator_out7189_out1            : std_logic;
  SIGNAL Logical_Operator_out7190_out1            : std_logic;
  SIGNAL Logical_Operator_out7191_out1            : std_logic;
  SIGNAL Logical_Operator_out7192_out1            : std_logic;
  SIGNAL Logical_Operator_out7193_out1            : std_logic;
  SIGNAL Logical_Operator_out7194_out1            : std_logic;
  SIGNAL Logical_Operator_out7195_out1            : std_logic;
  SIGNAL Logical_Operator_out7196_out1            : std_logic;
  SIGNAL Logical_Operator_out7197_out1            : std_logic;
  SIGNAL Logical_Operator_out7198_out1            : std_logic;
  SIGNAL Logical_Operator_out7199_out1            : std_logic;
  SIGNAL Logical_Operator_out7200_out1            : std_logic;
  SIGNAL Logical_Operator_out7201_out1            : std_logic;
  SIGNAL Logical_Operator_out7202_out1            : std_logic;
  SIGNAL Logical_Operator_out7203_out1            : std_logic;
  SIGNAL Logical_Operator_out7204_out1            : std_logic;
  SIGNAL Logical_Operator_out7205_out1            : std_logic;
  SIGNAL Logical_Operator_out7206_out1            : std_logic;
  SIGNAL Logical_Operator_out7207_out1            : std_logic;
  SIGNAL Logical_Operator_out7208_out1            : std_logic;
  SIGNAL Logical_Operator_out7209_out1            : std_logic;
  SIGNAL Logical_Operator_out7210_out1            : std_logic;
  SIGNAL Logical_Operator_out7211_out1            : std_logic;
  SIGNAL Logical_Operator_out7212_out1            : std_logic;
  SIGNAL Logical_Operator_out7213_out1            : std_logic;
  SIGNAL Logical_Operator_out7214_out1            : std_logic;
  SIGNAL Logical_Operator_out7215_out1            : std_logic;
  SIGNAL Logical_Operator_out7216_out1            : std_logic;
  SIGNAL Logical_Operator_out7217_out1            : std_logic;
  SIGNAL Logical_Operator_out7218_out1            : std_logic;
  SIGNAL Logical_Operator_out7219_out1            : std_logic;
  SIGNAL Logical_Operator_out7220_out1            : std_logic;
  SIGNAL Logical_Operator_out7221_out1            : std_logic;
  SIGNAL Logical_Operator_out7222_out1            : std_logic;
  SIGNAL Logical_Operator_out7223_out1            : std_logic;
  SIGNAL Logical_Operator_out7224_out1            : std_logic;
  SIGNAL Logical_Operator_out7225_out1            : std_logic;
  SIGNAL Logical_Operator_out7226_out1            : std_logic;
  SIGNAL Logical_Operator_out7227_out1            : std_logic;
  SIGNAL Logical_Operator_out7228_out1            : std_logic;
  SIGNAL Logical_Operator_out7229_out1            : std_logic;
  SIGNAL Logical_Operator_out7230_out1            : std_logic;
  SIGNAL Logical_Operator_out7231_out1            : std_logic;
  SIGNAL Logical_Operator_out7232_out1            : std_logic;
  SIGNAL Logical_Operator_out7233_out1            : std_logic;
  SIGNAL Logical_Operator_out7234_out1            : std_logic;
  SIGNAL Logical_Operator_out7235_out1            : std_logic;
  SIGNAL Logical_Operator_out7236_out1            : std_logic;
  SIGNAL Logical_Operator_out7237_out1            : std_logic;
  SIGNAL Logical_Operator_out7238_out1            : std_logic;
  SIGNAL Logical_Operator_out7239_out1            : std_logic;
  SIGNAL Logical_Operator_out7240_out1            : std_logic;
  SIGNAL Logical_Operator_out7241_out1            : std_logic;
  SIGNAL Logical_Operator_out7242_out1            : std_logic;
  SIGNAL Logical_Operator_out7243_out1            : std_logic;
  SIGNAL Logical_Operator_out7244_out1            : std_logic;
  SIGNAL Logical_Operator_out7245_out1            : std_logic;
  SIGNAL Logical_Operator_out7246_out1            : std_logic;
  SIGNAL Logical_Operator_out7247_out1            : std_logic;
  SIGNAL Logical_Operator_out7248_out1            : std_logic;
  SIGNAL Logical_Operator_out7249_out1            : std_logic;
  SIGNAL Logical_Operator_out7250_out1            : std_logic;
  SIGNAL Logical_Operator_out7251_out1            : std_logic;
  SIGNAL Logical_Operator_out7252_out1            : std_logic;
  SIGNAL Logical_Operator_out7253_out1            : std_logic;
  SIGNAL Logical_Operator_out7254_out1            : std_logic;
  SIGNAL Logical_Operator_out7255_out1            : std_logic;
  SIGNAL Logical_Operator_out7256_out1            : std_logic;
  SIGNAL Logical_Operator_out7257_out1            : std_logic;
  SIGNAL Logical_Operator_out7258_out1            : std_logic;
  SIGNAL Logical_Operator_out7259_out1            : std_logic;
  SIGNAL Logical_Operator_out7260_out1            : std_logic;
  SIGNAL Logical_Operator_out7261_out1            : std_logic;
  SIGNAL Logical_Operator_out7262_out1            : std_logic;
  SIGNAL Logical_Operator_out7263_out1            : std_logic;
  SIGNAL Logical_Operator_out7264_out1            : std_logic;
  SIGNAL Logical_Operator_out7265_out1            : std_logic;
  SIGNAL Logical_Operator_out7266_out1            : std_logic;
  SIGNAL Logical_Operator_out7267_out1            : std_logic;
  SIGNAL Logical_Operator_out7268_out1            : std_logic;
  SIGNAL Logical_Operator_out7269_out1            : std_logic;
  SIGNAL Logical_Operator_out7270_out1            : std_logic;
  SIGNAL Logical_Operator_out7271_out1            : std_logic;
  SIGNAL Logical_Operator_out7272_out1            : std_logic;
  SIGNAL Logical_Operator_out7273_out1            : std_logic;
  SIGNAL Logical_Operator_out7274_out1            : std_logic;
  SIGNAL Logical_Operator_out7275_out1            : std_logic;
  SIGNAL Logical_Operator_out7276_out1            : std_logic;
  SIGNAL Logical_Operator_out7277_out1            : std_logic;
  SIGNAL Logical_Operator_out7278_out1            : std_logic;
  SIGNAL Logical_Operator_out7279_out1            : std_logic;
  SIGNAL Logical_Operator_out7280_out1            : std_logic;
  SIGNAL Logical_Operator_out7281_out1            : std_logic;
  SIGNAL Logical_Operator_out7282_out1            : std_logic;
  SIGNAL Logical_Operator_out7283_out1            : std_logic;
  SIGNAL Logical_Operator_out7284_out1            : std_logic;
  SIGNAL Logical_Operator_out7285_out1            : std_logic;
  SIGNAL Logical_Operator_out7286_out1            : std_logic;
  SIGNAL Logical_Operator_out7287_out1            : std_logic;
  SIGNAL Logical_Operator_out7288_out1            : std_logic;
  SIGNAL Logical_Operator_out7289_out1            : std_logic;
  SIGNAL Logical_Operator_out7290_out1            : std_logic;
  SIGNAL Logical_Operator_out7291_out1            : std_logic;
  SIGNAL Logical_Operator_out7292_out1            : std_logic;
  SIGNAL Logical_Operator_out7293_out1            : std_logic;
  SIGNAL Logical_Operator_out7294_out1            : std_logic;
  SIGNAL Logical_Operator_out7295_out1            : std_logic;
  SIGNAL Logical_Operator_out7296_out1            : std_logic;
  SIGNAL Logical_Operator_out7297_out1            : std_logic;
  SIGNAL Logical_Operator_out7298_out1            : std_logic;
  SIGNAL Logical_Operator_out7299_out1            : std_logic;
  SIGNAL Logical_Operator_out7300_out1            : std_logic;
  SIGNAL Logical_Operator_out7301_out1            : std_logic;
  SIGNAL Logical_Operator_out7302_out1            : std_logic;
  SIGNAL Logical_Operator_out7303_out1            : std_logic;
  SIGNAL Logical_Operator_out7304_out1            : std_logic;
  SIGNAL Logical_Operator_out7305_out1            : std_logic;
  SIGNAL Logical_Operator_out7306_out1            : std_logic;
  SIGNAL Logical_Operator_out7307_out1            : std_logic;
  SIGNAL Logical_Operator_out7308_out1            : std_logic;
  SIGNAL Logical_Operator_out7309_out1            : std_logic;
  SIGNAL Logical_Operator_out7310_out1            : std_logic;
  SIGNAL Logical_Operator_out7311_out1            : std_logic;
  SIGNAL Logical_Operator_out7312_out1            : std_logic;
  SIGNAL Logical_Operator_out7313_out1            : std_logic;
  SIGNAL Logical_Operator_out7314_out1            : std_logic;
  SIGNAL Logical_Operator_out7315_out1            : std_logic;
  SIGNAL Logical_Operator_out7316_out1            : std_logic;
  SIGNAL Logical_Operator_out7317_out1            : std_logic;
  SIGNAL Logical_Operator_out7318_out1            : std_logic;
  SIGNAL Logical_Operator_out7319_out1            : std_logic;
  SIGNAL Logical_Operator_out7320_out1            : std_logic;
  SIGNAL Logical_Operator_out7321_out1            : std_logic;
  SIGNAL Logical_Operator_out7322_out1            : std_logic;
  SIGNAL Logical_Operator_out7323_out1            : std_logic;
  SIGNAL Logical_Operator_out7324_out1            : std_logic;
  SIGNAL Logical_Operator_out7325_out1            : std_logic;
  SIGNAL Logical_Operator_out7326_out1            : std_logic;
  SIGNAL Logical_Operator_out7327_out1            : std_logic;
  SIGNAL Logical_Operator_out7328_out1            : std_logic;
  SIGNAL Logical_Operator_out7329_out1            : std_logic;
  SIGNAL Logical_Operator_out7330_out1            : std_logic;
  SIGNAL Logical_Operator_out7331_out1            : std_logic;
  SIGNAL Logical_Operator_out7332_out1            : std_logic;
  SIGNAL Logical_Operator_out7333_out1            : std_logic;
  SIGNAL Logical_Operator_out7334_out1            : std_logic;
  SIGNAL Logical_Operator_out7335_out1            : std_logic;
  SIGNAL Logical_Operator_out7336_out1            : std_logic;
  SIGNAL Logical_Operator_out7337_out1            : std_logic;
  SIGNAL Logical_Operator_out7338_out1            : std_logic;
  SIGNAL Logical_Operator_out7339_out1            : std_logic;
  SIGNAL Logical_Operator_out7340_out1            : std_logic;
  SIGNAL Logical_Operator_out7341_out1            : std_logic;
  SIGNAL Logical_Operator_out7342_out1            : std_logic;
  SIGNAL Logical_Operator_out7343_out1            : std_logic;
  SIGNAL Logical_Operator_out7344_out1            : std_logic;
  SIGNAL Logical_Operator_out7345_out1            : std_logic;
  SIGNAL Logical_Operator_out7346_out1            : std_logic;
  SIGNAL Logical_Operator_out7347_out1            : std_logic;
  SIGNAL Logical_Operator_out7348_out1            : std_logic;
  SIGNAL Logical_Operator_out7349_out1            : std_logic;
  SIGNAL Logical_Operator_out7350_out1            : std_logic;
  SIGNAL Logical_Operator_out7351_out1            : std_logic;
  SIGNAL Logical_Operator_out7352_out1            : std_logic;
  SIGNAL Logical_Operator_out7353_out1            : std_logic;
  SIGNAL Logical_Operator_out7354_out1            : std_logic;
  SIGNAL Logical_Operator_out7355_out1            : std_logic;
  SIGNAL Logical_Operator_out7356_out1            : std_logic;
  SIGNAL Logical_Operator_out7357_out1            : std_logic;
  SIGNAL Logical_Operator_out7358_out1            : std_logic;
  SIGNAL Logical_Operator_out7359_out1            : std_logic;
  SIGNAL Logical_Operator_out7360_out1            : std_logic;
  SIGNAL Logical_Operator_out7361_out1            : std_logic;
  SIGNAL Logical_Operator_out7362_out1            : std_logic;
  SIGNAL Logical_Operator_out7363_out1            : std_logic;
  SIGNAL Logical_Operator_out7364_out1            : std_logic;
  SIGNAL Logical_Operator_out7365_out1            : std_logic;
  SIGNAL Logical_Operator_out7366_out1            : std_logic;
  SIGNAL Logical_Operator_out7367_out1            : std_logic;
  SIGNAL Logical_Operator_out7368_out1            : std_logic;
  SIGNAL Logical_Operator_out7369_out1            : std_logic;
  SIGNAL Logical_Operator_out7370_out1            : std_logic;
  SIGNAL Logical_Operator_out7371_out1            : std_logic;
  SIGNAL Logical_Operator_out7372_out1            : std_logic;
  SIGNAL Logical_Operator_out7373_out1            : std_logic;
  SIGNAL Logical_Operator_out7374_out1            : std_logic;
  SIGNAL Logical_Operator_out7375_out1            : std_logic;
  SIGNAL Logical_Operator_out7376_out1            : std_logic;
  SIGNAL Logical_Operator_out7377_out1            : std_logic;
  SIGNAL Logical_Operator_out7378_out1            : std_logic;
  SIGNAL Logical_Operator_out7379_out1            : std_logic;
  SIGNAL Logical_Operator_out7380_out1            : std_logic;
  SIGNAL Logical_Operator_out7381_out1            : std_logic;
  SIGNAL Logical_Operator_out7382_out1            : std_logic;
  SIGNAL Logical_Operator_out7383_out1            : std_logic;
  SIGNAL Logical_Operator_out7384_out1            : std_logic;
  SIGNAL Logical_Operator_out7385_out1            : std_logic;
  SIGNAL Logical_Operator_out7386_out1            : std_logic;
  SIGNAL Logical_Operator_out7387_out1            : std_logic;
  SIGNAL Logical_Operator_out7388_out1            : std_logic;
  SIGNAL Logical_Operator_out7389_out1            : std_logic;
  SIGNAL Logical_Operator_out7390_out1            : std_logic;
  SIGNAL Logical_Operator_out7391_out1            : std_logic;
  SIGNAL Logical_Operator_out7392_out1            : std_logic;
  SIGNAL Logical_Operator_out7393_out1            : std_logic;
  SIGNAL Logical_Operator_out7394_out1            : std_logic;
  SIGNAL Logical_Operator_out7395_out1            : std_logic;
  SIGNAL Logical_Operator_out7396_out1            : std_logic;
  SIGNAL Logical_Operator_out7397_out1            : std_logic;
  SIGNAL Logical_Operator_out7398_out1            : std_logic;
  SIGNAL Logical_Operator_out7399_out1            : std_logic;
  SIGNAL Logical_Operator_out7400_out1            : std_logic;
  SIGNAL Logical_Operator_out7401_out1            : std_logic;
  SIGNAL Logical_Operator_out7402_out1            : std_logic;
  SIGNAL Logical_Operator_out7403_out1            : std_logic;
  SIGNAL Logical_Operator_out7404_out1            : std_logic;
  SIGNAL Logical_Operator_out7405_out1            : std_logic;
  SIGNAL Logical_Operator_out7406_out1            : std_logic;
  SIGNAL Logical_Operator_out7407_out1            : std_logic;
  SIGNAL Logical_Operator_out7408_out1            : std_logic;
  SIGNAL Logical_Operator_out7409_out1            : std_logic;
  SIGNAL Logical_Operator_out7410_out1            : std_logic;
  SIGNAL Logical_Operator_out7411_out1            : std_logic;
  SIGNAL Logical_Operator_out7412_out1            : std_logic;
  SIGNAL Logical_Operator_out7413_out1            : std_logic;
  SIGNAL Logical_Operator_out7414_out1            : std_logic;
  SIGNAL Logical_Operator_out7415_out1            : std_logic;
  SIGNAL Logical_Operator_out7416_out1            : std_logic;
  SIGNAL Logical_Operator_out7417_out1            : std_logic;
  SIGNAL Logical_Operator_out7418_out1            : std_logic;
  SIGNAL Logical_Operator_out7419_out1            : std_logic;
  SIGNAL Logical_Operator_out7420_out1            : std_logic;
  SIGNAL Logical_Operator_out7421_out1            : std_logic;
  SIGNAL Logical_Operator_out7422_out1            : std_logic;
  SIGNAL Logical_Operator_out7423_out1            : std_logic;
  SIGNAL Logical_Operator_out7424_out1            : std_logic;
  SIGNAL Logical_Operator_out7425_out1            : std_logic;
  SIGNAL Logical_Operator_out7426_out1            : std_logic;
  SIGNAL Logical_Operator_out7427_out1            : std_logic;
  SIGNAL Logical_Operator_out7428_out1            : std_logic;
  SIGNAL Logical_Operator_out7429_out1            : std_logic;
  SIGNAL Logical_Operator_out7430_out1            : std_logic;
  SIGNAL Logical_Operator_out7431_out1            : std_logic;
  SIGNAL Logical_Operator_out7432_out1            : std_logic;
  SIGNAL Logical_Operator_out7433_out1            : std_logic;
  SIGNAL Logical_Operator_out7434_out1            : std_logic;
  SIGNAL Logical_Operator_out7435_out1            : std_logic;
  SIGNAL Logical_Operator_out7436_out1            : std_logic;
  SIGNAL Logical_Operator_out7437_out1            : std_logic;
  SIGNAL Logical_Operator_out7438_out1            : std_logic;
  SIGNAL Logical_Operator_out7439_out1            : std_logic;
  SIGNAL Logical_Operator_out7440_out1            : std_logic;
  SIGNAL Logical_Operator_out7441_out1            : std_logic;
  SIGNAL Logical_Operator_out7442_out1            : std_logic;
  SIGNAL Logical_Operator_out7443_out1            : std_logic;
  SIGNAL Logical_Operator_out7444_out1            : std_logic;
  SIGNAL Logical_Operator_out7445_out1            : std_logic;
  SIGNAL Logical_Operator_out7446_out1            : std_logic;
  SIGNAL Logical_Operator_out7447_out1            : std_logic;
  SIGNAL Logical_Operator_out7448_out1            : std_logic;
  SIGNAL Logical_Operator_out7449_out1            : std_logic;
  SIGNAL Logical_Operator_out7450_out1            : std_logic;
  SIGNAL Logical_Operator_out7451_out1            : std_logic;
  SIGNAL Logical_Operator_out7452_out1            : std_logic;
  SIGNAL Logical_Operator_out7453_out1            : std_logic;
  SIGNAL Logical_Operator_out7454_out1            : std_logic;
  SIGNAL Logical_Operator_out7455_out1            : std_logic;
  SIGNAL Logical_Operator_out7456_out1            : std_logic;
  SIGNAL Logical_Operator_out7457_out1            : std_logic;
  SIGNAL Logical_Operator_out7458_out1            : std_logic;
  SIGNAL Logical_Operator_out7459_out1            : std_logic;
  SIGNAL Logical_Operator_out7460_out1            : std_logic;
  SIGNAL Logical_Operator_out7461_out1            : std_logic;
  SIGNAL Logical_Operator_out7462_out1            : std_logic;
  SIGNAL Logical_Operator_out7463_out1            : std_logic;
  SIGNAL Logical_Operator_out7464_out1            : std_logic;
  SIGNAL Logical_Operator_out7465_out1            : std_logic;
  SIGNAL Logical_Operator_out7466_out1            : std_logic;
  SIGNAL Logical_Operator_out7467_out1            : std_logic;
  SIGNAL Logical_Operator_out7468_out1            : std_logic;
  SIGNAL Logical_Operator_out7469_out1            : std_logic;
  SIGNAL Logical_Operator_out7470_out1            : std_logic;
  SIGNAL Logical_Operator_out7471_out1            : std_logic;
  SIGNAL Logical_Operator_out7472_out1            : std_logic;
  SIGNAL Logical_Operator_out7473_out1            : std_logic;
  SIGNAL Logical_Operator_out7474_out1            : std_logic;
  SIGNAL Logical_Operator_out7475_out1            : std_logic;
  SIGNAL Logical_Operator_out7476_out1            : std_logic;
  SIGNAL Logical_Operator_out7477_out1            : std_logic;
  SIGNAL Logical_Operator_out7478_out1            : std_logic;
  SIGNAL Logical_Operator_out7479_out1            : std_logic;
  SIGNAL Logical_Operator_out7480_out1            : std_logic;
  SIGNAL Logical_Operator_out7481_out1            : std_logic;
  SIGNAL Logical_Operator_out7482_out1            : std_logic;
  SIGNAL Logical_Operator_out7483_out1            : std_logic;
  SIGNAL Logical_Operator_out7484_out1            : std_logic;
  SIGNAL Logical_Operator_out7485_out1            : std_logic;
  SIGNAL Logical_Operator_out7486_out1            : std_logic;
  SIGNAL Logical_Operator_out7487_out1            : std_logic;
  SIGNAL Logical_Operator_out7488_out1            : std_logic;
  SIGNAL Logical_Operator_out7489_out1            : std_logic;
  SIGNAL Logical_Operator_out7490_out1            : std_logic;
  SIGNAL Logical_Operator_out7491_out1            : std_logic;
  SIGNAL Logical_Operator_out7492_out1            : std_logic;
  SIGNAL Logical_Operator_out7493_out1            : std_logic;
  SIGNAL Logical_Operator_out7494_out1            : std_logic;
  SIGNAL Logical_Operator_out7495_out1            : std_logic;
  SIGNAL Logical_Operator_out7496_out1            : std_logic;
  SIGNAL Logical_Operator_out7497_out1            : std_logic;
  SIGNAL Logical_Operator_out7498_out1            : std_logic;
  SIGNAL Logical_Operator_out7499_out1            : std_logic;
  SIGNAL Logical_Operator_out7500_out1            : std_logic;
  SIGNAL Logical_Operator_out7501_out1            : std_logic;
  SIGNAL Logical_Operator_out7502_out1            : std_logic;
  SIGNAL Logical_Operator_out7503_out1            : std_logic;
  SIGNAL Logical_Operator_out7504_out1            : std_logic;
  SIGNAL Logical_Operator_out7505_out1            : std_logic;
  SIGNAL Logical_Operator_out7506_out1            : std_logic;
  SIGNAL Logical_Operator_out7507_out1            : std_logic;
  SIGNAL Logical_Operator_out7508_out1            : std_logic;
  SIGNAL Logical_Operator_out7509_out1            : std_logic;
  SIGNAL Logical_Operator_out7510_out1            : std_logic;
  SIGNAL Logical_Operator_out7511_out1            : std_logic;
  SIGNAL Logical_Operator_out7512_out1            : std_logic;
  SIGNAL Logical_Operator_out7513_out1            : std_logic;
  SIGNAL Logical_Operator_out7514_out1            : std_logic;
  SIGNAL Logical_Operator_out7515_out1            : std_logic;
  SIGNAL Logical_Operator_out7516_out1            : std_logic;
  SIGNAL Logical_Operator_out7517_out1            : std_logic;
  SIGNAL Logical_Operator_out7518_out1            : std_logic;
  SIGNAL Logical_Operator_out7519_out1            : std_logic;
  SIGNAL Logical_Operator_out7520_out1            : std_logic;
  SIGNAL Logical_Operator_out7521_out1            : std_logic;
  SIGNAL Logical_Operator_out7522_out1            : std_logic;
  SIGNAL Logical_Operator_out7523_out1            : std_logic;
  SIGNAL Logical_Operator_out7524_out1            : std_logic;
  SIGNAL Logical_Operator_out7525_out1            : std_logic;
  SIGNAL Logical_Operator_out7526_out1            : std_logic;
  SIGNAL Logical_Operator_out7527_out1            : std_logic;
  SIGNAL Logical_Operator_out7528_out1            : std_logic;
  SIGNAL Logical_Operator_out7529_out1            : std_logic;
  SIGNAL Logical_Operator_out7530_out1            : std_logic;
  SIGNAL Logical_Operator_out7531_out1            : std_logic;
  SIGNAL Logical_Operator_out7532_out1            : std_logic;
  SIGNAL Logical_Operator_out7533_out1            : std_logic;
  SIGNAL Logical_Operator_out7534_out1            : std_logic;
  SIGNAL Logical_Operator_out7535_out1            : std_logic;
  SIGNAL Logical_Operator_out7536_out1            : std_logic;
  SIGNAL Logical_Operator_out7537_out1            : std_logic;
  SIGNAL Logical_Operator_out7538_out1            : std_logic;
  SIGNAL Logical_Operator_out7539_out1            : std_logic;
  SIGNAL Logical_Operator_out7540_out1            : std_logic;
  SIGNAL Logical_Operator_out7541_out1            : std_logic;
  SIGNAL Logical_Operator_out7542_out1            : std_logic;
  SIGNAL Logical_Operator_out7543_out1            : std_logic;
  SIGNAL Logical_Operator_out7544_out1            : std_logic;
  SIGNAL Logical_Operator_out7545_out1            : std_logic;
  SIGNAL Logical_Operator_out7546_out1            : std_logic;
  SIGNAL Logical_Operator_out7547_out1            : std_logic;
  SIGNAL Logical_Operator_out7548_out1            : std_logic;
  SIGNAL Logical_Operator_out7549_out1            : std_logic;
  SIGNAL Logical_Operator_out7550_out1            : std_logic;
  SIGNAL Logical_Operator_out7551_out1            : std_logic;
  SIGNAL Logical_Operator_out7552_out1            : std_logic;
  SIGNAL Logical_Operator_out7553_out1            : std_logic;
  SIGNAL Logical_Operator_out7554_out1            : std_logic;
  SIGNAL Logical_Operator_out7555_out1            : std_logic;
  SIGNAL Logical_Operator_out7556_out1            : std_logic;
  SIGNAL Logical_Operator_out7557_out1            : std_logic;
  SIGNAL Logical_Operator_out7558_out1            : std_logic;
  SIGNAL Logical_Operator_out7559_out1            : std_logic;
  SIGNAL Logical_Operator_out7560_out1            : std_logic;
  SIGNAL Logical_Operator_out7561_out1            : std_logic;
  SIGNAL Logical_Operator_out7562_out1            : std_logic;
  SIGNAL Logical_Operator_out7563_out1            : std_logic;
  SIGNAL Logical_Operator_out7564_out1            : std_logic;
  SIGNAL Logical_Operator_out7565_out1            : std_logic;
  SIGNAL Logical_Operator_out7566_out1            : std_logic;
  SIGNAL Logical_Operator_out7567_out1            : std_logic;
  SIGNAL Logical_Operator_out7568_out1            : std_logic;
  SIGNAL Logical_Operator_out7569_out1            : std_logic;
  SIGNAL Logical_Operator_out7570_out1            : std_logic;
  SIGNAL Logical_Operator_out7571_out1            : std_logic;
  SIGNAL Logical_Operator_out7572_out1            : std_logic;
  SIGNAL Logical_Operator_out7573_out1            : std_logic;
  SIGNAL Logical_Operator_out7574_out1            : std_logic;
  SIGNAL Logical_Operator_out7575_out1            : std_logic;
  SIGNAL Logical_Operator_out7576_out1            : std_logic;
  SIGNAL Logical_Operator_out7577_out1            : std_logic;
  SIGNAL Logical_Operator_out7578_out1            : std_logic;
  SIGNAL Logical_Operator_out7579_out1            : std_logic;
  SIGNAL Logical_Operator_out7580_out1            : std_logic;
  SIGNAL Logical_Operator_out7581_out1            : std_logic;
  SIGNAL Logical_Operator_out7582_out1            : std_logic;
  SIGNAL Logical_Operator_out7583_out1            : std_logic;
  SIGNAL Logical_Operator_out7584_out1            : std_logic;
  SIGNAL Logical_Operator_out7585_out1            : std_logic;
  SIGNAL Logical_Operator_out7586_out1            : std_logic;
  SIGNAL Logical_Operator_out7587_out1            : std_logic;
  SIGNAL Logical_Operator_out7588_out1            : std_logic;
  SIGNAL Logical_Operator_out7589_out1            : std_logic;
  SIGNAL Logical_Operator_out7590_out1            : std_logic;
  SIGNAL Logical_Operator_out7591_out1            : std_logic;
  SIGNAL Logical_Operator_out7592_out1            : std_logic;
  SIGNAL Logical_Operator_out7593_out1            : std_logic;
  SIGNAL Logical_Operator_out7594_out1            : std_logic;
  SIGNAL Logical_Operator_out7595_out1            : std_logic;
  SIGNAL Logical_Operator_out7596_out1            : std_logic;
  SIGNAL Logical_Operator_out7597_out1            : std_logic;
  SIGNAL Logical_Operator_out7598_out1            : std_logic;
  SIGNAL Logical_Operator_out7599_out1            : std_logic;
  SIGNAL Logical_Operator_out7600_out1            : std_logic;
  SIGNAL Logical_Operator_out7601_out1            : std_logic;
  SIGNAL Logical_Operator_out7602_out1            : std_logic;
  SIGNAL Logical_Operator_out7603_out1            : std_logic;
  SIGNAL Logical_Operator_out7604_out1            : std_logic;
  SIGNAL Logical_Operator_out7605_out1            : std_logic;
  SIGNAL Logical_Operator_out7606_out1            : std_logic;
  SIGNAL Logical_Operator_out7607_out1            : std_logic;
  SIGNAL Logical_Operator_out7608_out1            : std_logic;
  SIGNAL Logical_Operator_out7609_out1            : std_logic;
  SIGNAL Logical_Operator_out7610_out1            : std_logic;
  SIGNAL Logical_Operator_out7611_out1            : std_logic;
  SIGNAL Logical_Operator_out7612_out1            : std_logic;
  SIGNAL Logical_Operator_out7613_out1            : std_logic;
  SIGNAL Logical_Operator_out7614_out1            : std_logic;
  SIGNAL Logical_Operator_out7615_out1            : std_logic;
  SIGNAL Logical_Operator_out7616_out1            : std_logic;
  SIGNAL Logical_Operator_out7617_out1            : std_logic;
  SIGNAL Logical_Operator_out7618_out1            : std_logic;
  SIGNAL Logical_Operator_out7619_out1            : std_logic;
  SIGNAL Logical_Operator_out7620_out1            : std_logic;
  SIGNAL Logical_Operator_out7621_out1            : std_logic;
  SIGNAL Logical_Operator_out7622_out1            : std_logic;
  SIGNAL Logical_Operator_out7623_out1            : std_logic;
  SIGNAL Logical_Operator_out7624_out1            : std_logic;
  SIGNAL Logical_Operator_out7625_out1            : std_logic;
  SIGNAL Logical_Operator_out7626_out1            : std_logic;
  SIGNAL Logical_Operator_out7627_out1            : std_logic;
  SIGNAL Logical_Operator_out7628_out1            : std_logic;
  SIGNAL Logical_Operator_out7629_out1            : std_logic;
  SIGNAL Logical_Operator_out7630_out1            : std_logic;
  SIGNAL Logical_Operator_out7631_out1            : std_logic;
  SIGNAL Logical_Operator_out7632_out1            : std_logic;
  SIGNAL Logical_Operator_out7633_out1            : std_logic;
  SIGNAL Logical_Operator_out7634_out1            : std_logic;
  SIGNAL Logical_Operator_out7635_out1            : std_logic;
  SIGNAL Logical_Operator_out7636_out1            : std_logic;
  SIGNAL Logical_Operator_out7637_out1            : std_logic;
  SIGNAL Logical_Operator_out7638_out1            : std_logic;
  SIGNAL Logical_Operator_out7639_out1            : std_logic;
  SIGNAL Logical_Operator_out7640_out1            : std_logic;
  SIGNAL Logical_Operator_out7641_out1            : std_logic;
  SIGNAL Logical_Operator_out7642_out1            : std_logic;
  SIGNAL Logical_Operator_out7643_out1            : std_logic;
  SIGNAL Logical_Operator_out7644_out1            : std_logic;
  SIGNAL Logical_Operator_out7645_out1            : std_logic;
  SIGNAL Logical_Operator_out7646_out1            : std_logic;
  SIGNAL Logical_Operator_out7647_out1            : std_logic;
  SIGNAL Logical_Operator_out7648_out1            : std_logic;
  SIGNAL Logical_Operator_out7649_out1            : std_logic;
  SIGNAL Logical_Operator_out7650_out1            : std_logic;
  SIGNAL Logical_Operator_out7651_out1            : std_logic;
  SIGNAL Logical_Operator_out7652_out1            : std_logic;
  SIGNAL Logical_Operator_out7653_out1            : std_logic;
  SIGNAL Logical_Operator_out7654_out1            : std_logic;
  SIGNAL Logical_Operator_out7655_out1            : std_logic;
  SIGNAL Logical_Operator_out7656_out1            : std_logic;
  SIGNAL Logical_Operator_out7657_out1            : std_logic;
  SIGNAL Logical_Operator_out7658_out1            : std_logic;
  SIGNAL Logical_Operator_out7659_out1            : std_logic;
  SIGNAL Logical_Operator_out7660_out1            : std_logic;
  SIGNAL Logical_Operator_out7661_out1            : std_logic;
  SIGNAL Logical_Operator_out7662_out1            : std_logic;
  SIGNAL Logical_Operator_out7663_out1            : std_logic;
  SIGNAL Logical_Operator_out7664_out1            : std_logic;
  SIGNAL Logical_Operator_out7665_out1            : std_logic;
  SIGNAL Logical_Operator_out7666_out1            : std_logic;
  SIGNAL Logical_Operator_out7667_out1            : std_logic;
  SIGNAL Logical_Operator_out7668_out1            : std_logic;
  SIGNAL Logical_Operator_out7669_out1            : std_logic;
  SIGNAL Logical_Operator_out7670_out1            : std_logic;
  SIGNAL Logical_Operator_out7671_out1            : std_logic;
  SIGNAL Logical_Operator_out7672_out1            : std_logic;
  SIGNAL Logical_Operator_out7673_out1            : std_logic;
  SIGNAL Logical_Operator_out7674_out1            : std_logic;
  SIGNAL Logical_Operator_out7675_out1            : std_logic;
  SIGNAL Logical_Operator_out7676_out1            : std_logic;
  SIGNAL Logical_Operator_out7677_out1            : std_logic;
  SIGNAL Logical_Operator_out7678_out1            : std_logic;
  SIGNAL Logical_Operator_out7679_out1            : std_logic;
  SIGNAL Logical_Operator_out7680_out1            : std_logic;
  SIGNAL Logical_Operator_out7681_out1            : std_logic;
  SIGNAL Logical_Operator_out7682_out1            : std_logic;
  SIGNAL Logical_Operator_out7683_out1            : std_logic;
  SIGNAL Logical_Operator_out7684_out1            : std_logic;
  SIGNAL Logical_Operator_out7685_out1            : std_logic;
  SIGNAL Logical_Operator_out7686_out1            : std_logic;
  SIGNAL Logical_Operator_out7687_out1            : std_logic;
  SIGNAL Logical_Operator_out7688_out1            : std_logic;
  SIGNAL Logical_Operator_out7689_out1            : std_logic;
  SIGNAL Logical_Operator_out7690_out1            : std_logic;
  SIGNAL Logical_Operator_out7691_out1            : std_logic;
  SIGNAL Logical_Operator_out7692_out1            : std_logic;
  SIGNAL Logical_Operator_out7693_out1            : std_logic;
  SIGNAL Logical_Operator_out7694_out1            : std_logic;
  SIGNAL Logical_Operator_out7695_out1            : std_logic;
  SIGNAL Logical_Operator_out7696_out1            : std_logic;
  SIGNAL Logical_Operator_out7697_out1            : std_logic;
  SIGNAL Logical_Operator_out7698_out1            : std_logic;
  SIGNAL Logical_Operator_out7699_out1            : std_logic;
  SIGNAL Logical_Operator_out7700_out1            : std_logic;
  SIGNAL Logical_Operator_out7701_out1            : std_logic;
  SIGNAL Logical_Operator_out7702_out1            : std_logic;
  SIGNAL Logical_Operator_out7703_out1            : std_logic;
  SIGNAL Logical_Operator_out7704_out1            : std_logic;
  SIGNAL Logical_Operator_out7705_out1            : std_logic;
  SIGNAL Logical_Operator_out7706_out1            : std_logic;
  SIGNAL Logical_Operator_out7707_out1            : std_logic;
  SIGNAL Logical_Operator_out7708_out1            : std_logic;
  SIGNAL Logical_Operator_out7709_out1            : std_logic;
  SIGNAL Logical_Operator_out7710_out1            : std_logic;
  SIGNAL Logical_Operator_out7711_out1            : std_logic;
  SIGNAL Logical_Operator_out7712_out1            : std_logic;
  SIGNAL Logical_Operator_out7713_out1            : std_logic;
  SIGNAL Logical_Operator_out7714_out1            : std_logic;
  SIGNAL Logical_Operator_out7715_out1            : std_logic;
  SIGNAL Logical_Operator_out7716_out1            : std_logic;
  SIGNAL Logical_Operator_out7717_out1            : std_logic;
  SIGNAL Logical_Operator_out7718_out1            : std_logic;
  SIGNAL Logical_Operator_out7719_out1            : std_logic;
  SIGNAL Logical_Operator_out7720_out1            : std_logic;
  SIGNAL Logical_Operator_out7721_out1            : std_logic;
  SIGNAL Logical_Operator_out7722_out1            : std_logic;
  SIGNAL Logical_Operator_out7723_out1            : std_logic;
  SIGNAL Logical_Operator_out7724_out1            : std_logic;
  SIGNAL Logical_Operator_out7725_out1            : std_logic;
  SIGNAL Logical_Operator_out7726_out1            : std_logic;
  SIGNAL Logical_Operator_out7727_out1            : std_logic;
  SIGNAL Logical_Operator_out7728_out1            : std_logic;
  SIGNAL Logical_Operator_out7729_out1            : std_logic;
  SIGNAL Logical_Operator_out7730_out1            : std_logic;
  SIGNAL Logical_Operator_out7731_out1            : std_logic;
  SIGNAL Logical_Operator_out7732_out1            : std_logic;
  SIGNAL Logical_Operator_out7733_out1            : std_logic;
  SIGNAL Logical_Operator_out7734_out1            : std_logic;
  SIGNAL Logical_Operator_out7735_out1            : std_logic;
  SIGNAL Logical_Operator_out7736_out1            : std_logic;
  SIGNAL Logical_Operator_out7737_out1            : std_logic;
  SIGNAL Logical_Operator_out7738_out1            : std_logic;
  SIGNAL Logical_Operator_out7739_out1            : std_logic;
  SIGNAL Logical_Operator_out7740_out1            : std_logic;
  SIGNAL Logical_Operator_out7741_out1            : std_logic;
  SIGNAL Logical_Operator_out7742_out1            : std_logic;
  SIGNAL Logical_Operator_out7743_out1            : std_logic;
  SIGNAL Logical_Operator_out7744_out1            : std_logic;
  SIGNAL Logical_Operator_out7745_out1            : std_logic;
  SIGNAL Logical_Operator_out7746_out1            : std_logic;
  SIGNAL Logical_Operator_out7747_out1            : std_logic;
  SIGNAL Logical_Operator_out7748_out1            : std_logic;
  SIGNAL Logical_Operator_out7749_out1            : std_logic;
  SIGNAL Logical_Operator_out7750_out1            : std_logic;
  SIGNAL Logical_Operator_out7751_out1            : std_logic;
  SIGNAL Logical_Operator_out7752_out1            : std_logic;
  SIGNAL Logical_Operator_out7753_out1            : std_logic;
  SIGNAL Logical_Operator_out7754_out1            : std_logic;
  SIGNAL Logical_Operator_out7755_out1            : std_logic;
  SIGNAL Logical_Operator_out7756_out1            : std_logic;
  SIGNAL Logical_Operator_out7757_out1            : std_logic;
  SIGNAL Logical_Operator_out7758_out1            : std_logic;
  SIGNAL Logical_Operator_out7759_out1            : std_logic;
  SIGNAL Logical_Operator_out7760_out1            : std_logic;
  SIGNAL Logical_Operator_out7761_out1            : std_logic;
  SIGNAL Logical_Operator_out7762_out1            : std_logic;
  SIGNAL Logical_Operator_out7763_out1            : std_logic;
  SIGNAL Logical_Operator_out7764_out1            : std_logic;
  SIGNAL Logical_Operator_out7765_out1            : std_logic;
  SIGNAL Logical_Operator_out7766_out1            : std_logic;
  SIGNAL Logical_Operator_out7767_out1            : std_logic;
  SIGNAL Logical_Operator_out7768_out1            : std_logic;
  SIGNAL Logical_Operator_out7769_out1            : std_logic;
  SIGNAL Logical_Operator_out7770_out1            : std_logic;
  SIGNAL Logical_Operator_out7771_out1            : std_logic;
  SIGNAL Logical_Operator_out7772_out1            : std_logic;
  SIGNAL Logical_Operator_out7773_out1            : std_logic;
  SIGNAL Logical_Operator_out7774_out1            : std_logic;
  SIGNAL Logical_Operator_out7775_out1            : std_logic;
  SIGNAL Logical_Operator_out7776_out1            : std_logic;
  SIGNAL Logical_Operator_out7777_out1            : std_logic;
  SIGNAL Logical_Operator_out7778_out1            : std_logic;
  SIGNAL Logical_Operator_out7779_out1            : std_logic;
  SIGNAL Logical_Operator_out7780_out1            : std_logic;
  SIGNAL Logical_Operator_out7781_out1            : std_logic;
  SIGNAL Logical_Operator_out7782_out1            : std_logic;
  SIGNAL Logical_Operator_out7783_out1            : std_logic;
  SIGNAL Logical_Operator_out7784_out1            : std_logic;
  SIGNAL Logical_Operator_out7785_out1            : std_logic;
  SIGNAL Logical_Operator_out7786_out1            : std_logic;
  SIGNAL Logical_Operator_out7787_out1            : std_logic;
  SIGNAL Logical_Operator_out7788_out1            : std_logic;
  SIGNAL Logical_Operator_out7789_out1            : std_logic;
  SIGNAL Logical_Operator_out7790_out1            : std_logic;
  SIGNAL Logical_Operator_out7791_out1            : std_logic;
  SIGNAL Logical_Operator_out7792_out1            : std_logic;
  SIGNAL Logical_Operator_out7793_out1            : std_logic;
  SIGNAL Logical_Operator_out7794_out1            : std_logic;
  SIGNAL Logical_Operator_out7795_out1            : std_logic;
  SIGNAL Logical_Operator_out7796_out1            : std_logic;
  SIGNAL Logical_Operator_out7797_out1            : std_logic;
  SIGNAL Logical_Operator_out7798_out1            : std_logic;
  SIGNAL Logical_Operator_out7799_out1            : std_logic;
  SIGNAL Logical_Operator_out7800_out1            : std_logic;
  SIGNAL Logical_Operator_out7801_out1            : std_logic;
  SIGNAL Logical_Operator_out7802_out1            : std_logic;
  SIGNAL Logical_Operator_out7803_out1            : std_logic;
  SIGNAL Logical_Operator_out7804_out1            : std_logic;
  SIGNAL Logical_Operator_out7805_out1            : std_logic;
  SIGNAL Logical_Operator_out7806_out1            : std_logic;
  SIGNAL Logical_Operator_out7807_out1            : std_logic;
  SIGNAL Logical_Operator_out7808_out1            : std_logic;
  SIGNAL Logical_Operator_out7809_out1            : std_logic;
  SIGNAL Logical_Operator_out7810_out1            : std_logic;
  SIGNAL Logical_Operator_out7811_out1            : std_logic;
  SIGNAL Logical_Operator_out7812_out1            : std_logic;
  SIGNAL Logical_Operator_out7813_out1            : std_logic;
  SIGNAL Logical_Operator_out7814_out1            : std_logic;
  SIGNAL Logical_Operator_out7815_out1            : std_logic;
  SIGNAL Logical_Operator_out7816_out1            : std_logic;
  SIGNAL Logical_Operator_out7817_out1            : std_logic;
  SIGNAL Logical_Operator_out7818_out1            : std_logic;
  SIGNAL Logical_Operator_out7819_out1            : std_logic;
  SIGNAL Logical_Operator_out7820_out1            : std_logic;
  SIGNAL Logical_Operator_out7821_out1            : std_logic;
  SIGNAL Logical_Operator_out7822_out1            : std_logic;
  SIGNAL Logical_Operator_out7823_out1            : std_logic;
  SIGNAL Logical_Operator_out7824_out1            : std_logic;
  SIGNAL Logical_Operator_out7825_out1            : std_logic;
  SIGNAL Logical_Operator_out7826_out1            : std_logic;
  SIGNAL Logical_Operator_out7827_out1            : std_logic;
  SIGNAL Logical_Operator_out7828_out1            : std_logic;
  SIGNAL Logical_Operator_out7829_out1            : std_logic;
  SIGNAL Logical_Operator_out7830_out1            : std_logic;
  SIGNAL Logical_Operator_out7831_out1            : std_logic;
  SIGNAL Logical_Operator_out7832_out1            : std_logic;
  SIGNAL Logical_Operator_out7833_out1            : std_logic;
  SIGNAL Logical_Operator_out7834_out1            : std_logic;
  SIGNAL Logical_Operator_out7835_out1            : std_logic;
  SIGNAL Logical_Operator_out7836_out1            : std_logic;
  SIGNAL Logical_Operator_out7837_out1            : std_logic;
  SIGNAL Logical_Operator_out7838_out1            : std_logic;
  SIGNAL Logical_Operator_out7839_out1            : std_logic;
  SIGNAL Logical_Operator_out7840_out1            : std_logic;
  SIGNAL Logical_Operator_out7841_out1            : std_logic;
  SIGNAL Logical_Operator_out7842_out1            : std_logic;
  SIGNAL Logical_Operator_out7843_out1            : std_logic;
  SIGNAL Logical_Operator_out7844_out1            : std_logic;
  SIGNAL Logical_Operator_out7845_out1            : std_logic;
  SIGNAL Logical_Operator_out7846_out1            : std_logic;
  SIGNAL Logical_Operator_out7847_out1            : std_logic;
  SIGNAL Logical_Operator_out7848_out1            : std_logic;
  SIGNAL Logical_Operator_out7849_out1            : std_logic;
  SIGNAL Logical_Operator_out7850_out1            : std_logic;
  SIGNAL Logical_Operator_out7851_out1            : std_logic;
  SIGNAL Logical_Operator_out7852_out1            : std_logic;
  SIGNAL Logical_Operator_out7853_out1            : std_logic;
  SIGNAL Logical_Operator_out7854_out1            : std_logic;
  SIGNAL Logical_Operator_out7855_out1            : std_logic;
  SIGNAL Logical_Operator_out7856_out1            : std_logic;
  SIGNAL Logical_Operator_out7857_out1            : std_logic;
  SIGNAL Logical_Operator_out7858_out1            : std_logic;
  SIGNAL Logical_Operator_out7859_out1            : std_logic;
  SIGNAL Logical_Operator_out7860_out1            : std_logic;
  SIGNAL Logical_Operator_out7861_out1            : std_logic;
  SIGNAL Logical_Operator_out7862_out1            : std_logic;
  SIGNAL Logical_Operator_out7863_out1            : std_logic;
  SIGNAL Logical_Operator_out7864_out1            : std_logic;
  SIGNAL Logical_Operator_out7865_out1            : std_logic;
  SIGNAL Logical_Operator_out7866_out1            : std_logic;
  SIGNAL Logical_Operator_out7867_out1            : std_logic;
  SIGNAL Logical_Operator_out7868_out1            : std_logic;
  SIGNAL Logical_Operator_out7869_out1            : std_logic;
  SIGNAL Logical_Operator_out7870_out1            : std_logic;
  SIGNAL Logical_Operator_out7871_out1            : std_logic;
  SIGNAL Logical_Operator_out7872_out1            : std_logic;
  SIGNAL Logical_Operator_out7873_out1            : std_logic;
  SIGNAL Logical_Operator_out7874_out1            : std_logic;
  SIGNAL Logical_Operator_out7875_out1            : std_logic;
  SIGNAL Logical_Operator_out7876_out1            : std_logic;
  SIGNAL Logical_Operator_out7877_out1            : std_logic;
  SIGNAL Logical_Operator_out7878_out1            : std_logic;
  SIGNAL Logical_Operator_out7879_out1            : std_logic;
  SIGNAL Logical_Operator_out7880_out1            : std_logic;
  SIGNAL Logical_Operator_out7881_out1            : std_logic;
  SIGNAL Logical_Operator_out7882_out1            : std_logic;
  SIGNAL Logical_Operator_out7883_out1            : std_logic;
  SIGNAL Logical_Operator_out7884_out1            : std_logic;
  SIGNAL Logical_Operator_out7885_out1            : std_logic;
  SIGNAL Logical_Operator_out7886_out1            : std_logic;
  SIGNAL Logical_Operator_out7887_out1            : std_logic;
  SIGNAL Logical_Operator_out7888_out1            : std_logic;
  SIGNAL Logical_Operator_out7889_out1            : std_logic;
  SIGNAL Logical_Operator_out7890_out1            : std_logic;
  SIGNAL Logical_Operator_out7891_out1            : std_logic;
  SIGNAL Logical_Operator_out7892_out1            : std_logic;
  SIGNAL Logical_Operator_out7893_out1            : std_logic;
  SIGNAL Logical_Operator_out7894_out1            : std_logic;
  SIGNAL Logical_Operator_out7895_out1            : std_logic;
  SIGNAL Logical_Operator_out7896_out1            : std_logic;
  SIGNAL Logical_Operator_out7897_out1            : std_logic;
  SIGNAL Logical_Operator_out7898_out1            : std_logic;
  SIGNAL Logical_Operator_out7899_out1            : std_logic;
  SIGNAL Logical_Operator_out7900_out1            : std_logic;
  SIGNAL Logical_Operator_out7901_out1            : std_logic;
  SIGNAL Logical_Operator_out7902_out1            : std_logic;
  SIGNAL Logical_Operator_out7903_out1            : std_logic;
  SIGNAL Logical_Operator_out7904_out1            : std_logic;
  SIGNAL Logical_Operator_out7905_out1            : std_logic;
  SIGNAL Logical_Operator_out7906_out1            : std_logic;
  SIGNAL Logical_Operator_out7907_out1            : std_logic;
  SIGNAL Logical_Operator_out7908_out1            : std_logic;
  SIGNAL Logical_Operator_out7909_out1            : std_logic;
  SIGNAL Logical_Operator_out7910_out1            : std_logic;
  SIGNAL Logical_Operator_out7911_out1            : std_logic;
  SIGNAL Logical_Operator_out7912_out1            : std_logic;
  SIGNAL Logical_Operator_out7913_out1            : std_logic;
  SIGNAL Logical_Operator_out7914_out1            : std_logic;
  SIGNAL Logical_Operator_out7915_out1            : std_logic;
  SIGNAL Logical_Operator_out7916_out1            : std_logic;
  SIGNAL Logical_Operator_out7917_out1            : std_logic;
  SIGNAL Logical_Operator_out7918_out1            : std_logic;
  SIGNAL Logical_Operator_out7919_out1            : std_logic;
  SIGNAL Logical_Operator_out7920_out1            : std_logic;
  SIGNAL Logical_Operator_out7921_out1            : std_logic;
  SIGNAL Logical_Operator_out7922_out1            : std_logic;
  SIGNAL Logical_Operator_out7923_out1            : std_logic;
  SIGNAL Logical_Operator_out7924_out1            : std_logic;
  SIGNAL Logical_Operator_out7925_out1            : std_logic;
  SIGNAL Logical_Operator_out7926_out1            : std_logic;
  SIGNAL Logical_Operator_out7927_out1            : std_logic;
  SIGNAL Logical_Operator_out7928_out1            : std_logic;
  SIGNAL Logical_Operator_out7929_out1            : std_logic;
  SIGNAL Logical_Operator_out7930_out1            : std_logic;
  SIGNAL Logical_Operator_out7931_out1            : std_logic;
  SIGNAL Logical_Operator_out7932_out1            : std_logic;
  SIGNAL Logical_Operator_out7933_out1            : std_logic;
  SIGNAL Logical_Operator_out7934_out1            : std_logic;
  SIGNAL Logical_Operator_out7935_out1            : std_logic;
  SIGNAL Logical_Operator_out7936_out1            : std_logic;
  SIGNAL Logical_Operator_out7937_out1            : std_logic;
  SIGNAL Logical_Operator_out7938_out1            : std_logic;
  SIGNAL Logical_Operator_out7939_out1            : std_logic;
  SIGNAL Logical_Operator_out7940_out1            : std_logic;
  SIGNAL Logical_Operator_out7941_out1            : std_logic;
  SIGNAL Logical_Operator_out7942_out1            : std_logic;
  SIGNAL Logical_Operator_out7943_out1            : std_logic;
  SIGNAL Logical_Operator_out7944_out1            : std_logic;
  SIGNAL Logical_Operator_out7945_out1            : std_logic;
  SIGNAL Logical_Operator_out7946_out1            : std_logic;
  SIGNAL Logical_Operator_out7947_out1            : std_logic;
  SIGNAL Logical_Operator_out7948_out1            : std_logic;
  SIGNAL Logical_Operator_out7949_out1            : std_logic;
  SIGNAL Logical_Operator_out7950_out1            : std_logic;
  SIGNAL Logical_Operator_out7951_out1            : std_logic;
  SIGNAL Logical_Operator_out7952_out1            : std_logic;
  SIGNAL Logical_Operator_out7953_out1            : std_logic;
  SIGNAL Logical_Operator_out7954_out1            : std_logic;
  SIGNAL Logical_Operator_out7955_out1            : std_logic;
  SIGNAL Logical_Operator_out7956_out1            : std_logic;
  SIGNAL Logical_Operator_out7957_out1            : std_logic;
  SIGNAL Logical_Operator_out7958_out1            : std_logic;
  SIGNAL Logical_Operator_out7959_out1            : std_logic;
  SIGNAL Logical_Operator_out7960_out1            : std_logic;
  SIGNAL Logical_Operator_out7961_out1            : std_logic;
  SIGNAL Logical_Operator_out7962_out1            : std_logic;
  SIGNAL Logical_Operator_out7963_out1            : std_logic;
  SIGNAL Logical_Operator_out7964_out1            : std_logic;
  SIGNAL Logical_Operator_out7965_out1            : std_logic;
  SIGNAL Logical_Operator_out7966_out1            : std_logic;
  SIGNAL Logical_Operator_out7967_out1            : std_logic;
  SIGNAL Logical_Operator_out7968_out1            : std_logic;
  SIGNAL Logical_Operator_out7969_out1            : std_logic;
  SIGNAL Logical_Operator_out7970_out1            : std_logic;
  SIGNAL Logical_Operator_out7971_out1            : std_logic;
  SIGNAL Logical_Operator_out7972_out1            : std_logic;
  SIGNAL Logical_Operator_out7973_out1            : std_logic;
  SIGNAL Logical_Operator_out7974_out1            : std_logic;
  SIGNAL Logical_Operator_out7975_out1            : std_logic;
  SIGNAL Logical_Operator_out7976_out1            : std_logic;
  SIGNAL Logical_Operator_out7977_out1            : std_logic;
  SIGNAL Logical_Operator_out7978_out1            : std_logic;
  SIGNAL Logical_Operator_out7979_out1            : std_logic;
  SIGNAL Logical_Operator_out7980_out1            : std_logic;
  SIGNAL Logical_Operator_out7981_out1            : std_logic;
  SIGNAL Logical_Operator_out7982_out1            : std_logic;
  SIGNAL Logical_Operator_out7983_out1            : std_logic;
  SIGNAL Logical_Operator_out7984_out1            : std_logic;
  SIGNAL Logical_Operator_out7985_out1            : std_logic;
  SIGNAL Logical_Operator_out7986_out1            : std_logic;
  SIGNAL Logical_Operator_out7987_out1            : std_logic;
  SIGNAL Logical_Operator_out7988_out1            : std_logic;
  SIGNAL Logical_Operator_out7989_out1            : std_logic;
  SIGNAL Logical_Operator_out7990_out1            : std_logic;
  SIGNAL Logical_Operator_out7991_out1            : std_logic;
  SIGNAL Logical_Operator_out7992_out1            : std_logic;
  SIGNAL Logical_Operator_out7993_out1            : std_logic;
  SIGNAL Logical_Operator_out7994_out1            : std_logic;
  SIGNAL Logical_Operator_out7995_out1            : std_logic;
  SIGNAL Logical_Operator_out7996_out1            : std_logic;
  SIGNAL Logical_Operator_out7997_out1            : std_logic;
  SIGNAL Logical_Operator_out7998_out1            : std_logic;
  SIGNAL Logical_Operator_out7999_out1            : std_logic;
  SIGNAL Logical_Operator_out8000_out1            : std_logic;
  SIGNAL Logical_Operator_out8001_out1            : std_logic;
  SIGNAL Logical_Operator_out8002_out1            : std_logic;
  SIGNAL Logical_Operator_out8003_out1            : std_logic;
  SIGNAL Logical_Operator_out8004_out1            : std_logic;
  SIGNAL Logical_Operator_out8005_out1            : std_logic;
  SIGNAL Logical_Operator_out8006_out1            : std_logic;
  SIGNAL Logical_Operator_out8007_out1            : std_logic;
  SIGNAL Logical_Operator_out8008_out1            : std_logic;
  SIGNAL Logical_Operator_out8009_out1            : std_logic;
  SIGNAL Logical_Operator_out8010_out1            : std_logic;
  SIGNAL Logical_Operator_out8011_out1            : std_logic;
  SIGNAL Logical_Operator_out8012_out1            : std_logic;
  SIGNAL Logical_Operator_out8013_out1            : std_logic;
  SIGNAL Logical_Operator_out8014_out1            : std_logic;
  SIGNAL Logical_Operator_out8015_out1            : std_logic;
  SIGNAL Logical_Operator_out8016_out1            : std_logic;
  SIGNAL Logical_Operator_out8017_out1            : std_logic;
  SIGNAL Logical_Operator_out8018_out1            : std_logic;
  SIGNAL Logical_Operator_out8019_out1            : std_logic;
  SIGNAL Logical_Operator_out8020_out1            : std_logic;
  SIGNAL Logical_Operator_out8021_out1            : std_logic;
  SIGNAL Logical_Operator_out8022_out1            : std_logic;
  SIGNAL Logical_Operator_out8023_out1            : std_logic;
  SIGNAL Logical_Operator_out8024_out1            : std_logic;
  SIGNAL Logical_Operator_out8025_out1            : std_logic;
  SIGNAL Logical_Operator_out8026_out1            : std_logic;
  SIGNAL Logical_Operator_out8027_out1            : std_logic;
  SIGNAL Logical_Operator_out8028_out1            : std_logic;
  SIGNAL Logical_Operator_out8029_out1            : std_logic;
  SIGNAL Logical_Operator_out8030_out1            : std_logic;
  SIGNAL Logical_Operator_out8031_out1            : std_logic;
  SIGNAL Logical_Operator_out8032_out1            : std_logic;
  SIGNAL Logical_Operator_out8033_out1            : std_logic;
  SIGNAL Logical_Operator_out8034_out1            : std_logic;
  SIGNAL Logical_Operator_out8035_out1            : std_logic;
  SIGNAL Logical_Operator_out8036_out1            : std_logic;
  SIGNAL Logical_Operator_out8037_out1            : std_logic;
  SIGNAL Logical_Operator_out8038_out1            : std_logic;
  SIGNAL Logical_Operator_out8039_out1            : std_logic;
  SIGNAL Logical_Operator_out8040_out1            : std_logic;
  SIGNAL Logical_Operator_out8041_out1            : std_logic;
  SIGNAL Logical_Operator_out8042_out1            : std_logic;
  SIGNAL Logical_Operator_out8043_out1            : std_logic;
  SIGNAL Logical_Operator_out8044_out1            : std_logic;
  SIGNAL Logical_Operator_out8045_out1            : std_logic;
  SIGNAL Logical_Operator_out8046_out1            : std_logic;
  SIGNAL Logical_Operator_out8047_out1            : std_logic;
  SIGNAL Logical_Operator_out8048_out1            : std_logic;
  SIGNAL Logical_Operator_out8049_out1            : std_logic;
  SIGNAL Logical_Operator_out8050_out1            : std_logic;
  SIGNAL Logical_Operator_out8051_out1            : std_logic;
  SIGNAL Logical_Operator_out8052_out1            : std_logic;
  SIGNAL Logical_Operator_out8053_out1            : std_logic;
  SIGNAL Logical_Operator_out8054_out1            : std_logic;
  SIGNAL Logical_Operator_out8055_out1            : std_logic;
  SIGNAL Logical_Operator_out8056_out1            : std_logic;
  SIGNAL Logical_Operator_out8057_out1            : std_logic;
  SIGNAL Logical_Operator_out8058_out1            : std_logic;
  SIGNAL Logical_Operator_out8059_out1            : std_logic;
  SIGNAL Logical_Operator_out8060_out1            : std_logic;
  SIGNAL Logical_Operator_out8061_out1            : std_logic;
  SIGNAL Logical_Operator_out8062_out1            : std_logic;
  SIGNAL Logical_Operator_out8063_out1            : std_logic;
  SIGNAL Logical_Operator_out8064_out1            : std_logic;
  SIGNAL Logical_Operator_out8065_out1            : std_logic;
  SIGNAL Logical_Operator_out8066_out1            : std_logic;
  SIGNAL Logical_Operator_out8067_out1            : std_logic;
  SIGNAL Logical_Operator_out8068_out1            : std_logic;
  SIGNAL Logical_Operator_out8069_out1            : std_logic;
  SIGNAL Logical_Operator_out8070_out1            : std_logic;
  SIGNAL Logical_Operator_out8071_out1            : std_logic;
  SIGNAL Logical_Operator_out8072_out1            : std_logic;
  SIGNAL Logical_Operator_out8073_out1            : std_logic;
  SIGNAL Logical_Operator_out8074_out1            : std_logic;
  SIGNAL Logical_Operator_out8075_out1            : std_logic;
  SIGNAL Logical_Operator_out8076_out1            : std_logic;
  SIGNAL Logical_Operator_out8077_out1            : std_logic;
  SIGNAL Logical_Operator_out8078_out1            : std_logic;
  SIGNAL Logical_Operator_out8079_out1            : std_logic;
  SIGNAL Logical_Operator_out8080_out1            : std_logic;
  SIGNAL Logical_Operator_out8081_out1            : std_logic;
  SIGNAL Logical_Operator_out8082_out1            : std_logic;
  SIGNAL Logical_Operator_out8083_out1            : std_logic;
  SIGNAL Logical_Operator_out8084_out1            : std_logic;
  SIGNAL Logical_Operator_out8085_out1            : std_logic;
  SIGNAL Logical_Operator_out8086_out1            : std_logic;
  SIGNAL Logical_Operator_out8087_out1            : std_logic;
  SIGNAL Logical_Operator_out8088_out1            : std_logic;
  SIGNAL Logical_Operator_out8089_out1            : std_logic;
  SIGNAL Logical_Operator_out8090_out1            : std_logic;
  SIGNAL Logical_Operator_out8091_out1            : std_logic;
  SIGNAL Logical_Operator_out8092_out1            : std_logic;
  SIGNAL Logical_Operator_out8093_out1            : std_logic;
  SIGNAL Logical_Operator_out8094_out1            : std_logic;
  SIGNAL Logical_Operator_out8095_out1            : std_logic;
  SIGNAL Logical_Operator_out8096_out1            : std_logic;
  SIGNAL Logical_Operator_out8097_out1            : std_logic;
  SIGNAL Logical_Operator_out8098_out1            : std_logic;
  SIGNAL Logical_Operator_out8099_out1            : std_logic;
  SIGNAL Logical_Operator_out8100_out1            : std_logic;
  SIGNAL Logical_Operator_out8101_out1            : std_logic;
  SIGNAL Logical_Operator_out8102_out1            : std_logic;
  SIGNAL Logical_Operator_out8103_out1            : std_logic;
  SIGNAL Logical_Operator_out8104_out1            : std_logic;
  SIGNAL Logical_Operator_out8105_out1            : std_logic;
  SIGNAL Logical_Operator_out8106_out1            : std_logic;
  SIGNAL Logical_Operator_out8107_out1            : std_logic;
  SIGNAL Logical_Operator_out8108_out1            : std_logic;
  SIGNAL Logical_Operator_out8109_out1            : std_logic;
  SIGNAL Logical_Operator_out8110_out1            : std_logic;
  SIGNAL Logical_Operator_out8111_out1            : std_logic;
  SIGNAL Logical_Operator_out8112_out1            : std_logic;
  SIGNAL Logical_Operator_out8113_out1            : std_logic;
  SIGNAL Logical_Operator_out8114_out1            : std_logic;
  SIGNAL Logical_Operator_out8115_out1            : std_logic;
  SIGNAL Logical_Operator_out8116_out1            : std_logic;
  SIGNAL Logical_Operator_out8117_out1            : std_logic;
  SIGNAL Logical_Operator_out8118_out1            : std_logic;
  SIGNAL Logical_Operator_out8119_out1            : std_logic;
  SIGNAL Logical_Operator_out8120_out1            : std_logic;
  SIGNAL Logical_Operator_out8121_out1            : std_logic;
  SIGNAL Logical_Operator_out8122_out1            : std_logic;
  SIGNAL Logical_Operator_out8123_out1            : std_logic;
  SIGNAL Logical_Operator_out8124_out1            : std_logic;
  SIGNAL Logical_Operator_out8125_out1            : std_logic;
  SIGNAL Logical_Operator_out8126_out1            : std_logic;
  SIGNAL Logical_Operator_out8127_out1            : std_logic;
  SIGNAL Logical_Operator_out8128_out1            : std_logic;
  SIGNAL Logical_Operator_out8129_out1            : std_logic;
  SIGNAL Logical_Operator_out8130_out1            : std_logic;
  SIGNAL Logical_Operator_out8131_out1            : std_logic;
  SIGNAL Logical_Operator_out8132_out1            : std_logic;
  SIGNAL Logical_Operator_out8133_out1            : std_logic;
  SIGNAL Logical_Operator_out8134_out1            : std_logic;
  SIGNAL Logical_Operator_out8135_out1            : std_logic;
  SIGNAL Logical_Operator_out8136_out1            : std_logic;
  SIGNAL Logical_Operator_out8137_out1            : std_logic;
  SIGNAL Logical_Operator_out8138_out1            : std_logic;
  SIGNAL Logical_Operator_out8139_out1            : std_logic;
  SIGNAL Logical_Operator_out8140_out1            : std_logic;
  SIGNAL Logical_Operator_out8141_out1            : std_logic;
  SIGNAL Logical_Operator_out8142_out1            : std_logic;
  SIGNAL Logical_Operator_out8143_out1            : std_logic;
  SIGNAL Logical_Operator_out8144_out1            : std_logic;
  SIGNAL Logical_Operator_out8145_out1            : std_logic;
  SIGNAL Logical_Operator_out8146_out1            : std_logic;
  SIGNAL Logical_Operator_out8147_out1            : std_logic;
  SIGNAL Logical_Operator_out8148_out1            : std_logic;
  SIGNAL Logical_Operator_out8149_out1            : std_logic;
  SIGNAL Logical_Operator_out8150_out1            : std_logic;
  SIGNAL Logical_Operator_out8151_out1            : std_logic;
  SIGNAL Logical_Operator_out8152_out1            : std_logic;
  SIGNAL Logical_Operator_out8153_out1            : std_logic;
  SIGNAL Logical_Operator_out8154_out1            : std_logic;
  SIGNAL Logical_Operator_out8155_out1            : std_logic;
  SIGNAL Logical_Operator_out8156_out1            : std_logic;
  SIGNAL Logical_Operator_out8157_out1            : std_logic;
  SIGNAL Logical_Operator_out8158_out1            : std_logic;
  SIGNAL Logical_Operator_out8159_out1            : std_logic;
  SIGNAL Logical_Operator_out8160_out1            : std_logic;
  SIGNAL Logical_Operator_out8161_out1            : std_logic;
  SIGNAL Logical_Operator_out8162_out1            : std_logic;
  SIGNAL Logical_Operator_out8163_out1            : std_logic;
  SIGNAL Logical_Operator_out8164_out1            : std_logic;
  SIGNAL Logical_Operator_out8165_out1            : std_logic;
  SIGNAL Logical_Operator_out8166_out1            : std_logic;
  SIGNAL Logical_Operator_out8167_out1            : std_logic;
  SIGNAL Logical_Operator_out8168_out1            : std_logic;
  SIGNAL Logical_Operator_out8169_out1            : std_logic;
  SIGNAL Logical_Operator_out8170_out1            : std_logic;
  SIGNAL Logical_Operator_out8171_out1            : std_logic;
  SIGNAL Logical_Operator_out8172_out1            : std_logic;
  SIGNAL Logical_Operator_out8173_out1            : std_logic;
  SIGNAL Logical_Operator_out8174_out1            : std_logic;
  SIGNAL Logical_Operator_out8175_out1            : std_logic;
  SIGNAL Logical_Operator_out8176_out1            : std_logic;
  SIGNAL Logical_Operator_out8177_out1            : std_logic;
  SIGNAL Logical_Operator_out8178_out1            : std_logic;
  SIGNAL Logical_Operator_out8179_out1            : std_logic;
  SIGNAL Logical_Operator_out8180_out1            : std_logic;
  SIGNAL Logical_Operator_out8181_out1            : std_logic;
  SIGNAL Logical_Operator_out8182_out1            : std_logic;
  SIGNAL Logical_Operator_out8183_out1            : std_logic;
  SIGNAL Logical_Operator_out8184_out1            : std_logic;
  SIGNAL Logical_Operator_out8185_out1            : std_logic;
  SIGNAL Logical_Operator_out8186_out1            : std_logic;
  SIGNAL Logical_Operator_out8187_out1            : std_logic;
  SIGNAL Logical_Operator_out8188_out1            : std_logic;
  SIGNAL Logical_Operator_out8189_out1            : std_logic;
  SIGNAL Logical_Operator_out8190_out1            : std_logic;
  SIGNAL Logical_Operator_out8191_out1            : std_logic;
  SIGNAL Logical_Operator_out8192_out1            : std_logic;
  SIGNAL Logical_Operator_out8193_out1            : std_logic;
  SIGNAL Logical_Operator_out8194_out1            : std_logic;
  SIGNAL Logical_Operator_out8195_out1            : std_logic;
  SIGNAL Logical_Operator_out8196_out1            : std_logic;
  SIGNAL Logical_Operator_out8197_out1            : std_logic;
  SIGNAL Logical_Operator_out8198_out1            : std_logic;
  SIGNAL Logical_Operator_out8199_out1            : std_logic;
  SIGNAL Logical_Operator_out8200_out1            : std_logic;
  SIGNAL Logical_Operator_out8201_out1            : std_logic;
  SIGNAL Logical_Operator_out8202_out1            : std_logic;
  SIGNAL Logical_Operator_out8203_out1            : std_logic;
  SIGNAL Logical_Operator_out8204_out1            : std_logic;
  SIGNAL Logical_Operator_out8205_out1            : std_logic;
  SIGNAL Logical_Operator_out8206_out1            : std_logic;
  SIGNAL Logical_Operator_out8207_out1            : std_logic;
  SIGNAL Logical_Operator_out8208_out1            : std_logic;
  SIGNAL Logical_Operator_out8209_out1            : std_logic;
  SIGNAL Logical_Operator_out8210_out1            : std_logic;
  SIGNAL Logical_Operator_out8211_out1            : std_logic;
  SIGNAL Logical_Operator_out8212_out1            : std_logic;
  SIGNAL Logical_Operator_out8213_out1            : std_logic;
  SIGNAL Logical_Operator_out8214_out1            : std_logic;
  SIGNAL Logical_Operator_out8215_out1            : std_logic;
  SIGNAL Logical_Operator_out8216_out1            : std_logic;
  SIGNAL Logical_Operator_out8217_out1            : std_logic;
  SIGNAL Logical_Operator_out8218_out1            : std_logic;
  SIGNAL Logical_Operator_out8219_out1            : std_logic;
  SIGNAL Logical_Operator_out8220_out1            : std_logic;
  SIGNAL Logical_Operator_out8221_out1            : std_logic;
  SIGNAL Logical_Operator_out8222_out1            : std_logic;
  SIGNAL Logical_Operator_out8223_out1            : std_logic;
  SIGNAL Logical_Operator_out8224_out1            : std_logic;
  SIGNAL Logical_Operator_out8225_out1            : std_logic;
  SIGNAL Logical_Operator_out8226_out1            : std_logic;
  SIGNAL Logical_Operator_out8227_out1            : std_logic;
  SIGNAL Logical_Operator_out8228_out1            : std_logic;
  SIGNAL Logical_Operator_out8229_out1            : std_logic;
  SIGNAL Logical_Operator_out8230_out1            : std_logic;
  SIGNAL Logical_Operator_out8231_out1            : std_logic;
  SIGNAL Logical_Operator_out8232_out1            : std_logic;
  SIGNAL Logical_Operator_out8233_out1            : std_logic;
  SIGNAL Logical_Operator_out8234_out1            : std_logic;
  SIGNAL Logical_Operator_out8235_out1            : std_logic;
  SIGNAL Logical_Operator_out8236_out1            : std_logic;
  SIGNAL Logical_Operator_out8237_out1            : std_logic;
  SIGNAL Logical_Operator_out8238_out1            : std_logic;
  SIGNAL Logical_Operator_out8239_out1            : std_logic;
  SIGNAL Logical_Operator_out8240_out1            : std_logic;
  SIGNAL Logical_Operator_out8241_out1            : std_logic;
  SIGNAL Logical_Operator_out8242_out1            : std_logic;
  SIGNAL Logical_Operator_out8243_out1            : std_logic;
  SIGNAL Logical_Operator_out8244_out1            : std_logic;
  SIGNAL Logical_Operator_out8245_out1            : std_logic;
  SIGNAL Logical_Operator_out8246_out1            : std_logic;
  SIGNAL Logical_Operator_out8247_out1            : std_logic;
  SIGNAL Logical_Operator_out8248_out1            : std_logic;
  SIGNAL Logical_Operator_out8249_out1            : std_logic;
  SIGNAL Logical_Operator_out8250_out1            : std_logic;
  SIGNAL Logical_Operator_out8251_out1            : std_logic;
  SIGNAL Logical_Operator_out8252_out1            : std_logic;
  SIGNAL Logical_Operator_out8253_out1            : std_logic;
  SIGNAL Logical_Operator_out8254_out1            : std_logic;
  SIGNAL Logical_Operator_out8255_out1            : std_logic;
  SIGNAL Logical_Operator_out8256_out1            : std_logic;
  SIGNAL Logical_Operator_out8257_out1            : std_logic;
  SIGNAL Logical_Operator_out8258_out1            : std_logic;
  SIGNAL Logical_Operator_out8259_out1            : std_logic;
  SIGNAL Logical_Operator_out8260_out1            : std_logic;
  SIGNAL Logical_Operator_out8261_out1            : std_logic;
  SIGNAL Logical_Operator_out8262_out1            : std_logic;
  SIGNAL Logical_Operator_out8263_out1            : std_logic;
  SIGNAL Logical_Operator_out8264_out1            : std_logic;
  SIGNAL Logical_Operator_out8265_out1            : std_logic;
  SIGNAL Logical_Operator_out8266_out1            : std_logic;
  SIGNAL Logical_Operator_out8267_out1            : std_logic;
  SIGNAL Logical_Operator_out8268_out1            : std_logic;
  SIGNAL Logical_Operator_out8269_out1            : std_logic;
  SIGNAL Logical_Operator_out8270_out1            : std_logic;
  SIGNAL Logical_Operator_out8271_out1            : std_logic;
  SIGNAL Logical_Operator_out8272_out1            : std_logic;
  SIGNAL Logical_Operator_out8273_out1            : std_logic;
  SIGNAL Logical_Operator_out8274_out1            : std_logic;
  SIGNAL Logical_Operator_out8275_out1            : std_logic;
  SIGNAL Logical_Operator_out8276_out1            : std_logic;
  SIGNAL Logical_Operator_out8277_out1            : std_logic;
  SIGNAL Logical_Operator_out8278_out1            : std_logic;
  SIGNAL Logical_Operator_out8279_out1            : std_logic;
  SIGNAL Logical_Operator_out8280_out1            : std_logic;
  SIGNAL Logical_Operator_out8281_out1            : std_logic;
  SIGNAL Logical_Operator_out8282_out1            : std_logic;
  SIGNAL Logical_Operator_out8283_out1            : std_logic;
  SIGNAL Logical_Operator_out8284_out1            : std_logic;
  SIGNAL Logical_Operator_out8285_out1            : std_logic;
  SIGNAL Logical_Operator_out8286_out1            : std_logic;
  SIGNAL Logical_Operator_out8287_out1            : std_logic;
  SIGNAL Logical_Operator_out8288_out1            : std_logic;
  SIGNAL Logical_Operator_out8289_out1            : std_logic;
  SIGNAL Logical_Operator_out8290_out1            : std_logic;
  SIGNAL Logical_Operator_out8291_out1            : std_logic;
  SIGNAL Logical_Operator_out8292_out1            : std_logic;
  SIGNAL Logical_Operator_out8293_out1            : std_logic;
  SIGNAL Logical_Operator_out8294_out1            : std_logic;
  SIGNAL Logical_Operator_out8295_out1            : std_logic;
  SIGNAL Logical_Operator_out8296_out1            : std_logic;
  SIGNAL Logical_Operator_out8297_out1            : std_logic;
  SIGNAL Logical_Operator_out8298_out1            : std_logic;
  SIGNAL Logical_Operator_out8299_out1            : std_logic;
  SIGNAL Logical_Operator_out8300_out1            : std_logic;
  SIGNAL Logical_Operator_out8301_out1            : std_logic;
  SIGNAL Logical_Operator_out8302_out1            : std_logic;
  SIGNAL Logical_Operator_out8303_out1            : std_logic;
  SIGNAL Logical_Operator_out8304_out1            : std_logic;
  SIGNAL Logical_Operator_out8305_out1            : std_logic;
  SIGNAL Logical_Operator_out8306_out1            : std_logic;
  SIGNAL Logical_Operator_out8307_out1            : std_logic;
  SIGNAL Logical_Operator_out8308_out1            : std_logic;
  SIGNAL Logical_Operator_out8309_out1            : std_logic;
  SIGNAL Logical_Operator_out8310_out1            : std_logic;
  SIGNAL Logical_Operator_out8311_out1            : std_logic;
  SIGNAL Logical_Operator_out8312_out1            : std_logic;
  SIGNAL Logical_Operator_out8313_out1            : std_logic;
  SIGNAL Logical_Operator_out8314_out1            : std_logic;
  SIGNAL Logical_Operator_out8315_out1            : std_logic;
  SIGNAL Logical_Operator_out8316_out1            : std_logic;
  SIGNAL Logical_Operator_out8317_out1            : std_logic;
  SIGNAL Logical_Operator_out8318_out1            : std_logic;
  SIGNAL Logical_Operator_out8319_out1            : std_logic;
  SIGNAL Logical_Operator_out8320_out1            : std_logic;
  SIGNAL Logical_Operator_out8321_out1            : std_logic;
  SIGNAL Logical_Operator_out8322_out1            : std_logic;
  SIGNAL Logical_Operator_out8323_out1            : std_logic;
  SIGNAL Logical_Operator_out8324_out1            : std_logic;
  SIGNAL Logical_Operator_out8325_out1            : std_logic;
  SIGNAL Logical_Operator_out8326_out1            : std_logic;
  SIGNAL Logical_Operator_out8327_out1            : std_logic;
  SIGNAL Logical_Operator_out8328_out1            : std_logic;
  SIGNAL Logical_Operator_out8329_out1            : std_logic;
  SIGNAL Logical_Operator_out8330_out1            : std_logic;
  SIGNAL Logical_Operator_out8331_out1            : std_logic;
  SIGNAL Logical_Operator_out8332_out1            : std_logic;
  SIGNAL Logical_Operator_out8333_out1            : std_logic;
  SIGNAL Logical_Operator_out8334_out1            : std_logic;
  SIGNAL Logical_Operator_out8335_out1            : std_logic;
  SIGNAL Logical_Operator_out8336_out1            : std_logic;
  SIGNAL Logical_Operator_out8337_out1            : std_logic;
  SIGNAL Logical_Operator_out8338_out1            : std_logic;
  SIGNAL Logical_Operator_out8339_out1            : std_logic;
  SIGNAL Logical_Operator_out8340_out1            : std_logic;
  SIGNAL Logical_Operator_out8341_out1            : std_logic;
  SIGNAL Logical_Operator_out8342_out1            : std_logic;
  SIGNAL Logical_Operator_out8343_out1            : std_logic;
  SIGNAL Logical_Operator_out8344_out1            : std_logic;
  SIGNAL Logical_Operator_out8345_out1            : std_logic;
  SIGNAL Logical_Operator_out8346_out1            : std_logic;
  SIGNAL Logical_Operator_out8347_out1            : std_logic;
  SIGNAL Logical_Operator_out8348_out1            : std_logic;
  SIGNAL Logical_Operator_out8349_out1            : std_logic;
  SIGNAL Logical_Operator_out8350_out1            : std_logic;
  SIGNAL Logical_Operator_out8351_out1            : std_logic;
  SIGNAL Logical_Operator_out8352_out1            : std_logic;
  SIGNAL Logical_Operator_out8353_out1            : std_logic;
  SIGNAL Logical_Operator_out8354_out1            : std_logic;
  SIGNAL Logical_Operator_out8355_out1            : std_logic;
  SIGNAL Logical_Operator_out8356_out1            : std_logic;
  SIGNAL Logical_Operator_out8357_out1            : std_logic;
  SIGNAL Logical_Operator_out8358_out1            : std_logic;
  SIGNAL Logical_Operator_out8359_out1            : std_logic;
  SIGNAL Logical_Operator_out8360_out1            : std_logic;
  SIGNAL Logical_Operator_out8361_out1            : std_logic;
  SIGNAL Logical_Operator_out8362_out1            : std_logic;
  SIGNAL Logical_Operator_out8363_out1            : std_logic;
  SIGNAL Logical_Operator_out8364_out1            : std_logic;
  SIGNAL Logical_Operator_out8365_out1            : std_logic;
  SIGNAL Logical_Operator_out8366_out1            : std_logic;
  SIGNAL Logical_Operator_out8367_out1            : std_logic;
  SIGNAL Logical_Operator_out8368_out1            : std_logic;
  SIGNAL Logical_Operator_out8369_out1            : std_logic;
  SIGNAL Logical_Operator_out8370_out1            : std_logic;
  SIGNAL Logical_Operator_out8371_out1            : std_logic;
  SIGNAL Logical_Operator_out8372_out1            : std_logic;
  SIGNAL Logical_Operator_out8373_out1            : std_logic;
  SIGNAL Logical_Operator_out8374_out1            : std_logic;
  SIGNAL Logical_Operator_out8375_out1            : std_logic;
  SIGNAL Logical_Operator_out8376_out1            : std_logic;
  SIGNAL Logical_Operator_out8377_out1            : std_logic;
  SIGNAL Logical_Operator_out8378_out1            : std_logic;
  SIGNAL Logical_Operator_out8379_out1            : std_logic;
  SIGNAL Logical_Operator_out8380_out1            : std_logic;
  SIGNAL Logical_Operator_out8381_out1            : std_logic;
  SIGNAL Logical_Operator_out8382_out1            : std_logic;
  SIGNAL Logical_Operator_out8383_out1            : std_logic;
  SIGNAL Logical_Operator_out8384_out1            : std_logic;
  SIGNAL Logical_Operator_out8385_out1            : std_logic;
  SIGNAL Logical_Operator_out8386_out1            : std_logic;
  SIGNAL Logical_Operator_out8387_out1            : std_logic;
  SIGNAL Logical_Operator_out8388_out1            : std_logic;
  SIGNAL Logical_Operator_out8389_out1            : std_logic;
  SIGNAL Logical_Operator_out8390_out1            : std_logic;
  SIGNAL Logical_Operator_out8391_out1            : std_logic;
  SIGNAL Logical_Operator_out8392_out1            : std_logic;
  SIGNAL Logical_Operator_out8393_out1            : std_logic;
  SIGNAL Logical_Operator_out8394_out1            : std_logic;
  SIGNAL Logical_Operator_out8395_out1            : std_logic;
  SIGNAL Logical_Operator_out8396_out1            : std_logic;
  SIGNAL Logical_Operator_out8397_out1            : std_logic;
  SIGNAL Logical_Operator_out8398_out1            : std_logic;
  SIGNAL Logical_Operator_out8399_out1            : std_logic;
  SIGNAL Logical_Operator_out8400_out1            : std_logic;
  SIGNAL Logical_Operator_out8401_out1            : std_logic;
  SIGNAL Logical_Operator_out8402_out1            : std_logic;
  SIGNAL Logical_Operator_out8403_out1            : std_logic;
  SIGNAL Logical_Operator_out8404_out1            : std_logic;
  SIGNAL Logical_Operator_out8405_out1            : std_logic;
  SIGNAL Logical_Operator_out8406_out1            : std_logic;
  SIGNAL Logical_Operator_out8407_out1            : std_logic;
  SIGNAL Logical_Operator_out8408_out1            : std_logic;
  SIGNAL Logical_Operator_out8409_out1            : std_logic;
  SIGNAL Logical_Operator_out8410_out1            : std_logic;
  SIGNAL Logical_Operator_out8411_out1            : std_logic;
  SIGNAL Logical_Operator_out8412_out1            : std_logic;
  SIGNAL Logical_Operator_out8413_out1            : std_logic;
  SIGNAL Logical_Operator_out8414_out1            : std_logic;
  SIGNAL Logical_Operator_out8415_out1            : std_logic;
  SIGNAL Logical_Operator_out8416_out1            : std_logic;
  SIGNAL Logical_Operator_out8417_out1            : std_logic;
  SIGNAL Logical_Operator_out8418_out1            : std_logic;
  SIGNAL Logical_Operator_out8419_out1            : std_logic;
  SIGNAL Logical_Operator_out8420_out1            : std_logic;
  SIGNAL Logical_Operator_out8421_out1            : std_logic;
  SIGNAL Logical_Operator_out8422_out1            : std_logic;
  SIGNAL Logical_Operator_out8423_out1            : std_logic;
  SIGNAL Logical_Operator_out8424_out1            : std_logic;
  SIGNAL Logical_Operator_out8425_out1            : std_logic;
  SIGNAL Logical_Operator_out8426_out1            : std_logic;
  SIGNAL Logical_Operator_out8427_out1            : std_logic;
  SIGNAL Logical_Operator_out8428_out1            : std_logic;
  SIGNAL Logical_Operator_out8429_out1            : std_logic;
  SIGNAL Logical_Operator_out8430_out1            : std_logic;
  SIGNAL Logical_Operator_out8431_out1            : std_logic;
  SIGNAL Logical_Operator_out8432_out1            : std_logic;
  SIGNAL Logical_Operator_out8433_out1            : std_logic;
  SIGNAL Logical_Operator_out8434_out1            : std_logic;
  SIGNAL Logical_Operator_out8435_out1            : std_logic;
  SIGNAL Logical_Operator_out8436_out1            : std_logic;
  SIGNAL Logical_Operator_out8437_out1            : std_logic;
  SIGNAL Logical_Operator_out8438_out1            : std_logic;
  SIGNAL Logical_Operator_out8439_out1            : std_logic;
  SIGNAL Logical_Operator_out8440_out1            : std_logic;
  SIGNAL Logical_Operator_out8441_out1            : std_logic;
  SIGNAL Logical_Operator_out8442_out1            : std_logic;
  SIGNAL Logical_Operator_out8443_out1            : std_logic;
  SIGNAL Logical_Operator_out8444_out1            : std_logic;
  SIGNAL Logical_Operator_out8445_out1            : std_logic;
  SIGNAL Logical_Operator_out8446_out1            : std_logic;
  SIGNAL Logical_Operator_out8447_out1            : std_logic;
  SIGNAL Logical_Operator_out8448_out1            : std_logic;
  SIGNAL Logical_Operator_out8449_out1            : std_logic;
  SIGNAL Logical_Operator_out8450_out1            : std_logic;
  SIGNAL Logical_Operator_out8451_out1            : std_logic;
  SIGNAL Logical_Operator_out8452_out1            : std_logic;
  SIGNAL Logical_Operator_out8453_out1            : std_logic;
  SIGNAL Logical_Operator_out8454_out1            : std_logic;
  SIGNAL Logical_Operator_out8455_out1            : std_logic;
  SIGNAL Logical_Operator_out8456_out1            : std_logic;
  SIGNAL Logical_Operator_out8457_out1            : std_logic;
  SIGNAL Logical_Operator_out8458_out1            : std_logic;
  SIGNAL Logical_Operator_out8459_out1            : std_logic;
  SIGNAL Logical_Operator_out8460_out1            : std_logic;
  SIGNAL Logical_Operator_out8461_out1            : std_logic;
  SIGNAL Logical_Operator_out8462_out1            : std_logic;
  SIGNAL Logical_Operator_out8463_out1            : std_logic;
  SIGNAL Logical_Operator_out8464_out1            : std_logic;
  SIGNAL Logical_Operator_out8465_out1            : std_logic;
  SIGNAL Logical_Operator_out8466_out1            : std_logic;
  SIGNAL Logical_Operator_out8467_out1            : std_logic;
  SIGNAL Logical_Operator_out8468_out1            : std_logic;
  SIGNAL Logical_Operator_out8469_out1            : std_logic;
  SIGNAL Logical_Operator_out8470_out1            : std_logic;
  SIGNAL Logical_Operator_out8471_out1            : std_logic;
  SIGNAL Logical_Operator_out8472_out1            : std_logic;
  SIGNAL Logical_Operator_out8473_out1            : std_logic;
  SIGNAL Logical_Operator_out8474_out1            : std_logic;
  SIGNAL Logical_Operator_out8475_out1            : std_logic;
  SIGNAL Logical_Operator_out8476_out1            : std_logic;
  SIGNAL Logical_Operator_out8477_out1            : std_logic;
  SIGNAL Logical_Operator_out8478_out1            : std_logic;
  SIGNAL Logical_Operator_out8479_out1            : std_logic;
  SIGNAL Logical_Operator_out8480_out1            : std_logic;
  SIGNAL Logical_Operator_out8481_out1            : std_logic;
  SIGNAL Logical_Operator_out8482_out1            : std_logic;
  SIGNAL Logical_Operator_out8483_out1            : std_logic;
  SIGNAL Logical_Operator_out8484_out1            : std_logic;
  SIGNAL Logical_Operator_out8485_out1            : std_logic;
  SIGNAL Logical_Operator_out8486_out1            : std_logic;
  SIGNAL Logical_Operator_out8487_out1            : std_logic;
  SIGNAL Logical_Operator_out8488_out1            : std_logic;
  SIGNAL Logical_Operator_out8489_out1            : std_logic;
  SIGNAL Logical_Operator_out8490_out1            : std_logic;
  SIGNAL Logical_Operator_out8491_out1            : std_logic;
  SIGNAL Logical_Operator_out8492_out1            : std_logic;
  SIGNAL Logical_Operator_out8493_out1            : std_logic;
  SIGNAL Logical_Operator_out8494_out1            : std_logic;
  SIGNAL Logical_Operator_out8495_out1            : std_logic;
  SIGNAL Logical_Operator_out8496_out1            : std_logic;
  SIGNAL Logical_Operator_out8497_out1            : std_logic;
  SIGNAL Logical_Operator_out8498_out1            : std_logic;
  SIGNAL Logical_Operator_out8499_out1            : std_logic;
  SIGNAL Logical_Operator_out8500_out1            : std_logic;
  SIGNAL Logical_Operator_out8501_out1            : std_logic;
  SIGNAL Logical_Operator_out8502_out1            : std_logic;
  SIGNAL Logical_Operator_out8503_out1            : std_logic;
  SIGNAL Logical_Operator_out8504_out1            : std_logic;
  SIGNAL Logical_Operator_out8505_out1            : std_logic;
  SIGNAL Logical_Operator_out8506_out1            : std_logic;
  SIGNAL Logical_Operator_out8507_out1            : std_logic;
  SIGNAL Logical_Operator_out8508_out1            : std_logic;
  SIGNAL Logical_Operator_out8509_out1            : std_logic;
  SIGNAL Logical_Operator_out8510_out1            : std_logic;
  SIGNAL Logical_Operator_out8511_out1            : std_logic;
  SIGNAL Logical_Operator_out8512_out1            : std_logic;
  SIGNAL Logical_Operator_out8513_out1            : std_logic;
  SIGNAL Logical_Operator_out8514_out1            : std_logic;
  SIGNAL Logical_Operator_out8515_out1            : std_logic;
  SIGNAL Logical_Operator_out8516_out1            : std_logic;
  SIGNAL Logical_Operator_out8517_out1            : std_logic;
  SIGNAL Logical_Operator_out8518_out1            : std_logic;
  SIGNAL Logical_Operator_out8519_out1            : std_logic;
  SIGNAL Logical_Operator_out8520_out1            : std_logic;
  SIGNAL Logical_Operator_out8521_out1            : std_logic;
  SIGNAL Logical_Operator_out8522_out1            : std_logic;
  SIGNAL Logical_Operator_out8523_out1            : std_logic;
  SIGNAL Logical_Operator_out8524_out1            : std_logic;
  SIGNAL Logical_Operator_out8525_out1            : std_logic;
  SIGNAL Logical_Operator_out8526_out1            : std_logic;
  SIGNAL Logical_Operator_out8527_out1            : std_logic;
  SIGNAL Logical_Operator_out8528_out1            : std_logic;
  SIGNAL Logical_Operator_out8529_out1            : std_logic;
  SIGNAL Logical_Operator_out8530_out1            : std_logic;
  SIGNAL Logical_Operator_out8531_out1            : std_logic;
  SIGNAL Logical_Operator_out8532_out1            : std_logic;
  SIGNAL Logical_Operator_out8533_out1            : std_logic;
  SIGNAL Logical_Operator_out8534_out1            : std_logic;
  SIGNAL Logical_Operator_out8535_out1            : std_logic;
  SIGNAL Logical_Operator_out8536_out1            : std_logic;
  SIGNAL Logical_Operator_out8537_out1            : std_logic;
  SIGNAL Logical_Operator_out8538_out1            : std_logic;
  SIGNAL Logical_Operator_out8539_out1            : std_logic;
  SIGNAL Logical_Operator_out8540_out1            : std_logic;
  SIGNAL Logical_Operator_out8541_out1            : std_logic;
  SIGNAL Logical_Operator_out8542_out1            : std_logic;
  SIGNAL Logical_Operator_out8543_out1            : std_logic;
  SIGNAL Logical_Operator_out8544_out1            : std_logic;
  SIGNAL Logical_Operator_out8545_out1            : std_logic;
  SIGNAL Logical_Operator_out8546_out1            : std_logic;
  SIGNAL Logical_Operator_out8547_out1            : std_logic;
  SIGNAL Logical_Operator_out8548_out1            : std_logic;
  SIGNAL Logical_Operator_out8549_out1            : std_logic;
  SIGNAL Logical_Operator_out8550_out1            : std_logic;
  SIGNAL Logical_Operator_out8551_out1            : std_logic;
  SIGNAL Logical_Operator_out8552_out1            : std_logic;
  SIGNAL Logical_Operator_out8553_out1            : std_logic;
  SIGNAL Logical_Operator_out8554_out1            : std_logic;
  SIGNAL Logical_Operator_out8555_out1            : std_logic;
  SIGNAL Logical_Operator_out8556_out1            : std_logic;
  SIGNAL Logical_Operator_out8557_out1            : std_logic;
  SIGNAL Logical_Operator_out8558_out1            : std_logic;
  SIGNAL Logical_Operator_out8559_out1            : std_logic;
  SIGNAL Logical_Operator_out8560_out1            : std_logic;
  SIGNAL Logical_Operator_out8561_out1            : std_logic;
  SIGNAL Logical_Operator_out8562_out1            : std_logic;
  SIGNAL Logical_Operator_out8563_out1            : std_logic;
  SIGNAL Logical_Operator_out8564_out1            : std_logic;
  SIGNAL Logical_Operator_out8565_out1            : std_logic;
  SIGNAL Logical_Operator_out8566_out1            : std_logic;
  SIGNAL Logical_Operator_out8567_out1            : std_logic;
  SIGNAL Logical_Operator_out8568_out1            : std_logic;
  SIGNAL Logical_Operator_out8569_out1            : std_logic;
  SIGNAL Logical_Operator_out8570_out1            : std_logic;
  SIGNAL Logical_Operator_out8571_out1            : std_logic;
  SIGNAL Logical_Operator_out8572_out1            : std_logic;
  SIGNAL Logical_Operator_out8573_out1            : std_logic;
  SIGNAL Logical_Operator_out8574_out1            : std_logic;
  SIGNAL Logical_Operator_out8575_out1            : std_logic;
  SIGNAL Logical_Operator_out8576_out1            : std_logic;
  SIGNAL Logical_Operator_out8577_out1            : std_logic;
  SIGNAL Logical_Operator_out8578_out1            : std_logic;
  SIGNAL Logical_Operator_out8579_out1            : std_logic;
  SIGNAL Logical_Operator_out8580_out1            : std_logic;
  SIGNAL Logical_Operator_out8581_out1            : std_logic;
  SIGNAL Logical_Operator_out8582_out1            : std_logic;
  SIGNAL Logical_Operator_out8583_out1            : std_logic;
  SIGNAL Logical_Operator_out8584_out1            : std_logic;
  SIGNAL Logical_Operator_out8585_out1            : std_logic;
  SIGNAL Logical_Operator_out8586_out1            : std_logic;
  SIGNAL Logical_Operator_out8587_out1            : std_logic;
  SIGNAL Logical_Operator_out8588_out1            : std_logic;
  SIGNAL Logical_Operator_out8589_out1            : std_logic;
  SIGNAL Logical_Operator_out8590_out1            : std_logic;
  SIGNAL Logical_Operator_out8591_out1            : std_logic;
  SIGNAL Logical_Operator_out8592_out1            : std_logic;
  SIGNAL Logical_Operator_out8593_out1            : std_logic;
  SIGNAL Logical_Operator_out8594_out1            : std_logic;
  SIGNAL Logical_Operator_out8595_out1            : std_logic;
  SIGNAL Logical_Operator_out8596_out1            : std_logic;
  SIGNAL Logical_Operator_out8597_out1            : std_logic;
  SIGNAL Logical_Operator_out8598_out1            : std_logic;
  SIGNAL Logical_Operator_out8599_out1            : std_logic;
  SIGNAL Logical_Operator_out8600_out1            : std_logic;
  SIGNAL Logical_Operator_out8601_out1            : std_logic;
  SIGNAL Logical_Operator_out8602_out1            : std_logic;
  SIGNAL Logical_Operator_out8603_out1            : std_logic;
  SIGNAL Logical_Operator_out8604_out1            : std_logic;
  SIGNAL Logical_Operator_out8605_out1            : std_logic;
  SIGNAL Logical_Operator_out8606_out1            : std_logic;
  SIGNAL Logical_Operator_out8607_out1            : std_logic;
  SIGNAL Logical_Operator_out8608_out1            : std_logic;
  SIGNAL Logical_Operator_out8609_out1            : std_logic;
  SIGNAL Logical_Operator_out8610_out1            : std_logic;
  SIGNAL Logical_Operator_out8611_out1            : std_logic;
  SIGNAL Logical_Operator_out8612_out1            : std_logic;
  SIGNAL Logical_Operator_out8613_out1            : std_logic;
  SIGNAL Logical_Operator_out8614_out1            : std_logic;
  SIGNAL Logical_Operator_out8615_out1            : std_logic;
  SIGNAL Logical_Operator_out8616_out1            : std_logic;
  SIGNAL Logical_Operator_out8617_out1            : std_logic;
  SIGNAL Logical_Operator_out8618_out1            : std_logic;
  SIGNAL Logical_Operator_out8619_out1            : std_logic;
  SIGNAL Logical_Operator_out8620_out1            : std_logic;
  SIGNAL Logical_Operator_out8621_out1            : std_logic;
  SIGNAL Logical_Operator_out8622_out1            : std_logic;
  SIGNAL Logical_Operator_out8623_out1            : std_logic;
  SIGNAL Logical_Operator_out8624_out1            : std_logic;
  SIGNAL Logical_Operator_out8625_out1            : std_logic;
  SIGNAL Logical_Operator_out8626_out1            : std_logic;
  SIGNAL Logical_Operator_out8627_out1            : std_logic;
  SIGNAL Logical_Operator_out8628_out1            : std_logic;
  SIGNAL Logical_Operator_out8629_out1            : std_logic;
  SIGNAL Logical_Operator_out8630_out1            : std_logic;
  SIGNAL Logical_Operator_out8631_out1            : std_logic;
  SIGNAL Logical_Operator_out8632_out1            : std_logic;
  SIGNAL Logical_Operator_out8633_out1            : std_logic;
  SIGNAL Logical_Operator_out8634_out1            : std_logic;
  SIGNAL Logical_Operator_out8635_out1            : std_logic;
  SIGNAL Logical_Operator_out8636_out1            : std_logic;
  SIGNAL Logical_Operator_out8637_out1            : std_logic;
  SIGNAL Logical_Operator_out8638_out1            : std_logic;
  SIGNAL Logical_Operator_out8639_out1            : std_logic;
  SIGNAL Logical_Operator_out8640_out1            : std_logic;
  SIGNAL Logical_Operator_out8641_out1            : std_logic;
  SIGNAL Logical_Operator_out8642_out1            : std_logic;
  SIGNAL Logical_Operator_out8643_out1            : std_logic;
  SIGNAL Logical_Operator_out8644_out1            : std_logic;
  SIGNAL Logical_Operator_out8645_out1            : std_logic;
  SIGNAL Logical_Operator_out8646_out1            : std_logic;
  SIGNAL Logical_Operator_out8647_out1            : std_logic;
  SIGNAL Logical_Operator_out8648_out1            : std_logic;
  SIGNAL Logical_Operator_out8649_out1            : std_logic;
  SIGNAL Logical_Operator_out8650_out1            : std_logic;
  SIGNAL Logical_Operator_out8651_out1            : std_logic;
  SIGNAL Logical_Operator_out8652_out1            : std_logic;
  SIGNAL Logical_Operator_out8653_out1            : std_logic;
  SIGNAL Logical_Operator_out8654_out1            : std_logic;
  SIGNAL Logical_Operator_out8655_out1            : std_logic;
  SIGNAL Logical_Operator_out8656_out1            : std_logic;
  SIGNAL Logical_Operator_out8657_out1            : std_logic;
  SIGNAL Logical_Operator_out8658_out1            : std_logic;
  SIGNAL Logical_Operator_out8659_out1            : std_logic;
  SIGNAL Logical_Operator_out8660_out1            : std_logic;
  SIGNAL Logical_Operator_out8661_out1            : std_logic;
  SIGNAL Logical_Operator_out8662_out1            : std_logic;
  SIGNAL Logical_Operator_out8663_out1            : std_logic;
  SIGNAL Logical_Operator_out8664_out1            : std_logic;
  SIGNAL Logical_Operator_out8665_out1            : std_logic;
  SIGNAL Logical_Operator_out8666_out1            : std_logic;
  SIGNAL Logical_Operator_out8667_out1            : std_logic;
  SIGNAL Logical_Operator_out8668_out1            : std_logic;
  SIGNAL Logical_Operator_out8669_out1            : std_logic;
  SIGNAL Logical_Operator_out8670_out1            : std_logic;
  SIGNAL Logical_Operator_out8671_out1            : std_logic;
  SIGNAL Logical_Operator_out8672_out1            : std_logic;
  SIGNAL Logical_Operator_out8673_out1            : std_logic;
  SIGNAL Logical_Operator_out8674_out1            : std_logic;
  SIGNAL Logical_Operator_out8675_out1            : std_logic;
  SIGNAL Logical_Operator_out8676_out1            : std_logic;
  SIGNAL Logical_Operator_out8677_out1            : std_logic;
  SIGNAL Logical_Operator_out8678_out1            : std_logic;
  SIGNAL Logical_Operator_out8679_out1            : std_logic;
  SIGNAL Logical_Operator_out8680_out1            : std_logic;
  SIGNAL Logical_Operator_out8681_out1            : std_logic;
  SIGNAL Logical_Operator_out8682_out1            : std_logic;
  SIGNAL Logical_Operator_out8683_out1            : std_logic;
  SIGNAL Logical_Operator_out8684_out1            : std_logic;
  SIGNAL Logical_Operator_out8685_out1            : std_logic;
  SIGNAL Logical_Operator_out8686_out1            : std_logic;
  SIGNAL Logical_Operator_out8687_out1            : std_logic;
  SIGNAL Logical_Operator_out8688_out1            : std_logic;
  SIGNAL Logical_Operator_out8689_out1            : std_logic;
  SIGNAL Logical_Operator_out8690_out1            : std_logic;
  SIGNAL Logical_Operator_out8691_out1            : std_logic;
  SIGNAL Logical_Operator_out8692_out1            : std_logic;
  SIGNAL Logical_Operator_out8693_out1            : std_logic;
  SIGNAL Logical_Operator_out8694_out1            : std_logic;
  SIGNAL Logical_Operator_out8695_out1            : std_logic;
  SIGNAL Logical_Operator_out8696_out1            : std_logic;
  SIGNAL Logical_Operator_out8697_out1            : std_logic;
  SIGNAL Logical_Operator_out8698_out1            : std_logic;
  SIGNAL Logical_Operator_out8699_out1            : std_logic;
  SIGNAL Logical_Operator_out8700_out1            : std_logic;
  SIGNAL Logical_Operator_out8701_out1            : std_logic;
  SIGNAL Logical_Operator_out8702_out1            : std_logic;
  SIGNAL Logical_Operator_out8703_out1            : std_logic;
  SIGNAL Logical_Operator_out8704_out1            : std_logic;
  SIGNAL Logical_Operator_out8705_out1            : std_logic;
  SIGNAL Logical_Operator_out8706_out1            : std_logic;
  SIGNAL Logical_Operator_out8707_out1            : std_logic;
  SIGNAL Logical_Operator_out8708_out1            : std_logic;
  SIGNAL Logical_Operator_out8709_out1            : std_logic;
  SIGNAL Logical_Operator_out8710_out1            : std_logic;
  SIGNAL Logical_Operator_out8711_out1            : std_logic;
  SIGNAL Logical_Operator_out8712_out1            : std_logic;
  SIGNAL Logical_Operator_out8713_out1            : std_logic;
  SIGNAL Logical_Operator_out8714_out1            : std_logic;
  SIGNAL Logical_Operator_out8715_out1            : std_logic;
  SIGNAL Logical_Operator_out8716_out1            : std_logic;
  SIGNAL Logical_Operator_out8717_out1            : std_logic;
  SIGNAL Logical_Operator_out8718_out1            : std_logic;
  SIGNAL Logical_Operator_out8719_out1            : std_logic;
  SIGNAL Logical_Operator_out8720_out1            : std_logic;
  SIGNAL Logical_Operator_out8721_out1            : std_logic;
  SIGNAL Logical_Operator_out8722_out1            : std_logic;
  SIGNAL Logical_Operator_out8723_out1            : std_logic;
  SIGNAL Logical_Operator_out8724_out1            : std_logic;
  SIGNAL Logical_Operator_out8725_out1            : std_logic;
  SIGNAL Logical_Operator_out8726_out1            : std_logic;
  SIGNAL Logical_Operator_out8727_out1            : std_logic;
  SIGNAL Logical_Operator_out8728_out1            : std_logic;
  SIGNAL Logical_Operator_out8729_out1            : std_logic;
  SIGNAL Logical_Operator_out8730_out1            : std_logic;
  SIGNAL Logical_Operator_out8731_out1            : std_logic;
  SIGNAL Logical_Operator_out8732_out1            : std_logic;
  SIGNAL Logical_Operator_out8733_out1            : std_logic;
  SIGNAL Logical_Operator_out8734_out1            : std_logic;
  SIGNAL Logical_Operator_out8735_out1            : std_logic;
  SIGNAL Logical_Operator_out8736_out1            : std_logic;
  SIGNAL Logical_Operator_out8737_out1            : std_logic;
  SIGNAL Logical_Operator_out8738_out1            : std_logic;
  SIGNAL Logical_Operator_out8739_out1            : std_logic;
  SIGNAL Logical_Operator_out8740_out1            : std_logic;
  SIGNAL Logical_Operator_out8741_out1            : std_logic;
  SIGNAL Logical_Operator_out8742_out1            : std_logic;
  SIGNAL Logical_Operator_out8743_out1            : std_logic;
  SIGNAL Logical_Operator_out8744_out1            : std_logic;
  SIGNAL Logical_Operator_out8745_out1            : std_logic;
  SIGNAL Logical_Operator_out8746_out1            : std_logic;
  SIGNAL Logical_Operator_out8747_out1            : std_logic;
  SIGNAL Logical_Operator_out8748_out1            : std_logic;
  SIGNAL Logical_Operator_out8749_out1            : std_logic;
  SIGNAL Logical_Operator_out8750_out1            : std_logic;
  SIGNAL Logical_Operator_out8751_out1            : std_logic;
  SIGNAL Logical_Operator_out8752_out1            : std_logic;
  SIGNAL Logical_Operator_out8753_out1            : std_logic;
  SIGNAL Logical_Operator_out8754_out1            : std_logic;
  SIGNAL Logical_Operator_out8755_out1            : std_logic;
  SIGNAL Logical_Operator_out8756_out1            : std_logic;
  SIGNAL Logical_Operator_out8757_out1            : std_logic;
  SIGNAL Logical_Operator_out8758_out1            : std_logic;
  SIGNAL Logical_Operator_out8759_out1            : std_logic;
  SIGNAL Logical_Operator_out8760_out1            : std_logic;
  SIGNAL Logical_Operator_out8761_out1            : std_logic;
  SIGNAL Logical_Operator_out8762_out1            : std_logic;
  SIGNAL Logical_Operator_out8763_out1            : std_logic;
  SIGNAL Logical_Operator_out8764_out1            : std_logic;
  SIGNAL Logical_Operator_out8765_out1            : std_logic;
  SIGNAL Logical_Operator_out8766_out1            : std_logic;
  SIGNAL Logical_Operator_out8767_out1            : std_logic;
  SIGNAL Logical_Operator_out8768_out1            : std_logic;
  SIGNAL Logical_Operator_out8769_out1            : std_logic;
  SIGNAL Logical_Operator_out8770_out1            : std_logic;
  SIGNAL Logical_Operator_out8771_out1            : std_logic;
  SIGNAL Logical_Operator_out8772_out1            : std_logic;
  SIGNAL Logical_Operator_out8773_out1            : std_logic;
  SIGNAL Logical_Operator_out8774_out1            : std_logic;
  SIGNAL Logical_Operator_out8775_out1            : std_logic;
  SIGNAL Logical_Operator_out8776_out1            : std_logic;
  SIGNAL Logical_Operator_out8777_out1            : std_logic;
  SIGNAL Logical_Operator_out8778_out1            : std_logic;
  SIGNAL Logical_Operator_out8779_out1            : std_logic;
  SIGNAL Logical_Operator_out8780_out1            : std_logic;
  SIGNAL Logical_Operator_out8781_out1            : std_logic;
  SIGNAL Logical_Operator_out8782_out1            : std_logic;
  SIGNAL Logical_Operator_out8783_out1            : std_logic;
  SIGNAL Logical_Operator_out8784_out1            : std_logic;
  SIGNAL Logical_Operator_out8785_out1            : std_logic;
  SIGNAL Logical_Operator_out8786_out1            : std_logic;
  SIGNAL Logical_Operator_out8787_out1            : std_logic;
  SIGNAL Logical_Operator_out8788_out1            : std_logic;
  SIGNAL Logical_Operator_out8789_out1            : std_logic;
  SIGNAL Logical_Operator_out8790_out1            : std_logic;
  SIGNAL Logical_Operator_out8791_out1            : std_logic;
  SIGNAL Logical_Operator_out8792_out1            : std_logic;
  SIGNAL Logical_Operator_out8793_out1            : std_logic;
  SIGNAL Logical_Operator_out8794_out1            : std_logic;
  SIGNAL Logical_Operator_out8795_out1            : std_logic;
  SIGNAL Logical_Operator_out8796_out1            : std_logic;
  SIGNAL Logical_Operator_out8797_out1            : std_logic;
  SIGNAL Logical_Operator_out8798_out1            : std_logic;
  SIGNAL Logical_Operator_out8799_out1            : std_logic;
  SIGNAL Logical_Operator_out8800_out1            : std_logic;
  SIGNAL Logical_Operator_out8801_out1            : std_logic;
  SIGNAL Logical_Operator_out8802_out1            : std_logic;
  SIGNAL Logical_Operator_out8803_out1            : std_logic;
  SIGNAL Logical_Operator_out8804_out1            : std_logic;
  SIGNAL Logical_Operator_out8805_out1            : std_logic;
  SIGNAL Logical_Operator_out8806_out1            : std_logic;
  SIGNAL Logical_Operator_out8807_out1            : std_logic;
  SIGNAL Logical_Operator_out8808_out1            : std_logic;
  SIGNAL Logical_Operator_out8809_out1            : std_logic;
  SIGNAL Logical_Operator_out8810_out1            : std_logic;
  SIGNAL Logical_Operator_out8811_out1            : std_logic;
  SIGNAL Logical_Operator_out8812_out1            : std_logic;
  SIGNAL Logical_Operator_out8813_out1            : std_logic;
  SIGNAL Logical_Operator_out8814_out1            : std_logic;
  SIGNAL Logical_Operator_out8815_out1            : std_logic;
  SIGNAL Logical_Operator_out8816_out1            : std_logic;
  SIGNAL Logical_Operator_out8817_out1            : std_logic;
  SIGNAL Logical_Operator_out8818_out1            : std_logic;
  SIGNAL Logical_Operator_out8819_out1            : std_logic;
  SIGNAL Logical_Operator_out8820_out1            : std_logic;
  SIGNAL Logical_Operator_out8821_out1            : std_logic;
  SIGNAL Logical_Operator_out8822_out1            : std_logic;
  SIGNAL Logical_Operator_out8823_out1            : std_logic;
  SIGNAL Logical_Operator_out8824_out1            : std_logic;
  SIGNAL Logical_Operator_out8825_out1            : std_logic;
  SIGNAL Logical_Operator_out8826_out1            : std_logic;
  SIGNAL Logical_Operator_out8827_out1            : std_logic;
  SIGNAL Logical_Operator_out8828_out1            : std_logic;
  SIGNAL Logical_Operator_out8829_out1            : std_logic;
  SIGNAL Logical_Operator_out8830_out1            : std_logic;
  SIGNAL Logical_Operator_out8831_out1            : std_logic;
  SIGNAL Logical_Operator_out8832_out1            : std_logic;
  SIGNAL Logical_Operator_out8833_out1            : std_logic;
  SIGNAL Logical_Operator_out8834_out1            : std_logic;
  SIGNAL Logical_Operator_out8835_out1            : std_logic;
  SIGNAL Logical_Operator_out8836_out1            : std_logic;
  SIGNAL Logical_Operator_out8837_out1            : std_logic;
  SIGNAL Logical_Operator_out8838_out1            : std_logic;
  SIGNAL Logical_Operator_out8839_out1            : std_logic;
  SIGNAL Logical_Operator_out8840_out1            : std_logic;
  SIGNAL Logical_Operator_out8841_out1            : std_logic;
  SIGNAL Logical_Operator_out8842_out1            : std_logic;
  SIGNAL Logical_Operator_out8843_out1            : std_logic;
  SIGNAL Logical_Operator_out8844_out1            : std_logic;
  SIGNAL Logical_Operator_out8845_out1            : std_logic;
  SIGNAL Logical_Operator_out8846_out1            : std_logic;
  SIGNAL Logical_Operator_out8847_out1            : std_logic;
  SIGNAL Logical_Operator_out8848_out1            : std_logic;
  SIGNAL Logical_Operator_out8849_out1            : std_logic;
  SIGNAL Logical_Operator_out8850_out1            : std_logic;
  SIGNAL Logical_Operator_out8851_out1            : std_logic;
  SIGNAL Logical_Operator_out8852_out1            : std_logic;
  SIGNAL Logical_Operator_out8853_out1            : std_logic;
  SIGNAL Logical_Operator_out8854_out1            : std_logic;
  SIGNAL Logical_Operator_out8855_out1            : std_logic;
  SIGNAL Logical_Operator_out8856_out1            : std_logic;
  SIGNAL Logical_Operator_out8857_out1            : std_logic;
  SIGNAL Logical_Operator_out8858_out1            : std_logic;
  SIGNAL Logical_Operator_out8859_out1            : std_logic;
  SIGNAL Logical_Operator_out8860_out1            : std_logic;
  SIGNAL Logical_Operator_out8861_out1            : std_logic;
  SIGNAL Logical_Operator_out8862_out1            : std_logic;
  SIGNAL Logical_Operator_out8863_out1            : std_logic;
  SIGNAL Logical_Operator_out8864_out1            : std_logic;
  SIGNAL Logical_Operator_out8865_out1            : std_logic;
  SIGNAL Logical_Operator_out8866_out1            : std_logic;
  SIGNAL Logical_Operator_out8867_out1            : std_logic;
  SIGNAL Logical_Operator_out8868_out1            : std_logic;
  SIGNAL Logical_Operator_out8869_out1            : std_logic;
  SIGNAL Logical_Operator_out8870_out1            : std_logic;
  SIGNAL Logical_Operator_out8871_out1            : std_logic;
  SIGNAL Logical_Operator_out8872_out1            : std_logic;
  SIGNAL Logical_Operator_out8873_out1            : std_logic;
  SIGNAL Logical_Operator_out8874_out1            : std_logic;
  SIGNAL Logical_Operator_out8875_out1            : std_logic;
  SIGNAL Logical_Operator_out8876_out1            : std_logic;
  SIGNAL Logical_Operator_out8877_out1            : std_logic;
  SIGNAL Logical_Operator_out8878_out1            : std_logic;
  SIGNAL Logical_Operator_out8879_out1            : std_logic;
  SIGNAL Logical_Operator_out8880_out1            : std_logic;
  SIGNAL Logical_Operator_out8881_out1            : std_logic;
  SIGNAL Logical_Operator_out8882_out1            : std_logic;
  SIGNAL Logical_Operator_out8883_out1            : std_logic;
  SIGNAL Logical_Operator_out8884_out1            : std_logic;
  SIGNAL Logical_Operator_out8885_out1            : std_logic;
  SIGNAL Logical_Operator_out8886_out1            : std_logic;
  SIGNAL Logical_Operator_out8887_out1            : std_logic;
  SIGNAL Logical_Operator_out8888_out1            : std_logic;
  SIGNAL Logical_Operator_out8889_out1            : std_logic;
  SIGNAL Logical_Operator_out8890_out1            : std_logic;
  SIGNAL Logical_Operator_out8891_out1            : std_logic;
  SIGNAL Logical_Operator_out8892_out1            : std_logic;
  SIGNAL Logical_Operator_out8893_out1            : std_logic;
  SIGNAL Logical_Operator_out8894_out1            : std_logic;
  SIGNAL Logical_Operator_out8895_out1            : std_logic;
  SIGNAL Logical_Operator_out8896_out1            : std_logic;
  SIGNAL Logical_Operator_out8897_out1            : std_logic;
  SIGNAL Logical_Operator_out8898_out1            : std_logic;
  SIGNAL Logical_Operator_out8899_out1            : std_logic;
  SIGNAL Logical_Operator_out8900_out1            : std_logic;
  SIGNAL Logical_Operator_out8901_out1            : std_logic;
  SIGNAL Logical_Operator_out8902_out1            : std_logic;
  SIGNAL Logical_Operator_out8903_out1            : std_logic;
  SIGNAL Logical_Operator_out8904_out1            : std_logic;
  SIGNAL Logical_Operator_out8905_out1            : std_logic;
  SIGNAL Logical_Operator_out8906_out1            : std_logic;
  SIGNAL Logical_Operator_out8907_out1            : std_logic;
  SIGNAL Logical_Operator_out8908_out1            : std_logic;
  SIGNAL Logical_Operator_out8909_out1            : std_logic;
  SIGNAL Logical_Operator_out8910_out1            : std_logic;
  SIGNAL Logical_Operator_out8911_out1            : std_logic;
  SIGNAL Logical_Operator_out8912_out1            : std_logic;
  SIGNAL Logical_Operator_out8913_out1            : std_logic;
  SIGNAL Logical_Operator_out8914_out1            : std_logic;
  SIGNAL Logical_Operator_out8915_out1            : std_logic;
  SIGNAL Logical_Operator_out8916_out1            : std_logic;
  SIGNAL Logical_Operator_out8917_out1            : std_logic;
  SIGNAL Logical_Operator_out8918_out1            : std_logic;
  SIGNAL Logical_Operator_out8919_out1            : std_logic;
  SIGNAL Logical_Operator_out8920_out1            : std_logic;
  SIGNAL Logical_Operator_out8921_out1            : std_logic;
  SIGNAL Logical_Operator_out8922_out1            : std_logic;
  SIGNAL Logical_Operator_out8923_out1            : std_logic;
  SIGNAL Logical_Operator_out8924_out1            : std_logic;
  SIGNAL Logical_Operator_out8925_out1            : std_logic;
  SIGNAL Logical_Operator_out8926_out1            : std_logic;
  SIGNAL Logical_Operator_out8927_out1            : std_logic;
  SIGNAL Logical_Operator_out8928_out1            : std_logic;
  SIGNAL Logical_Operator_out8929_out1            : std_logic;
  SIGNAL Logical_Operator_out8930_out1            : std_logic;
  SIGNAL Logical_Operator_out8931_out1            : std_logic;
  SIGNAL Logical_Operator_out8932_out1            : std_logic;
  SIGNAL Logical_Operator_out8933_out1            : std_logic;
  SIGNAL Logical_Operator_out8934_out1            : std_logic;
  SIGNAL Logical_Operator_out8935_out1            : std_logic;
  SIGNAL Logical_Operator_out8936_out1            : std_logic;
  SIGNAL Logical_Operator_out8937_out1            : std_logic;
  SIGNAL Logical_Operator_out8938_out1            : std_logic;
  SIGNAL Logical_Operator_out8939_out1            : std_logic;
  SIGNAL Logical_Operator_out8940_out1            : std_logic;
  SIGNAL Logical_Operator_out8941_out1            : std_logic;
  SIGNAL Logical_Operator_out8942_out1            : std_logic;
  SIGNAL Logical_Operator_out8943_out1            : std_logic;
  SIGNAL Logical_Operator_out8944_out1            : std_logic;
  SIGNAL Logical_Operator_out8945_out1            : std_logic;
  SIGNAL Logical_Operator_out8946_out1            : std_logic;
  SIGNAL Logical_Operator_out8947_out1            : std_logic;
  SIGNAL Logical_Operator_out8948_out1            : std_logic;
  SIGNAL Logical_Operator_out8949_out1            : std_logic;
  SIGNAL Logical_Operator_out8950_out1            : std_logic;
  SIGNAL Logical_Operator_out8951_out1            : std_logic;
  SIGNAL Logical_Operator_out8952_out1            : std_logic;
  SIGNAL Logical_Operator_out8953_out1            : std_logic;
  SIGNAL Logical_Operator_out8954_out1            : std_logic;
  SIGNAL Logical_Operator_out8955_out1            : std_logic;
  SIGNAL Logical_Operator_out8956_out1            : std_logic;
  SIGNAL Logical_Operator_out8957_out1            : std_logic;
  SIGNAL Logical_Operator_out8958_out1            : std_logic;
  SIGNAL Logical_Operator_out8959_out1            : std_logic;
  SIGNAL Logical_Operator_out8960_out1            : std_logic;
  SIGNAL Logical_Operator_out8961_out1            : std_logic;
  SIGNAL Logical_Operator_out8962_out1            : std_logic;
  SIGNAL Logical_Operator_out8963_out1            : std_logic;
  SIGNAL Logical_Operator_out8964_out1            : std_logic;
  SIGNAL Logical_Operator_out8965_out1            : std_logic;
  SIGNAL Logical_Operator_out8966_out1            : std_logic;
  SIGNAL Logical_Operator_out8967_out1            : std_logic;
  SIGNAL Logical_Operator_out8968_out1            : std_logic;
  SIGNAL Logical_Operator_out8969_out1            : std_logic;
  SIGNAL Logical_Operator_out8970_out1            : std_logic;
  SIGNAL Logical_Operator_out8971_out1            : std_logic;
  SIGNAL Logical_Operator_out8972_out1            : std_logic;
  SIGNAL Logical_Operator_out8973_out1            : std_logic;
  SIGNAL Logical_Operator_out8974_out1            : std_logic;
  SIGNAL Logical_Operator_out8975_out1            : std_logic;
  SIGNAL Logical_Operator_out8976_out1            : std_logic;
  SIGNAL Logical_Operator_out8977_out1            : std_logic;
  SIGNAL Logical_Operator_out8978_out1            : std_logic;
  SIGNAL Logical_Operator_out8979_out1            : std_logic;
  SIGNAL Logical_Operator_out8980_out1            : std_logic;
  SIGNAL Logical_Operator_out8981_out1            : std_logic;
  SIGNAL Logical_Operator_out8982_out1            : std_logic;
  SIGNAL Logical_Operator_out8983_out1            : std_logic;
  SIGNAL Logical_Operator_out8984_out1            : std_logic;
  SIGNAL Logical_Operator_out8985_out1            : std_logic;
  SIGNAL Logical_Operator_out8986_out1            : std_logic;
  SIGNAL Logical_Operator_out8987_out1            : std_logic;
  SIGNAL Logical_Operator_out8988_out1            : std_logic;
  SIGNAL Logical_Operator_out8989_out1            : std_logic;
  SIGNAL Logical_Operator_out8990_out1            : std_logic;
  SIGNAL Logical_Operator_out8991_out1            : std_logic;
  SIGNAL Logical_Operator_out8992_out1            : std_logic;
  SIGNAL Logical_Operator_out8993_out1            : std_logic;
  SIGNAL Logical_Operator_out8994_out1            : std_logic;
  SIGNAL Logical_Operator_out8995_out1            : std_logic;
  SIGNAL Logical_Operator_out8996_out1            : std_logic;
  SIGNAL Logical_Operator_out8997_out1            : std_logic;
  SIGNAL Logical_Operator_out8998_out1            : std_logic;
  SIGNAL Logical_Operator_out8999_out1            : std_logic;
  SIGNAL Logical_Operator_out9000_out1            : std_logic;
  SIGNAL Logical_Operator_out9001_out1            : std_logic;
  SIGNAL Logical_Operator_out9002_out1            : std_logic;
  SIGNAL Logical_Operator_out9003_out1            : std_logic;
  SIGNAL Logical_Operator_out9004_out1            : std_logic;
  SIGNAL Logical_Operator_out9005_out1            : std_logic;
  SIGNAL Logical_Operator_out9006_out1            : std_logic;
  SIGNAL Logical_Operator_out9007_out1            : std_logic;
  SIGNAL Logical_Operator_out9008_out1            : std_logic;
  SIGNAL Logical_Operator_out9009_out1            : std_logic;
  SIGNAL Logical_Operator_out9010_out1            : std_logic;
  SIGNAL Logical_Operator_out9011_out1            : std_logic;
  SIGNAL Logical_Operator_out9012_out1            : std_logic;
  SIGNAL Logical_Operator_out9013_out1            : std_logic;
  SIGNAL Logical_Operator_out9014_out1            : std_logic;
  SIGNAL Logical_Operator_out9015_out1            : std_logic;
  SIGNAL Logical_Operator_out9016_out1            : std_logic;
  SIGNAL Logical_Operator_out9017_out1            : std_logic;
  SIGNAL Logical_Operator_out9018_out1            : std_logic;
  SIGNAL Logical_Operator_out9019_out1            : std_logic;
  SIGNAL Logical_Operator_out9020_out1            : std_logic;
  SIGNAL Logical_Operator_out9021_out1            : std_logic;
  SIGNAL Logical_Operator_out9022_out1            : std_logic;
  SIGNAL Logical_Operator_out9023_out1            : std_logic;
  SIGNAL Logical_Operator_out9024_out1            : std_logic;
  SIGNAL Logical_Operator_out9025_out1            : std_logic;
  SIGNAL Logical_Operator_out9026_out1            : std_logic;
  SIGNAL Logical_Operator_out9027_out1            : std_logic;
  SIGNAL Logical_Operator_out9028_out1            : std_logic;
  SIGNAL Logical_Operator_out9029_out1            : std_logic;
  SIGNAL Logical_Operator_out9030_out1            : std_logic;
  SIGNAL Logical_Operator_out9031_out1            : std_logic;
  SIGNAL Logical_Operator_out9032_out1            : std_logic;
  SIGNAL Logical_Operator_out9033_out1            : std_logic;
  SIGNAL Logical_Operator_out9034_out1            : std_logic;
  SIGNAL Logical_Operator_out9035_out1            : std_logic;
  SIGNAL Logical_Operator_out9036_out1            : std_logic;
  SIGNAL Logical_Operator_out9037_out1            : std_logic;
  SIGNAL Logical_Operator_out9038_out1            : std_logic;
  SIGNAL Logical_Operator_out9039_out1            : std_logic;
  SIGNAL Logical_Operator_out9040_out1            : std_logic;
  SIGNAL Logical_Operator_out9041_out1            : std_logic;
  SIGNAL Logical_Operator_out9042_out1            : std_logic;
  SIGNAL Logical_Operator_out9043_out1            : std_logic;
  SIGNAL Logical_Operator_out9044_out1            : std_logic;
  SIGNAL Logical_Operator_out9045_out1            : std_logic;
  SIGNAL Logical_Operator_out9046_out1            : std_logic;
  SIGNAL Logical_Operator_out9047_out1            : std_logic;
  SIGNAL Logical_Operator_out9048_out1            : std_logic;
  SIGNAL Logical_Operator_out9049_out1            : std_logic;
  SIGNAL Logical_Operator_out9050_out1            : std_logic;
  SIGNAL Logical_Operator_out9051_out1            : std_logic;
  SIGNAL Logical_Operator_out9052_out1            : std_logic;
  SIGNAL Logical_Operator_out9053_out1            : std_logic;
  SIGNAL Logical_Operator_out9054_out1            : std_logic;
  SIGNAL Logical_Operator_out9055_out1            : std_logic;
  SIGNAL Logical_Operator_out9056_out1            : std_logic;
  SIGNAL Logical_Operator_out9057_out1            : std_logic;
  SIGNAL Logical_Operator_out9058_out1            : std_logic;
  SIGNAL Logical_Operator_out9059_out1            : std_logic;
  SIGNAL Logical_Operator_out9060_out1            : std_logic;
  SIGNAL Logical_Operator_out9061_out1            : std_logic;
  SIGNAL Logical_Operator_out9062_out1            : std_logic;
  SIGNAL Logical_Operator_out9063_out1            : std_logic;
  SIGNAL Logical_Operator_out9064_out1            : std_logic;
  SIGNAL Logical_Operator_out9065_out1            : std_logic;
  SIGNAL Logical_Operator_out9066_out1            : std_logic;
  SIGNAL Logical_Operator_out9067_out1            : std_logic;
  SIGNAL Logical_Operator_out9068_out1            : std_logic;
  SIGNAL Logical_Operator_out9069_out1            : std_logic;
  SIGNAL Logical_Operator_out9070_out1            : std_logic;
  SIGNAL Logical_Operator_out9071_out1            : std_logic;
  SIGNAL Logical_Operator_out9072_out1            : std_logic;
  SIGNAL Logical_Operator_out9073_out1            : std_logic;
  SIGNAL Logical_Operator_out9074_out1            : std_logic;
  SIGNAL Logical_Operator_out9075_out1            : std_logic;
  SIGNAL Logical_Operator_out9076_out1            : std_logic;
  SIGNAL Logical_Operator_out9077_out1            : std_logic;
  SIGNAL Logical_Operator_out9078_out1            : std_logic;
  SIGNAL Logical_Operator_out9079_out1            : std_logic;
  SIGNAL Logical_Operator_out9080_out1            : std_logic;
  SIGNAL Logical_Operator_out9081_out1            : std_logic;
  SIGNAL Logical_Operator_out9082_out1            : std_logic;
  SIGNAL Logical_Operator_out9083_out1            : std_logic;
  SIGNAL Logical_Operator_out9084_out1            : std_logic;
  SIGNAL Logical_Operator_out9085_out1            : std_logic;
  SIGNAL Logical_Operator_out9086_out1            : std_logic;
  SIGNAL Logical_Operator_out9087_out1            : std_logic;
  SIGNAL Logical_Operator_out9088_out1            : std_logic;
  SIGNAL Logical_Operator_out9089_out1            : std_logic;
  SIGNAL Logical_Operator_out9090_out1            : std_logic;
  SIGNAL Logical_Operator_out9091_out1            : std_logic;
  SIGNAL Logical_Operator_out9092_out1            : std_logic;
  SIGNAL Logical_Operator_out9093_out1            : std_logic;
  SIGNAL Logical_Operator_out9094_out1            : std_logic;
  SIGNAL Logical_Operator_out9095_out1            : std_logic;
  SIGNAL Logical_Operator_out9096_out1            : std_logic;
  SIGNAL Logical_Operator_out9097_out1            : std_logic;
  SIGNAL Logical_Operator_out9098_out1            : std_logic;
  SIGNAL Logical_Operator_out9099_out1            : std_logic;
  SIGNAL Logical_Operator_out9100_out1            : std_logic;
  SIGNAL Logical_Operator_out9101_out1            : std_logic;
  SIGNAL Logical_Operator_out9102_out1            : std_logic;
  SIGNAL Logical_Operator_out9103_out1            : std_logic;
  SIGNAL Logical_Operator_out9104_out1            : std_logic;
  SIGNAL Logical_Operator_out9105_out1            : std_logic;
  SIGNAL Logical_Operator_out9106_out1            : std_logic;
  SIGNAL Logical_Operator_out9107_out1            : std_logic;
  SIGNAL Logical_Operator_out9108_out1            : std_logic;
  SIGNAL Logical_Operator_out9109_out1            : std_logic;
  SIGNAL Logical_Operator_out9110_out1            : std_logic;
  SIGNAL Logical_Operator_out9111_out1            : std_logic;
  SIGNAL Logical_Operator_out9112_out1            : std_logic;
  SIGNAL Logical_Operator_out9113_out1            : std_logic;
  SIGNAL Logical_Operator_out9114_out1            : std_logic;
  SIGNAL Logical_Operator_out9115_out1            : std_logic;
  SIGNAL Logical_Operator_out9116_out1            : std_logic;
  SIGNAL Logical_Operator_out9117_out1            : std_logic;
  SIGNAL Logical_Operator_out9118_out1            : std_logic;
  SIGNAL Logical_Operator_out9119_out1            : std_logic;
  SIGNAL Logical_Operator_out9120_out1            : std_logic;
  SIGNAL Logical_Operator_out9121_out1            : std_logic;
  SIGNAL Logical_Operator_out9122_out1            : std_logic;
  SIGNAL Logical_Operator_out9123_out1            : std_logic;
  SIGNAL Logical_Operator_out9124_out1            : std_logic;
  SIGNAL Logical_Operator_out9125_out1            : std_logic;
  SIGNAL Logical_Operator_out9126_out1            : std_logic;
  SIGNAL Logical_Operator_out9127_out1            : std_logic;
  SIGNAL Logical_Operator_out9128_out1            : std_logic;
  SIGNAL Logical_Operator_out9129_out1            : std_logic;
  SIGNAL Logical_Operator_out9130_out1            : std_logic;
  SIGNAL Logical_Operator_out9131_out1            : std_logic;
  SIGNAL Logical_Operator_out9132_out1            : std_logic;
  SIGNAL Logical_Operator_out9133_out1            : std_logic;
  SIGNAL Logical_Operator_out9134_out1            : std_logic;
  SIGNAL Logical_Operator_out9135_out1            : std_logic;
  SIGNAL Logical_Operator_out9136_out1            : std_logic;
  SIGNAL Logical_Operator_out9137_out1            : std_logic;
  SIGNAL Logical_Operator_out9138_out1            : std_logic;
  SIGNAL Logical_Operator_out9139_out1            : std_logic;
  SIGNAL Logical_Operator_out9140_out1            : std_logic;
  SIGNAL Logical_Operator_out9141_out1            : std_logic;
  SIGNAL Logical_Operator_out9142_out1            : std_logic;
  SIGNAL Logical_Operator_out9143_out1            : std_logic;
  SIGNAL Logical_Operator_out9144_out1            : std_logic;
  SIGNAL Logical_Operator_out9145_out1            : std_logic;
  SIGNAL Logical_Operator_out9146_out1            : std_logic;
  SIGNAL Logical_Operator_out9147_out1            : std_logic;
  SIGNAL Logical_Operator_out9148_out1            : std_logic;
  SIGNAL Logical_Operator_out9149_out1            : std_logic;
  SIGNAL Logical_Operator_out9150_out1            : std_logic;
  SIGNAL Logical_Operator_out9151_out1            : std_logic;
  SIGNAL Logical_Operator_out9152_out1            : std_logic;
  SIGNAL Logical_Operator_out9153_out1            : std_logic;
  SIGNAL Logical_Operator_out9154_out1            : std_logic;
  SIGNAL Logical_Operator_out9155_out1            : std_logic;
  SIGNAL Logical_Operator_out9156_out1            : std_logic;
  SIGNAL Logical_Operator_out9157_out1            : std_logic;
  SIGNAL Logical_Operator_out9158_out1            : std_logic;
  SIGNAL Logical_Operator_out9159_out1            : std_logic;
  SIGNAL Logical_Operator_out9160_out1            : std_logic;
  SIGNAL Logical_Operator_out9161_out1            : std_logic;
  SIGNAL Logical_Operator_out9162_out1            : std_logic;
  SIGNAL Logical_Operator_out9163_out1            : std_logic;
  SIGNAL Logical_Operator_out9164_out1            : std_logic;
  SIGNAL Logical_Operator_out9165_out1            : std_logic;
  SIGNAL Logical_Operator_out9166_out1            : std_logic;
  SIGNAL Logical_Operator_out9167_out1            : std_logic;
  SIGNAL Logical_Operator_out9168_out1            : std_logic;
  SIGNAL Logical_Operator_out9169_out1            : std_logic;
  SIGNAL Logical_Operator_out9170_out1            : std_logic;
  SIGNAL Logical_Operator_out9171_out1            : std_logic;
  SIGNAL Logical_Operator_out9172_out1            : std_logic;
  SIGNAL Logical_Operator_out9173_out1            : std_logic;
  SIGNAL Logical_Operator_out9174_out1            : std_logic;
  SIGNAL Logical_Operator_out9175_out1            : std_logic;
  SIGNAL Logical_Operator_out9176_out1            : std_logic;
  SIGNAL Logical_Operator_out9177_out1            : std_logic;
  SIGNAL Logical_Operator_out9178_out1            : std_logic;
  SIGNAL Logical_Operator_out9179_out1            : std_logic;
  SIGNAL Logical_Operator_out9180_out1            : std_logic;
  SIGNAL Logical_Operator_out9181_out1            : std_logic;
  SIGNAL Logical_Operator_out9182_out1            : std_logic;
  SIGNAL Logical_Operator_out9183_out1            : std_logic;
  SIGNAL Logical_Operator_out9184_out1            : std_logic;
  SIGNAL Logical_Operator_out9185_out1            : std_logic;
  SIGNAL Logical_Operator_out9186_out1            : std_logic;
  SIGNAL Logical_Operator_out9187_out1            : std_logic;
  SIGNAL Logical_Operator_out9188_out1            : std_logic;
  SIGNAL Logical_Operator_out9189_out1            : std_logic;
  SIGNAL Logical_Operator_out9190_out1            : std_logic;
  SIGNAL Logical_Operator_out9191_out1            : std_logic;
  SIGNAL Logical_Operator_out9192_out1            : std_logic;
  SIGNAL Logical_Operator_out9193_out1            : std_logic;
  SIGNAL Logical_Operator_out9194_out1            : std_logic;
  SIGNAL Logical_Operator_out9195_out1            : std_logic;
  SIGNAL Logical_Operator_out9196_out1            : std_logic;
  SIGNAL Logical_Operator_out9197_out1            : std_logic;
  SIGNAL Logical_Operator_out9198_out1            : std_logic;
  SIGNAL Logical_Operator_out9199_out1            : std_logic;
  SIGNAL Logical_Operator_out9200_out1            : std_logic;
  SIGNAL Logical_Operator_out9201_out1            : std_logic;
  SIGNAL Logical_Operator_out9202_out1            : std_logic;
  SIGNAL Logical_Operator_out9203_out1            : std_logic;
  SIGNAL Logical_Operator_out9204_out1            : std_logic;
  SIGNAL Logical_Operator_out9205_out1            : std_logic;
  SIGNAL Logical_Operator_out9206_out1            : std_logic;
  SIGNAL Logical_Operator_out9207_out1            : std_logic;
  SIGNAL Logical_Operator_out9208_out1            : std_logic;
  SIGNAL Logical_Operator_out9209_out1            : std_logic;
  SIGNAL Logical_Operator_out9210_out1            : std_logic;
  SIGNAL Logical_Operator_out9211_out1            : std_logic;
  SIGNAL Logical_Operator_out9212_out1            : std_logic;
  SIGNAL Logical_Operator_out9213_out1            : std_logic;
  SIGNAL Logical_Operator_out9214_out1            : std_logic;
  SIGNAL Logical_Operator_out9215_out1            : std_logic;
  SIGNAL Logical_Operator_out9216_out1            : std_logic;
  SIGNAL Logical_Operator_out9217_out1            : std_logic;
  SIGNAL Logical_Operator_out9218_out1            : std_logic;
  SIGNAL Logical_Operator_out9219_out1            : std_logic;
  SIGNAL Logical_Operator_out9220_out1            : std_logic;
  SIGNAL Logical_Operator_out9221_out1            : std_logic;
  SIGNAL Logical_Operator_out9222_out1            : std_logic;
  SIGNAL Logical_Operator_out9223_out1            : std_logic;
  SIGNAL Logical_Operator_out9224_out1            : std_logic;
  SIGNAL Logical_Operator_out9225_out1            : std_logic;
  SIGNAL Logical_Operator_out9226_out1            : std_logic;
  SIGNAL Logical_Operator_out9227_out1            : std_logic;
  SIGNAL Logical_Operator_out9228_out1            : std_logic;
  SIGNAL Logical_Operator_out9229_out1            : std_logic;
  SIGNAL Logical_Operator_out9230_out1            : std_logic;
  SIGNAL Logical_Operator_out9231_out1            : std_logic;
  SIGNAL Logical_Operator_out9232_out1            : std_logic;
  SIGNAL Logical_Operator_out9233_out1            : std_logic;
  SIGNAL Logical_Operator_out9234_out1            : std_logic;
  SIGNAL Logical_Operator_out9235_out1            : std_logic;
  SIGNAL Logical_Operator_out9236_out1            : std_logic;
  SIGNAL Logical_Operator_out9237_out1            : std_logic;
  SIGNAL Logical_Operator_out9238_out1            : std_logic;
  SIGNAL Logical_Operator_out9239_out1            : std_logic;
  SIGNAL Logical_Operator_out9240_out1            : std_logic;
  SIGNAL Logical_Operator_out9241_out1            : std_logic;
  SIGNAL Logical_Operator_out9242_out1            : std_logic;
  SIGNAL Logical_Operator_out9243_out1            : std_logic;
  SIGNAL Logical_Operator_out9244_out1            : std_logic;
  SIGNAL Logical_Operator_out9245_out1            : std_logic;
  SIGNAL Logical_Operator_out9246_out1            : std_logic;
  SIGNAL Logical_Operator_out9247_out1            : std_logic;
  SIGNAL Logical_Operator_out9248_out1            : std_logic;
  SIGNAL Logical_Operator_out9249_out1            : std_logic;
  SIGNAL Logical_Operator_out9250_out1            : std_logic;
  SIGNAL Logical_Operator_out9251_out1            : std_logic;
  SIGNAL Logical_Operator_out9252_out1            : std_logic;
  SIGNAL Logical_Operator_out9253_out1            : std_logic;
  SIGNAL Logical_Operator_out9254_out1            : std_logic;
  SIGNAL Logical_Operator_out9255_out1            : std_logic;
  SIGNAL Logical_Operator_out9256_out1            : std_logic;
  SIGNAL Logical_Operator_out9257_out1            : std_logic;
  SIGNAL Logical_Operator_out9258_out1            : std_logic;
  SIGNAL Logical_Operator_out9259_out1            : std_logic;
  SIGNAL Logical_Operator_out9260_out1            : std_logic;
  SIGNAL Logical_Operator_out9261_out1            : std_logic;
  SIGNAL Logical_Operator_out9262_out1            : std_logic;
  SIGNAL Logical_Operator_out9263_out1            : std_logic;
  SIGNAL Logical_Operator_out9264_out1            : std_logic;
  SIGNAL Logical_Operator_out9265_out1            : std_logic;
  SIGNAL Logical_Operator_out9266_out1            : std_logic;
  SIGNAL Logical_Operator_out9267_out1            : std_logic;
  SIGNAL Logical_Operator_out9268_out1            : std_logic;
  SIGNAL Logical_Operator_out9269_out1            : std_logic;
  SIGNAL Logical_Operator_out9270_out1            : std_logic;
  SIGNAL Logical_Operator_out9271_out1            : std_logic;
  SIGNAL Logical_Operator_out9272_out1            : std_logic;
  SIGNAL Logical_Operator_out9273_out1            : std_logic;
  SIGNAL Logical_Operator_out9274_out1            : std_logic;
  SIGNAL Logical_Operator_out9275_out1            : std_logic;
  SIGNAL Logical_Operator_out9276_out1            : std_logic;
  SIGNAL Logical_Operator_out9277_out1            : std_logic;
  SIGNAL Logical_Operator_out9278_out1            : std_logic;
  SIGNAL Logical_Operator_out9279_out1            : std_logic;
  SIGNAL Logical_Operator_out9280_out1            : std_logic;
  SIGNAL Logical_Operator_out9281_out1            : std_logic;
  SIGNAL Logical_Operator_out9282_out1            : std_logic;
  SIGNAL Logical_Operator_out9283_out1            : std_logic;
  SIGNAL Logical_Operator_out9284_out1            : std_logic;
  SIGNAL Logical_Operator_out9285_out1            : std_logic;
  SIGNAL Logical_Operator_out9286_out1            : std_logic;
  SIGNAL Logical_Operator_out9287_out1            : std_logic;
  SIGNAL Logical_Operator_out9288_out1            : std_logic;
  SIGNAL Logical_Operator_out9289_out1            : std_logic;
  SIGNAL Logical_Operator_out9290_out1            : std_logic;
  SIGNAL Logical_Operator_out9291_out1            : std_logic;
  SIGNAL Logical_Operator_out9292_out1            : std_logic;
  SIGNAL Logical_Operator_out9293_out1            : std_logic;
  SIGNAL Logical_Operator_out9294_out1            : std_logic;
  SIGNAL Logical_Operator_out9295_out1            : std_logic;
  SIGNAL Logical_Operator_out9296_out1            : std_logic;
  SIGNAL Logical_Operator_out9297_out1            : std_logic;
  SIGNAL Logical_Operator_out9298_out1            : std_logic;
  SIGNAL Logical_Operator_out9299_out1            : std_logic;
  SIGNAL Logical_Operator_out9300_out1            : std_logic;
  SIGNAL Logical_Operator_out9301_out1            : std_logic;
  SIGNAL Logical_Operator_out9302_out1            : std_logic;
  SIGNAL Logical_Operator_out9303_out1            : std_logic;
  SIGNAL Logical_Operator_out9304_out1            : std_logic;
  SIGNAL Logical_Operator_out9305_out1            : std_logic;
  SIGNAL Logical_Operator_out9306_out1            : std_logic;
  SIGNAL Logical_Operator_out9307_out1            : std_logic;
  SIGNAL Logical_Operator_out9308_out1            : std_logic;
  SIGNAL Logical_Operator_out9309_out1            : std_logic;
  SIGNAL Logical_Operator_out9310_out1            : std_logic;
  SIGNAL Logical_Operator_out9311_out1            : std_logic;
  SIGNAL Logical_Operator_out9312_out1            : std_logic;
  SIGNAL Logical_Operator_out9313_out1            : std_logic;
  SIGNAL Logical_Operator_out9314_out1            : std_logic;
  SIGNAL Logical_Operator_out9315_out1            : std_logic;
  SIGNAL Logical_Operator_out9316_out1            : std_logic;
  SIGNAL Logical_Operator_out9317_out1            : std_logic;
  SIGNAL Logical_Operator_out9318_out1            : std_logic;
  SIGNAL Logical_Operator_out9319_out1            : std_logic;
  SIGNAL Logical_Operator_out9320_out1            : std_logic;
  SIGNAL Logical_Operator_out9321_out1            : std_logic;
  SIGNAL Logical_Operator_out9322_out1            : std_logic;
  SIGNAL Logical_Operator_out9323_out1            : std_logic;
  SIGNAL Logical_Operator_out9324_out1            : std_logic;
  SIGNAL Logical_Operator_out9325_out1            : std_logic;
  SIGNAL Logical_Operator_out9326_out1            : std_logic;
  SIGNAL Logical_Operator_out9327_out1            : std_logic;
  SIGNAL Logical_Operator_out9328_out1            : std_logic;
  SIGNAL Logical_Operator_out9329_out1            : std_logic;
  SIGNAL Logical_Operator_out9330_out1            : std_logic;
  SIGNAL Logical_Operator_out9331_out1            : std_logic;
  SIGNAL Logical_Operator_out9332_out1            : std_logic;
  SIGNAL Logical_Operator_out9333_out1            : std_logic;
  SIGNAL Logical_Operator_out9334_out1            : std_logic;
  SIGNAL Logical_Operator_out9335_out1            : std_logic;
  SIGNAL Logical_Operator_out9336_out1            : std_logic;
  SIGNAL Logical_Operator_out9337_out1            : std_logic;
  SIGNAL Logical_Operator_out9338_out1            : std_logic;
  SIGNAL Logical_Operator_out9339_out1            : std_logic;
  SIGNAL Logical_Operator_out9340_out1            : std_logic;
  SIGNAL Logical_Operator_out9341_out1            : std_logic;
  SIGNAL Logical_Operator_out9342_out1            : std_logic;
  SIGNAL Logical_Operator_out9343_out1            : std_logic;
  SIGNAL Logical_Operator_out9344_out1            : std_logic;
  SIGNAL Logical_Operator_out9345_out1            : std_logic;
  SIGNAL Logical_Operator_out9346_out1            : std_logic;
  SIGNAL Logical_Operator_out9347_out1            : std_logic;
  SIGNAL Logical_Operator_out9348_out1            : std_logic;
  SIGNAL Logical_Operator_out9349_out1            : std_logic;
  SIGNAL Logical_Operator_out9350_out1            : std_logic;
  SIGNAL Logical_Operator_out9351_out1            : std_logic;
  SIGNAL Logical_Operator_out9352_out1            : std_logic;
  SIGNAL Logical_Operator_out9353_out1            : std_logic;
  SIGNAL Logical_Operator_out9354_out1            : std_logic;
  SIGNAL Logical_Operator_out9355_out1            : std_logic;
  SIGNAL Logical_Operator_out9356_out1            : std_logic;
  SIGNAL Logical_Operator_out9357_out1            : std_logic;
  SIGNAL Logical_Operator_out9358_out1            : std_logic;
  SIGNAL Logical_Operator_out9359_out1            : std_logic;
  SIGNAL Logical_Operator_out9360_out1            : std_logic;
  SIGNAL Logical_Operator_out9361_out1            : std_logic;
  SIGNAL Logical_Operator_out9362_out1            : std_logic;
  SIGNAL Logical_Operator_out9363_out1            : std_logic;
  SIGNAL Logical_Operator_out9364_out1            : std_logic;
  SIGNAL Logical_Operator_out9365_out1            : std_logic;
  SIGNAL Logical_Operator_out9366_out1            : std_logic;
  SIGNAL Logical_Operator_out9367_out1            : std_logic;
  SIGNAL Logical_Operator_out9368_out1            : std_logic;
  SIGNAL Logical_Operator_out9369_out1            : std_logic;
  SIGNAL Logical_Operator_out9370_out1            : std_logic;
  SIGNAL Logical_Operator_out9371_out1            : std_logic;
  SIGNAL Logical_Operator_out9372_out1            : std_logic;
  SIGNAL Logical_Operator_out9373_out1            : std_logic;
  SIGNAL Logical_Operator_out9374_out1            : std_logic;
  SIGNAL Logical_Operator_out9375_out1            : std_logic;
  SIGNAL Logical_Operator_out9376_out1            : std_logic;
  SIGNAL Logical_Operator_out9377_out1            : std_logic;
  SIGNAL Logical_Operator_out9378_out1            : std_logic;
  SIGNAL Logical_Operator_out9379_out1            : std_logic;
  SIGNAL Logical_Operator_out9380_out1            : std_logic;
  SIGNAL Logical_Operator_out9381_out1            : std_logic;
  SIGNAL Logical_Operator_out9382_out1            : std_logic;
  SIGNAL Logical_Operator_out9383_out1            : std_logic;
  SIGNAL Logical_Operator_out9384_out1            : std_logic;
  SIGNAL Logical_Operator_out9385_out1            : std_logic;
  SIGNAL Logical_Operator_out9386_out1            : std_logic;
  SIGNAL Logical_Operator_out9387_out1            : std_logic;
  SIGNAL Logical_Operator_out9388_out1            : std_logic;
  SIGNAL Logical_Operator_out9389_out1            : std_logic;
  SIGNAL Logical_Operator_out9390_out1            : std_logic;
  SIGNAL Logical_Operator_out9391_out1            : std_logic;
  SIGNAL Logical_Operator_out9392_out1            : std_logic;
  SIGNAL Logical_Operator_out9393_out1            : std_logic;
  SIGNAL Logical_Operator_out9394_out1            : std_logic;
  SIGNAL Logical_Operator_out9395_out1            : std_logic;
  SIGNAL Logical_Operator_out9396_out1            : std_logic;
  SIGNAL Logical_Operator_out9397_out1            : std_logic;
  SIGNAL Logical_Operator_out9398_out1            : std_logic;
  SIGNAL Logical_Operator_out9399_out1            : std_logic;
  SIGNAL Logical_Operator_out9400_out1            : std_logic;
  SIGNAL Logical_Operator_out9401_out1            : std_logic;
  SIGNAL Logical_Operator_out9402_out1            : std_logic;
  SIGNAL Logical_Operator_out9403_out1            : std_logic;
  SIGNAL Logical_Operator_out9404_out1            : std_logic;
  SIGNAL Logical_Operator_out9405_out1            : std_logic;
  SIGNAL Logical_Operator_out9406_out1            : std_logic;
  SIGNAL Logical_Operator_out9407_out1            : std_logic;
  SIGNAL Logical_Operator_out9408_out1            : std_logic;
  SIGNAL Logical_Operator_out9409_out1            : std_logic;
  SIGNAL Logical_Operator_out9410_out1            : std_logic;
  SIGNAL Logical_Operator_out9411_out1            : std_logic;
  SIGNAL Logical_Operator_out9412_out1            : std_logic;
  SIGNAL Logical_Operator_out9413_out1            : std_logic;
  SIGNAL Logical_Operator_out9414_out1            : std_logic;
  SIGNAL Logical_Operator_out9415_out1            : std_logic;
  SIGNAL Logical_Operator_out9416_out1            : std_logic;
  SIGNAL Logical_Operator_out9417_out1            : std_logic;
  SIGNAL Logical_Operator_out9418_out1            : std_logic;
  SIGNAL Logical_Operator_out9419_out1            : std_logic;
  SIGNAL Logical_Operator_out9420_out1            : std_logic;
  SIGNAL Logical_Operator_out9421_out1            : std_logic;
  SIGNAL Logical_Operator_out9422_out1            : std_logic;
  SIGNAL Logical_Operator_out9423_out1            : std_logic;
  SIGNAL Logical_Operator_out9424_out1            : std_logic;
  SIGNAL Logical_Operator_out9425_out1            : std_logic;
  SIGNAL Logical_Operator_out9426_out1            : std_logic;
  SIGNAL Logical_Operator_out9427_out1            : std_logic;
  SIGNAL Logical_Operator_out9428_out1            : std_logic;
  SIGNAL Logical_Operator_out9429_out1            : std_logic;
  SIGNAL Logical_Operator_out9430_out1            : std_logic;
  SIGNAL Logical_Operator_out9431_out1            : std_logic;
  SIGNAL Logical_Operator_out9432_out1            : std_logic;
  SIGNAL Logical_Operator_out9433_out1            : std_logic;
  SIGNAL Logical_Operator_out9434_out1            : std_logic;
  SIGNAL Logical_Operator_out9435_out1            : std_logic;
  SIGNAL Logical_Operator_out9436_out1            : std_logic;
  SIGNAL Logical_Operator_out9437_out1            : std_logic;
  SIGNAL Logical_Operator_out9438_out1            : std_logic;
  SIGNAL Logical_Operator_out9439_out1            : std_logic;
  SIGNAL Logical_Operator_out9440_out1            : std_logic;
  SIGNAL Logical_Operator_out9441_out1            : std_logic;
  SIGNAL Logical_Operator_out9442_out1            : std_logic;
  SIGNAL Logical_Operator_out9443_out1            : std_logic;
  SIGNAL Logical_Operator_out9444_out1            : std_logic;
  SIGNAL Logical_Operator_out9445_out1            : std_logic;
  SIGNAL Logical_Operator_out9446_out1            : std_logic;
  SIGNAL Logical_Operator_out9447_out1            : std_logic;
  SIGNAL Logical_Operator_out9448_out1            : std_logic;
  SIGNAL Logical_Operator_out9449_out1            : std_logic;
  SIGNAL Logical_Operator_out9450_out1            : std_logic;
  SIGNAL Logical_Operator_out9451_out1            : std_logic;
  SIGNAL Logical_Operator_out9452_out1            : std_logic;
  SIGNAL Logical_Operator_out9453_out1            : std_logic;
  SIGNAL Logical_Operator_out9454_out1            : std_logic;
  SIGNAL Logical_Operator_out9455_out1            : std_logic;
  SIGNAL Logical_Operator_out9456_out1            : std_logic;
  SIGNAL Logical_Operator_out9457_out1            : std_logic;
  SIGNAL Logical_Operator_out9458_out1            : std_logic;
  SIGNAL Logical_Operator_out9459_out1            : std_logic;
  SIGNAL Logical_Operator_out9460_out1            : std_logic;
  SIGNAL Logical_Operator_out9461_out1            : std_logic;
  SIGNAL Logical_Operator_out9462_out1            : std_logic;
  SIGNAL Logical_Operator_out9463_out1            : std_logic;
  SIGNAL Logical_Operator_out9464_out1            : std_logic;
  SIGNAL Logical_Operator_out9465_out1            : std_logic;
  SIGNAL Logical_Operator_out9466_out1            : std_logic;
  SIGNAL Logical_Operator_out9467_out1            : std_logic;
  SIGNAL Logical_Operator_out9468_out1            : std_logic;
  SIGNAL Logical_Operator_out9469_out1            : std_logic;
  SIGNAL Logical_Operator_out9470_out1            : std_logic;
  SIGNAL Logical_Operator_out9471_out1            : std_logic;
  SIGNAL Logical_Operator_out9472_out1            : std_logic;
  SIGNAL Logical_Operator_out9473_out1            : std_logic;
  SIGNAL Logical_Operator_out9474_out1            : std_logic;
  SIGNAL Logical_Operator_out9475_out1            : std_logic;
  SIGNAL Logical_Operator_out9476_out1            : std_logic;
  SIGNAL Logical_Operator_out9477_out1            : std_logic;
  SIGNAL Logical_Operator_out9478_out1            : std_logic;
  SIGNAL Logical_Operator_out9479_out1            : std_logic;
  SIGNAL Logical_Operator_out9480_out1            : std_logic;
  SIGNAL Logical_Operator_out9481_out1            : std_logic;
  SIGNAL Logical_Operator_out9482_out1            : std_logic;
  SIGNAL Logical_Operator_out9483_out1            : std_logic;
  SIGNAL Logical_Operator_out9484_out1            : std_logic;
  SIGNAL Logical_Operator_out9485_out1            : std_logic;
  SIGNAL Logical_Operator_out9486_out1            : std_logic;
  SIGNAL Logical_Operator_out9487_out1            : std_logic;
  SIGNAL Logical_Operator_out9488_out1            : std_logic;
  SIGNAL Logical_Operator_out9489_out1            : std_logic;
  SIGNAL Logical_Operator_out9490_out1            : std_logic;
  SIGNAL Logical_Operator_out9491_out1            : std_logic;
  SIGNAL Logical_Operator_out9492_out1            : std_logic;
  SIGNAL Logical_Operator_out9493_out1            : std_logic;
  SIGNAL Logical_Operator_out9494_out1            : std_logic;
  SIGNAL Logical_Operator_out9495_out1            : std_logic;
  SIGNAL Logical_Operator_out9496_out1            : std_logic;
  SIGNAL Logical_Operator_out9497_out1            : std_logic;
  SIGNAL Logical_Operator_out9498_out1            : std_logic;
  SIGNAL Logical_Operator_out9499_out1            : std_logic;
  SIGNAL Logical_Operator_out9500_out1            : std_logic;
  SIGNAL Logical_Operator_out9501_out1            : std_logic;
  SIGNAL Logical_Operator_out9502_out1            : std_logic;
  SIGNAL Logical_Operator_out9503_out1            : std_logic;
  SIGNAL Logical_Operator_out9504_out1            : std_logic;
  SIGNAL Logical_Operator_out9505_out1            : std_logic;
  SIGNAL Logical_Operator_out9506_out1            : std_logic;
  SIGNAL Logical_Operator_out9507_out1            : std_logic;
  SIGNAL Logical_Operator_out9508_out1            : std_logic;
  SIGNAL Logical_Operator_out9509_out1            : std_logic;
  SIGNAL Logical_Operator_out9510_out1            : std_logic;
  SIGNAL Logical_Operator_out9511_out1            : std_logic;
  SIGNAL Logical_Operator_out9512_out1            : std_logic;
  SIGNAL Logical_Operator_out9513_out1            : std_logic;
  SIGNAL Logical_Operator_out9514_out1            : std_logic;
  SIGNAL Logical_Operator_out9515_out1            : std_logic;
  SIGNAL Logical_Operator_out9516_out1            : std_logic;
  SIGNAL Logical_Operator_out9517_out1            : std_logic;
  SIGNAL Logical_Operator_out9518_out1            : std_logic;
  SIGNAL Logical_Operator_out9519_out1            : std_logic;
  SIGNAL Logical_Operator_out9520_out1            : std_logic;
  SIGNAL Logical_Operator_out9521_out1            : std_logic;
  SIGNAL Logical_Operator_out9522_out1            : std_logic;
  SIGNAL Logical_Operator_out9523_out1            : std_logic;
  SIGNAL Logical_Operator_out9524_out1            : std_logic;
  SIGNAL Logical_Operator_out9525_out1            : std_logic;
  SIGNAL Logical_Operator_out9526_out1            : std_logic;
  SIGNAL Logical_Operator_out9527_out1            : std_logic;
  SIGNAL Logical_Operator_out9528_out1            : std_logic;
  SIGNAL Logical_Operator_out9529_out1            : std_logic;
  SIGNAL Logical_Operator_out9530_out1            : std_logic;
  SIGNAL Logical_Operator_out9531_out1            : std_logic;
  SIGNAL Logical_Operator_out9532_out1            : std_logic;
  SIGNAL Logical_Operator_out9533_out1            : std_logic;
  SIGNAL Logical_Operator_out9534_out1            : std_logic;
  SIGNAL Logical_Operator_out9535_out1            : std_logic;
  SIGNAL Logical_Operator_out9536_out1            : std_logic;
  SIGNAL Logical_Operator_out9537_out1            : std_logic;
  SIGNAL Logical_Operator_out9538_out1            : std_logic;
  SIGNAL Logical_Operator_out9539_out1            : std_logic;
  SIGNAL Logical_Operator_out9540_out1            : std_logic;
  SIGNAL Logical_Operator_out9541_out1            : std_logic;
  SIGNAL Logical_Operator_out9542_out1            : std_logic;
  SIGNAL Logical_Operator_out9543_out1            : std_logic;
  SIGNAL Logical_Operator_out9544_out1            : std_logic;
  SIGNAL Logical_Operator_out9545_out1            : std_logic;
  SIGNAL Logical_Operator_out9546_out1            : std_logic;
  SIGNAL Logical_Operator_out9547_out1            : std_logic;
  SIGNAL Logical_Operator_out9548_out1            : std_logic;
  SIGNAL Logical_Operator_out9549_out1            : std_logic;
  SIGNAL Logical_Operator_out9550_out1            : std_logic;
  SIGNAL Logical_Operator_out9551_out1            : std_logic;
  SIGNAL Logical_Operator_out9552_out1            : std_logic;
  SIGNAL Logical_Operator_out9553_out1            : std_logic;
  SIGNAL Logical_Operator_out9554_out1            : std_logic;
  SIGNAL Logical_Operator_out9555_out1            : std_logic;
  SIGNAL Logical_Operator_out9556_out1            : std_logic;
  SIGNAL Logical_Operator_out9557_out1            : std_logic;
  SIGNAL Logical_Operator_out9558_out1            : std_logic;
  SIGNAL Logical_Operator_out9559_out1            : std_logic;
  SIGNAL Logical_Operator_out9560_out1            : std_logic;
  SIGNAL Logical_Operator_out9561_out1            : std_logic;
  SIGNAL Logical_Operator_out9562_out1            : std_logic;
  SIGNAL Logical_Operator_out9563_out1            : std_logic;
  SIGNAL Logical_Operator_out9564_out1            : std_logic;
  SIGNAL Logical_Operator_out9565_out1            : std_logic;
  SIGNAL Logical_Operator_out9566_out1            : std_logic;
  SIGNAL Logical_Operator_out9567_out1            : std_logic;
  SIGNAL Logical_Operator_out9568_out1            : std_logic;
  SIGNAL Logical_Operator_out9569_out1            : std_logic;
  SIGNAL Logical_Operator_out9570_out1            : std_logic;
  SIGNAL Logical_Operator_out9571_out1            : std_logic;
  SIGNAL Logical_Operator_out9572_out1            : std_logic;
  SIGNAL Logical_Operator_out9573_out1            : std_logic;
  SIGNAL Logical_Operator_out9574_out1            : std_logic;
  SIGNAL Logical_Operator_out9575_out1            : std_logic;
  SIGNAL Logical_Operator_out9576_out1            : std_logic;
  SIGNAL Logical_Operator_out9577_out1            : std_logic;
  SIGNAL Logical_Operator_out9578_out1            : std_logic;
  SIGNAL Logical_Operator_out9579_out1            : std_logic;
  SIGNAL Logical_Operator_out9580_out1            : std_logic;
  SIGNAL Logical_Operator_out9581_out1            : std_logic;
  SIGNAL Logical_Operator_out9582_out1            : std_logic;
  SIGNAL Logical_Operator_out9583_out1            : std_logic;
  SIGNAL Logical_Operator_out9584_out1            : std_logic;
  SIGNAL Logical_Operator_out9585_out1            : std_logic;
  SIGNAL Logical_Operator_out9586_out1            : std_logic;
  SIGNAL Logical_Operator_out9587_out1            : std_logic;
  SIGNAL Logical_Operator_out9588_out1            : std_logic;
  SIGNAL Logical_Operator_out9589_out1            : std_logic;
  SIGNAL Logical_Operator_out9590_out1            : std_logic;
  SIGNAL Logical_Operator_out9591_out1            : std_logic;
  SIGNAL Logical_Operator_out9592_out1            : std_logic;
  SIGNAL Logical_Operator_out9593_out1            : std_logic;
  SIGNAL Logical_Operator_out9594_out1            : std_logic;
  SIGNAL Logical_Operator_out9595_out1            : std_logic;
  SIGNAL Logical_Operator_out9596_out1            : std_logic;
  SIGNAL Logical_Operator_out9597_out1            : std_logic;
  SIGNAL Logical_Operator_out9598_out1            : std_logic;
  SIGNAL Logical_Operator_out9599_out1            : std_logic;
  SIGNAL Logical_Operator_out9600_out1            : std_logic;
  SIGNAL Logical_Operator_out9601_out1            : std_logic;
  SIGNAL Logical_Operator_out9602_out1            : std_logic;
  SIGNAL Logical_Operator_out9603_out1            : std_logic;
  SIGNAL Logical_Operator_out9604_out1            : std_logic;
  SIGNAL Logical_Operator_out9605_out1            : std_logic;
  SIGNAL Logical_Operator_out9606_out1            : std_logic;
  SIGNAL Logical_Operator_out9607_out1            : std_logic;
  SIGNAL Logical_Operator_out9608_out1            : std_logic;
  SIGNAL Logical_Operator_out9609_out1            : std_logic;
  SIGNAL Logical_Operator_out9610_out1            : std_logic;
  SIGNAL Logical_Operator_out9611_out1            : std_logic;
  SIGNAL Logical_Operator_out9612_out1            : std_logic;
  SIGNAL Logical_Operator_out9613_out1            : std_logic;
  SIGNAL Logical_Operator_out9614_out1            : std_logic;
  SIGNAL Logical_Operator_out9615_out1            : std_logic;
  SIGNAL Logical_Operator_out9616_out1            : std_logic;
  SIGNAL Logical_Operator_out9617_out1            : std_logic;
  SIGNAL Logical_Operator_out9618_out1            : std_logic;
  SIGNAL Logical_Operator_out9619_out1            : std_logic;
  SIGNAL Logical_Operator_out9620_out1            : std_logic;
  SIGNAL Logical_Operator_out9621_out1            : std_logic;
  SIGNAL Logical_Operator_out9622_out1            : std_logic;
  SIGNAL Logical_Operator_out9623_out1            : std_logic;
  SIGNAL Logical_Operator_out9624_out1            : std_logic;
  SIGNAL Logical_Operator_out9625_out1            : std_logic;
  SIGNAL Logical_Operator_out9626_out1            : std_logic;
  SIGNAL Logical_Operator_out9627_out1            : std_logic;
  SIGNAL Logical_Operator_out9628_out1            : std_logic;
  SIGNAL Logical_Operator_out9629_out1            : std_logic;
  SIGNAL Logical_Operator_out9630_out1            : std_logic;
  SIGNAL Logical_Operator_out9631_out1            : std_logic;
  SIGNAL Logical_Operator_out9632_out1            : std_logic;
  SIGNAL Logical_Operator_out9633_out1            : std_logic;
  SIGNAL Logical_Operator_out9634_out1            : std_logic;
  SIGNAL Logical_Operator_out9635_out1            : std_logic;
  SIGNAL Logical_Operator_out9636_out1            : std_logic;
  SIGNAL Logical_Operator_out9637_out1            : std_logic;
  SIGNAL Logical_Operator_out9638_out1            : std_logic;
  SIGNAL Logical_Operator_out9639_out1            : std_logic;
  SIGNAL Logical_Operator_out9640_out1            : std_logic;
  SIGNAL Logical_Operator_out9641_out1            : std_logic;
  SIGNAL Logical_Operator_out9642_out1            : std_logic;
  SIGNAL Logical_Operator_out9643_out1            : std_logic;
  SIGNAL Logical_Operator_out9644_out1            : std_logic;
  SIGNAL Logical_Operator_out9645_out1            : std_logic;
  SIGNAL Logical_Operator_out9646_out1            : std_logic;
  SIGNAL Logical_Operator_out9647_out1            : std_logic;
  SIGNAL Logical_Operator_out9648_out1            : std_logic;
  SIGNAL Logical_Operator_out9649_out1            : std_logic;
  SIGNAL Logical_Operator_out9650_out1            : std_logic;
  SIGNAL Logical_Operator_out9651_out1            : std_logic;
  SIGNAL Logical_Operator_out9652_out1            : std_logic;
  SIGNAL Logical_Operator_out9653_out1            : std_logic;
  SIGNAL Logical_Operator_out9654_out1            : std_logic;
  SIGNAL Logical_Operator_out9655_out1            : std_logic;
  SIGNAL Logical_Operator_out9656_out1            : std_logic;
  SIGNAL Logical_Operator_out9657_out1            : std_logic;
  SIGNAL Logical_Operator_out9658_out1            : std_logic;
  SIGNAL Logical_Operator_out9659_out1            : std_logic;
  SIGNAL Logical_Operator_out9660_out1            : std_logic;
  SIGNAL Logical_Operator_out9661_out1            : std_logic;
  SIGNAL Logical_Operator_out9662_out1            : std_logic;
  SIGNAL Logical_Operator_out9663_out1            : std_logic;
  SIGNAL Logical_Operator_out9664_out1            : std_logic;
  SIGNAL Logical_Operator_out9665_out1            : std_logic;
  SIGNAL Logical_Operator_out9666_out1            : std_logic;
  SIGNAL Logical_Operator_out9667_out1            : std_logic;
  SIGNAL Logical_Operator_out9668_out1            : std_logic;
  SIGNAL Logical_Operator_out9669_out1            : std_logic;
  SIGNAL Logical_Operator_out9670_out1            : std_logic;
  SIGNAL Logical_Operator_out9671_out1            : std_logic;
  SIGNAL Logical_Operator_out9672_out1            : std_logic;
  SIGNAL Logical_Operator_out9673_out1            : std_logic;
  SIGNAL Logical_Operator_out9674_out1            : std_logic;
  SIGNAL Logical_Operator_out9675_out1            : std_logic;
  SIGNAL Logical_Operator_out9676_out1            : std_logic;
  SIGNAL Logical_Operator_out9677_out1            : std_logic;
  SIGNAL Logical_Operator_out9678_out1            : std_logic;
  SIGNAL Logical_Operator_out9679_out1            : std_logic;
  SIGNAL Logical_Operator_out9680_out1            : std_logic;
  SIGNAL Logical_Operator_out9681_out1            : std_logic;
  SIGNAL Logical_Operator_out9682_out1            : std_logic;
  SIGNAL Logical_Operator_out9683_out1            : std_logic;
  SIGNAL Logical_Operator_out9684_out1            : std_logic;
  SIGNAL Logical_Operator_out9685_out1            : std_logic;
  SIGNAL Logical_Operator_out9686_out1            : std_logic;
  SIGNAL Logical_Operator_out9687_out1            : std_logic;
  SIGNAL Logical_Operator_out9688_out1            : std_logic;
  SIGNAL Logical_Operator_out9689_out1            : std_logic;
  SIGNAL Logical_Operator_out9690_out1            : std_logic;
  SIGNAL Logical_Operator_out9691_out1            : std_logic;
  SIGNAL Logical_Operator_out9692_out1            : std_logic;
  SIGNAL Logical_Operator_out9693_out1            : std_logic;
  SIGNAL Logical_Operator_out9694_out1            : std_logic;
  SIGNAL Logical_Operator_out9695_out1            : std_logic;
  SIGNAL Logical_Operator_out9696_out1            : std_logic;
  SIGNAL Logical_Operator_out9697_out1            : std_logic;
  SIGNAL Logical_Operator_out9698_out1            : std_logic;
  SIGNAL Logical_Operator_out9699_out1            : std_logic;
  SIGNAL Logical_Operator_out9700_out1            : std_logic;
  SIGNAL Logical_Operator_out9701_out1            : std_logic;
  SIGNAL Logical_Operator_out9702_out1            : std_logic;
  SIGNAL Logical_Operator_out9703_out1            : std_logic;
  SIGNAL Logical_Operator_out9704_out1            : std_logic;
  SIGNAL Logical_Operator_out9705_out1            : std_logic;
  SIGNAL Logical_Operator_out9706_out1            : std_logic;
  SIGNAL Logical_Operator_out9707_out1            : std_logic;
  SIGNAL Logical_Operator_out9708_out1            : std_logic;
  SIGNAL Logical_Operator_out9709_out1            : std_logic;
  SIGNAL Logical_Operator_out9710_out1            : std_logic;
  SIGNAL Logical_Operator_out9711_out1            : std_logic;
  SIGNAL Logical_Operator_out9712_out1            : std_logic;
  SIGNAL Logical_Operator_out9713_out1            : std_logic;
  SIGNAL Logical_Operator_out9714_out1            : std_logic;
  SIGNAL Logical_Operator_out9715_out1            : std_logic;
  SIGNAL Logical_Operator_out9716_out1            : std_logic;
  SIGNAL Logical_Operator_out9717_out1            : std_logic;
  SIGNAL Logical_Operator_out9718_out1            : std_logic;
  SIGNAL Logical_Operator_out9719_out1            : std_logic;
  SIGNAL Logical_Operator_out9720_out1            : std_logic;
  SIGNAL Logical_Operator_out9721_out1            : std_logic;
  SIGNAL Logical_Operator_out9722_out1            : std_logic;
  SIGNAL Logical_Operator_out9723_out1            : std_logic;
  SIGNAL Logical_Operator_out9724_out1            : std_logic;
  SIGNAL Logical_Operator_out9725_out1            : std_logic;
  SIGNAL Logical_Operator_out9726_out1            : std_logic;
  SIGNAL Logical_Operator_out9727_out1            : std_logic;
  SIGNAL Logical_Operator_out9728_out1            : std_logic;
  SIGNAL Logical_Operator_out9729_out1            : std_logic;
  SIGNAL Logical_Operator_out9730_out1            : std_logic;
  SIGNAL Logical_Operator_out9731_out1            : std_logic;
  SIGNAL Logical_Operator_out9732_out1            : std_logic;
  SIGNAL Logical_Operator_out9733_out1            : std_logic;
  SIGNAL Logical_Operator_out9734_out1            : std_logic;
  SIGNAL Logical_Operator_out9735_out1            : std_logic;
  SIGNAL Logical_Operator_out9736_out1            : std_logic;
  SIGNAL Logical_Operator_out9737_out1            : std_logic;
  SIGNAL Logical_Operator_out9738_out1            : std_logic;
  SIGNAL Logical_Operator_out9739_out1            : std_logic;
  SIGNAL Logical_Operator_out9740_out1            : std_logic;
  SIGNAL Logical_Operator_out9741_out1            : std_logic;
  SIGNAL Logical_Operator_out9742_out1            : std_logic;
  SIGNAL Logical_Operator_out9743_out1            : std_logic;
  SIGNAL Logical_Operator_out9744_out1            : std_logic;
  SIGNAL Logical_Operator_out9745_out1            : std_logic;
  SIGNAL Logical_Operator_out9746_out1            : std_logic;
  SIGNAL Logical_Operator_out9747_out1            : std_logic;
  SIGNAL Logical_Operator_out9748_out1            : std_logic;
  SIGNAL Logical_Operator_out9749_out1            : std_logic;
  SIGNAL Logical_Operator_out9750_out1            : std_logic;
  SIGNAL Logical_Operator_out9751_out1            : std_logic;
  SIGNAL Logical_Operator_out9752_out1            : std_logic;
  SIGNAL Logical_Operator_out9753_out1            : std_logic;
  SIGNAL Logical_Operator_out9754_out1            : std_logic;
  SIGNAL Logical_Operator_out9755_out1            : std_logic;
  SIGNAL Logical_Operator_out9756_out1            : std_logic;
  SIGNAL Logical_Operator_out9757_out1            : std_logic;
  SIGNAL Logical_Operator_out9758_out1            : std_logic;
  SIGNAL Logical_Operator_out9759_out1            : std_logic;
  SIGNAL Logical_Operator_out9760_out1            : std_logic;
  SIGNAL Logical_Operator_out9761_out1            : std_logic;
  SIGNAL Logical_Operator_out9762_out1            : std_logic;
  SIGNAL Logical_Operator_out9763_out1            : std_logic;
  SIGNAL Logical_Operator_out9764_out1            : std_logic;
  SIGNAL Logical_Operator_out9765_out1            : std_logic;
  SIGNAL Logical_Operator_out9766_out1            : std_logic;
  SIGNAL Logical_Operator_out9767_out1            : std_logic;
  SIGNAL Logical_Operator_out9768_out1            : std_logic;
  SIGNAL Logical_Operator_out9769_out1            : std_logic;
  SIGNAL Logical_Operator_out9770_out1            : std_logic;
  SIGNAL Logical_Operator_out9771_out1            : std_logic;
  SIGNAL Logical_Operator_out9772_out1            : std_logic;
  SIGNAL Logical_Operator_out9773_out1            : std_logic;
  SIGNAL Logical_Operator_out9774_out1            : std_logic;
  SIGNAL Logical_Operator_out9775_out1            : std_logic;
  SIGNAL Logical_Operator_out9776_out1            : std_logic;
  SIGNAL Logical_Operator_out9777_out1            : std_logic;
  SIGNAL Logical_Operator_out9778_out1            : std_logic;
  SIGNAL Logical_Operator_out9779_out1            : std_logic;
  SIGNAL Logical_Operator_out9780_out1            : std_logic;
  SIGNAL Logical_Operator_out9781_out1            : std_logic;
  SIGNAL Logical_Operator_out9782_out1            : std_logic;
  SIGNAL Logical_Operator_out9783_out1            : std_logic;
  SIGNAL Logical_Operator_out9784_out1            : std_logic;
  SIGNAL Logical_Operator_out9785_out1            : std_logic;
  SIGNAL Logical_Operator_out9786_out1            : std_logic;
  SIGNAL Logical_Operator_out9787_out1            : std_logic;
  SIGNAL Logical_Operator_out9788_out1            : std_logic;
  SIGNAL Logical_Operator_out9789_out1            : std_logic;
  SIGNAL Logical_Operator_out9790_out1            : std_logic;
  SIGNAL Logical_Operator_out9791_out1            : std_logic;
  SIGNAL Logical_Operator_out9792_out1            : std_logic;
  SIGNAL Logical_Operator_out9793_out1            : std_logic;
  SIGNAL Logical_Operator_out9794_out1            : std_logic;
  SIGNAL Logical_Operator_out9795_out1            : std_logic;
  SIGNAL Logical_Operator_out9796_out1            : std_logic;
  SIGNAL Logical_Operator_out9797_out1            : std_logic;
  SIGNAL Logical_Operator_out9798_out1            : std_logic;
  SIGNAL Logical_Operator_out9799_out1            : std_logic;
  SIGNAL Logical_Operator_out9800_out1            : std_logic;
  SIGNAL Logical_Operator_out9801_out1            : std_logic;
  SIGNAL Logical_Operator_out9802_out1            : std_logic;
  SIGNAL Logical_Operator_out9803_out1            : std_logic;
  SIGNAL Logical_Operator_out9804_out1            : std_logic;
  SIGNAL Logical_Operator_out9805_out1            : std_logic;
  SIGNAL Logical_Operator_out9806_out1            : std_logic;
  SIGNAL Logical_Operator_out9807_out1            : std_logic;
  SIGNAL Logical_Operator_out9808_out1            : std_logic;
  SIGNAL Logical_Operator_out9809_out1            : std_logic;
  SIGNAL Logical_Operator_out9810_out1            : std_logic;
  SIGNAL Logical_Operator_out9811_out1            : std_logic;
  SIGNAL Logical_Operator_out9812_out1            : std_logic;
  SIGNAL Logical_Operator_out9813_out1            : std_logic;
  SIGNAL Logical_Operator_out9814_out1            : std_logic;
  SIGNAL Logical_Operator_out9815_out1            : std_logic;
  SIGNAL Logical_Operator_out9816_out1            : std_logic;
  SIGNAL Logical_Operator_out9817_out1            : std_logic;
  SIGNAL Logical_Operator_out9818_out1            : std_logic;
  SIGNAL Logical_Operator_out9819_out1            : std_logic;
  SIGNAL Logical_Operator_out9820_out1            : std_logic;
  SIGNAL Logical_Operator_out9821_out1            : std_logic;
  SIGNAL Logical_Operator_out9822_out1            : std_logic;
  SIGNAL Logical_Operator_out9823_out1            : std_logic;
  SIGNAL Logical_Operator_out9824_out1            : std_logic;
  SIGNAL Logical_Operator_out9825_out1            : std_logic;
  SIGNAL Logical_Operator_out9826_out1            : std_logic;
  SIGNAL Logical_Operator_out9827_out1            : std_logic;
  SIGNAL Logical_Operator_out9828_out1            : std_logic;
  SIGNAL Logical_Operator_out9829_out1            : std_logic;
  SIGNAL Logical_Operator_out9830_out1            : std_logic;
  SIGNAL Logical_Operator_out9831_out1            : std_logic;
  SIGNAL Logical_Operator_out9832_out1            : std_logic;
  SIGNAL Logical_Operator_out9833_out1            : std_logic;
  SIGNAL Logical_Operator_out9834_out1            : std_logic;
  SIGNAL Logical_Operator_out9835_out1            : std_logic;
  SIGNAL Logical_Operator_out9836_out1            : std_logic;
  SIGNAL Logical_Operator_out9837_out1            : std_logic;
  SIGNAL Logical_Operator_out9838_out1            : std_logic;
  SIGNAL Logical_Operator_out9839_out1            : std_logic;
  SIGNAL Logical_Operator_out9840_out1            : std_logic;
  SIGNAL Logical_Operator_out9841_out1            : std_logic;
  SIGNAL Logical_Operator_out9842_out1            : std_logic;
  SIGNAL Logical_Operator_out9843_out1            : std_logic;
  SIGNAL Logical_Operator_out9844_out1            : std_logic;
  SIGNAL Logical_Operator_out9845_out1            : std_logic;
  SIGNAL Logical_Operator_out9846_out1            : std_logic;
  SIGNAL Logical_Operator_out9847_out1            : std_logic;
  SIGNAL Logical_Operator_out9848_out1            : std_logic;
  SIGNAL Logical_Operator_out9849_out1            : std_logic;
  SIGNAL Logical_Operator_out9850_out1            : std_logic;
  SIGNAL Logical_Operator_out9851_out1            : std_logic;
  SIGNAL Logical_Operator_out9852_out1            : std_logic;
  SIGNAL Logical_Operator_out9853_out1            : std_logic;
  SIGNAL Logical_Operator_out9854_out1            : std_logic;
  SIGNAL Logical_Operator_out9855_out1            : std_logic;
  SIGNAL Logical_Operator_out9856_out1            : std_logic;
  SIGNAL Logical_Operator_out9857_out1            : std_logic;
  SIGNAL Logical_Operator_out9858_out1            : std_logic;
  SIGNAL Logical_Operator_out9859_out1            : std_logic;
  SIGNAL Logical_Operator_out9860_out1            : std_logic;
  SIGNAL Logical_Operator_out9861_out1            : std_logic;
  SIGNAL Logical_Operator_out9862_out1            : std_logic;
  SIGNAL Logical_Operator_out9863_out1            : std_logic;
  SIGNAL Logical_Operator_out9864_out1            : std_logic;
  SIGNAL Logical_Operator_out9865_out1            : std_logic;
  SIGNAL Logical_Operator_out9866_out1            : std_logic;
  SIGNAL Logical_Operator_out9867_out1            : std_logic;
  SIGNAL Logical_Operator_out9868_out1            : std_logic;
  SIGNAL Logical_Operator_out9869_out1            : std_logic;
  SIGNAL Logical_Operator_out9870_out1            : std_logic;
  SIGNAL Logical_Operator_out9871_out1            : std_logic;
  SIGNAL Logical_Operator_out9872_out1            : std_logic;
  SIGNAL Logical_Operator_out9873_out1            : std_logic;
  SIGNAL Logical_Operator_out9874_out1            : std_logic;
  SIGNAL Logical_Operator_out9875_out1            : std_logic;
  SIGNAL Logical_Operator_out9876_out1            : std_logic;
  SIGNAL Logical_Operator_out9877_out1            : std_logic;
  SIGNAL Logical_Operator_out9878_out1            : std_logic;
  SIGNAL Logical_Operator_out9879_out1            : std_logic;
  SIGNAL Logical_Operator_out9880_out1            : std_logic;
  SIGNAL Logical_Operator_out9881_out1            : std_logic;
  SIGNAL Logical_Operator_out9882_out1            : std_logic;
  SIGNAL Logical_Operator_out9883_out1            : std_logic;
  SIGNAL Logical_Operator_out9884_out1            : std_logic;
  SIGNAL Logical_Operator_out9885_out1            : std_logic;
  SIGNAL Logical_Operator_out9886_out1            : std_logic;
  SIGNAL Logical_Operator_out9887_out1            : std_logic;
  SIGNAL Logical_Operator_out9888_out1            : std_logic;
  SIGNAL Logical_Operator_out9889_out1            : std_logic;
  SIGNAL Logical_Operator_out9890_out1            : std_logic;
  SIGNAL Logical_Operator_out9891_out1            : std_logic;
  SIGNAL Logical_Operator_out9892_out1            : std_logic;
  SIGNAL Logical_Operator_out9893_out1            : std_logic;
  SIGNAL Logical_Operator_out9894_out1            : std_logic;
  SIGNAL Logical_Operator_out9895_out1            : std_logic;
  SIGNAL Logical_Operator_out9896_out1            : std_logic;
  SIGNAL Logical_Operator_out9897_out1            : std_logic;
  SIGNAL Logical_Operator_out9898_out1            : std_logic;
  SIGNAL Logical_Operator_out9899_out1            : std_logic;
  SIGNAL Logical_Operator_out9900_out1            : std_logic;
  SIGNAL Logical_Operator_out9901_out1            : std_logic;
  SIGNAL Logical_Operator_out9902_out1            : std_logic;
  SIGNAL Logical_Operator_out9903_out1            : std_logic;
  SIGNAL Logical_Operator_out9904_out1            : std_logic;
  SIGNAL Logical_Operator_out9905_out1            : std_logic;
  SIGNAL Logical_Operator_out9906_out1            : std_logic;
  SIGNAL Logical_Operator_out9907_out1            : std_logic;
  SIGNAL Logical_Operator_out9908_out1            : std_logic;
  SIGNAL Logical_Operator_out9909_out1            : std_logic;
  SIGNAL Logical_Operator_out9910_out1            : std_logic;
  SIGNAL Logical_Operator_out9911_out1            : std_logic;
  SIGNAL Logical_Operator_out9912_out1            : std_logic;
  SIGNAL Logical_Operator_out9913_out1            : std_logic;
  SIGNAL Logical_Operator_out9914_out1            : std_logic;
  SIGNAL Logical_Operator_out9915_out1            : std_logic;
  SIGNAL Logical_Operator_out9916_out1            : std_logic;
  SIGNAL Logical_Operator_out9917_out1            : std_logic;
  SIGNAL Logical_Operator_out9918_out1            : std_logic;
  SIGNAL Logical_Operator_out9919_out1            : std_logic;
  SIGNAL Logical_Operator_out9920_out1            : std_logic;
  SIGNAL Logical_Operator_out9921_out1            : std_logic;
  SIGNAL Logical_Operator_out9922_out1            : std_logic;
  SIGNAL Logical_Operator_out9923_out1            : std_logic;
  SIGNAL Logical_Operator_out9924_out1            : std_logic;
  SIGNAL Logical_Operator_out9925_out1            : std_logic;
  SIGNAL Logical_Operator_out9926_out1            : std_logic;
  SIGNAL Logical_Operator_out9927_out1            : std_logic;
  SIGNAL Logical_Operator_out9928_out1            : std_logic;
  SIGNAL Logical_Operator_out9929_out1            : std_logic;
  SIGNAL Logical_Operator_out9930_out1            : std_logic;
  SIGNAL Logical_Operator_out9931_out1            : std_logic;
  SIGNAL Logical_Operator_out9932_out1            : std_logic;
  SIGNAL Logical_Operator_out9933_out1            : std_logic;
  SIGNAL Logical_Operator_out9934_out1            : std_logic;
  SIGNAL Logical_Operator_out9935_out1            : std_logic;
  SIGNAL Logical_Operator_out9936_out1            : std_logic;
  SIGNAL Logical_Operator_out9937_out1            : std_logic;
  SIGNAL Logical_Operator_out9938_out1            : std_logic;
  SIGNAL Logical_Operator_out9939_out1            : std_logic;
  SIGNAL Logical_Operator_out9940_out1            : std_logic;
  SIGNAL Logical_Operator_out9941_out1            : std_logic;
  SIGNAL Logical_Operator_out9942_out1            : std_logic;
  SIGNAL Logical_Operator_out9943_out1            : std_logic;
  SIGNAL Logical_Operator_out9944_out1            : std_logic;
  SIGNAL Logical_Operator_out9945_out1            : std_logic;
  SIGNAL Logical_Operator_out9946_out1            : std_logic;
  SIGNAL Logical_Operator_out9947_out1            : std_logic;
  SIGNAL Logical_Operator_out9948_out1            : std_logic;
  SIGNAL Logical_Operator_out9949_out1            : std_logic;
  SIGNAL Logical_Operator_out9950_out1            : std_logic;
  SIGNAL Logical_Operator_out9951_out1            : std_logic;
  SIGNAL Logical_Operator_out9952_out1            : std_logic;
  SIGNAL Logical_Operator_out9953_out1            : std_logic;
  SIGNAL Logical_Operator_out9954_out1            : std_logic;
  SIGNAL Logical_Operator_out9955_out1            : std_logic;
  SIGNAL Logical_Operator_out9956_out1            : std_logic;
  SIGNAL Logical_Operator_out9957_out1            : std_logic;
  SIGNAL Logical_Operator_out9958_out1            : std_logic;
  SIGNAL Logical_Operator_out9959_out1            : std_logic;
  SIGNAL Logical_Operator_out9960_out1            : std_logic;
  SIGNAL Logical_Operator_out9961_out1            : std_logic;
  SIGNAL Logical_Operator_out9962_out1            : std_logic;
  SIGNAL Logical_Operator_out9963_out1            : std_logic;
  SIGNAL Logical_Operator_out9964_out1            : std_logic;
  SIGNAL Logical_Operator_out9965_out1            : std_logic;
  SIGNAL Logical_Operator_out9966_out1            : std_logic;
  SIGNAL Logical_Operator_out9967_out1            : std_logic;
  SIGNAL Logical_Operator_out9968_out1            : std_logic;
  SIGNAL Logical_Operator_out9969_out1            : std_logic;
  SIGNAL Logical_Operator_out9970_out1            : std_logic;
  SIGNAL Logical_Operator_out9971_out1            : std_logic;
  SIGNAL Logical_Operator_out9972_out1            : std_logic;
  SIGNAL Logical_Operator_out9973_out1            : std_logic;
  SIGNAL Logical_Operator_out9974_out1            : std_logic;
  SIGNAL Logical_Operator_out9975_out1            : std_logic;
  SIGNAL Logical_Operator_out9976_out1            : std_logic;
  SIGNAL Logical_Operator_out9977_out1            : std_logic;
  SIGNAL Logical_Operator_out9978_out1            : std_logic;
  SIGNAL Logical_Operator_out9979_out1            : std_logic;
  SIGNAL Logical_Operator_out9980_out1            : std_logic;
  SIGNAL Logical_Operator_out9981_out1            : std_logic;
  SIGNAL Logical_Operator_out9982_out1            : std_logic;
  SIGNAL Logical_Operator_out9983_out1            : std_logic;
  SIGNAL Logical_Operator_out9984_out1            : std_logic;
  SIGNAL Logical_Operator_out9985_out1            : std_logic;
  SIGNAL Logical_Operator_out9986_out1            : std_logic;
  SIGNAL Logical_Operator_out9987_out1            : std_logic;
  SIGNAL Logical_Operator_out9988_out1            : std_logic;
  SIGNAL Logical_Operator_out9989_out1            : std_logic;
  SIGNAL Logical_Operator_out9990_out1            : std_logic;
  SIGNAL Logical_Operator_out9991_out1            : std_logic;
  SIGNAL Logical_Operator_out9992_out1            : std_logic;
  SIGNAL Logical_Operator_out9993_out1            : std_logic;
  SIGNAL Logical_Operator_out9994_out1            : std_logic;
  SIGNAL Logical_Operator_out9995_out1            : std_logic;
  SIGNAL Logical_Operator_out9996_out1            : std_logic;
  SIGNAL Logical_Operator_out9997_out1            : std_logic;
  SIGNAL Logical_Operator_out9998_out1            : std_logic;
  SIGNAL Logical_Operator_out9999_out1            : std_logic;
  SIGNAL Logical_Operator_out10000_out1            : std_logic;
  SIGNAL Logical_Operator_out10001_out1            : std_logic;
  SIGNAL Logical_Operator_out10002_out1            : std_logic;
  SIGNAL Logical_Operator_out10003_out1            : std_logic;
  SIGNAL Logical_Operator_out10004_out1            : std_logic;
  SIGNAL Logical_Operator_out10005_out1            : std_logic;
  SIGNAL Logical_Operator_out10006_out1            : std_logic;
  SIGNAL Logical_Operator_out10007_out1            : std_logic;
  SIGNAL Logical_Operator_out10008_out1            : std_logic;
  SIGNAL Logical_Operator_out10009_out1            : std_logic;
  SIGNAL Logical_Operator_out10010_out1            : std_logic;
  SIGNAL Logical_Operator_out10011_out1            : std_logic;
  SIGNAL Logical_Operator_out10012_out1            : std_logic;
  SIGNAL Logical_Operator_out10013_out1            : std_logic;
  SIGNAL Logical_Operator_out10014_out1            : std_logic;
  SIGNAL Logical_Operator_out10015_out1            : std_logic;
  SIGNAL Logical_Operator_out10016_out1            : std_logic;
  SIGNAL Logical_Operator_out10017_out1            : std_logic;
  SIGNAL Logical_Operator_out10018_out1            : std_logic;
  SIGNAL Logical_Operator_out10019_out1            : std_logic;
  SIGNAL Logical_Operator_out10020_out1            : std_logic;
  SIGNAL Logical_Operator_out10021_out1            : std_logic;
  SIGNAL Logical_Operator_out10022_out1            : std_logic;
  SIGNAL Logical_Operator_out10023_out1            : std_logic;
  SIGNAL Logical_Operator_out10024_out1            : std_logic;
  SIGNAL Logical_Operator_out10025_out1            : std_logic;
  SIGNAL Logical_Operator_out10026_out1            : std_logic;
  SIGNAL Logical_Operator_out10027_out1            : std_logic;
  SIGNAL Logical_Operator_out10028_out1            : std_logic;
  SIGNAL Logical_Operator_out10029_out1            : std_logic;
  SIGNAL Logical_Operator_out10030_out1            : std_logic;
  SIGNAL Logical_Operator_out10031_out1            : std_logic;
  SIGNAL Logical_Operator_out10032_out1            : std_logic;
  SIGNAL Logical_Operator_out10033_out1            : std_logic;
  SIGNAL Logical_Operator_out10034_out1            : std_logic;
  SIGNAL Logical_Operator_out10035_out1            : std_logic;
  SIGNAL Logical_Operator_out10036_out1            : std_logic;
  SIGNAL Logical_Operator_out10037_out1            : std_logic;
  SIGNAL Logical_Operator_out10038_out1            : std_logic;
  SIGNAL Logical_Operator_out10039_out1            : std_logic;
  SIGNAL Logical_Operator_out10040_out1            : std_logic;
  SIGNAL Logical_Operator_out10041_out1            : std_logic;
  SIGNAL Logical_Operator_out10042_out1            : std_logic;
  SIGNAL Logical_Operator_out10043_out1            : std_logic;
  SIGNAL Logical_Operator_out10044_out1            : std_logic;
  SIGNAL Logical_Operator_out10045_out1            : std_logic;
  SIGNAL Logical_Operator_out10046_out1            : std_logic;
  SIGNAL Logical_Operator_out10047_out1            : std_logic;
  SIGNAL Logical_Operator_out10048_out1            : std_logic;
  SIGNAL Logical_Operator_out10049_out1            : std_logic;
  SIGNAL Logical_Operator_out10050_out1            : std_logic;
  SIGNAL Logical_Operator_out10051_out1            : std_logic;
  SIGNAL Logical_Operator_out10052_out1            : std_logic;
  SIGNAL Logical_Operator_out10053_out1            : std_logic;
  SIGNAL Logical_Operator_out10054_out1            : std_logic;
  SIGNAL Logical_Operator_out10055_out1            : std_logic;
  SIGNAL Logical_Operator_out10056_out1            : std_logic;
  SIGNAL Logical_Operator_out10057_out1            : std_logic;
  SIGNAL Logical_Operator_out10058_out1            : std_logic;
  SIGNAL Logical_Operator_out10059_out1            : std_logic;
  SIGNAL Logical_Operator_out10060_out1            : std_logic;
  SIGNAL Logical_Operator_out10061_out1            : std_logic;
  SIGNAL Logical_Operator_out10062_out1            : std_logic;
  SIGNAL Logical_Operator_out10063_out1            : std_logic;
  SIGNAL Logical_Operator_out10064_out1            : std_logic;
  SIGNAL Logical_Operator_out10065_out1            : std_logic;
  SIGNAL Logical_Operator_out10066_out1            : std_logic;
  SIGNAL Logical_Operator_out10067_out1            : std_logic;
  SIGNAL Logical_Operator_out10068_out1            : std_logic;
  SIGNAL Logical_Operator_out10069_out1            : std_logic;
  SIGNAL Logical_Operator_out10070_out1            : std_logic;
  SIGNAL Logical_Operator_out10071_out1            : std_logic;
  SIGNAL Logical_Operator_out10072_out1            : std_logic;
  SIGNAL Logical_Operator_out10073_out1            : std_logic;
  SIGNAL Logical_Operator_out10074_out1            : std_logic;
  SIGNAL Logical_Operator_out10075_out1            : std_logic;
  SIGNAL Logical_Operator_out10076_out1            : std_logic;
  SIGNAL Logical_Operator_out10077_out1            : std_logic;
  SIGNAL Logical_Operator_out10078_out1            : std_logic;
  SIGNAL Logical_Operator_out10079_out1            : std_logic;
  SIGNAL Logical_Operator_out10080_out1            : std_logic;
  SIGNAL Logical_Operator_out10081_out1            : std_logic;
  SIGNAL Logical_Operator_out10082_out1            : std_logic;
  SIGNAL Logical_Operator_out10083_out1            : std_logic;
  SIGNAL Logical_Operator_out10084_out1            : std_logic;
  SIGNAL Logical_Operator_out10085_out1            : std_logic;
  SIGNAL Logical_Operator_out10086_out1            : std_logic;
  SIGNAL Logical_Operator_out10087_out1            : std_logic;
  SIGNAL Logical_Operator_out10088_out1            : std_logic;
  SIGNAL Logical_Operator_out10089_out1            : std_logic;
  SIGNAL Logical_Operator_out10090_out1            : std_logic;
  SIGNAL Logical_Operator_out10091_out1            : std_logic;
  SIGNAL Logical_Operator_out10092_out1            : std_logic;
  SIGNAL Logical_Operator_out10093_out1            : std_logic;
  SIGNAL Logical_Operator_out10094_out1            : std_logic;
  SIGNAL Logical_Operator_out10095_out1            : std_logic;
  SIGNAL Logical_Operator_out10096_out1            : std_logic;
  SIGNAL Logical_Operator_out10097_out1            : std_logic;
  SIGNAL Logical_Operator_out10098_out1            : std_logic;
  SIGNAL Logical_Operator_out10099_out1            : std_logic;
  SIGNAL Logical_Operator_out10100_out1            : std_logic;
  SIGNAL Logical_Operator_out10101_out1            : std_logic;
  SIGNAL Logical_Operator_out10102_out1            : std_logic;
  SIGNAL Logical_Operator_out10103_out1            : std_logic;
  SIGNAL Logical_Operator_out10104_out1            : std_logic;
  SIGNAL Logical_Operator_out10105_out1            : std_logic;
  SIGNAL Logical_Operator_out10106_out1            : std_logic;
  SIGNAL Logical_Operator_out10107_out1            : std_logic;
  SIGNAL Logical_Operator_out10108_out1            : std_logic;
  SIGNAL Logical_Operator_out10109_out1            : std_logic;
  SIGNAL Logical_Operator_out10110_out1            : std_logic;
  SIGNAL Logical_Operator_out10111_out1            : std_logic;
  SIGNAL Logical_Operator_out10112_out1            : std_logic;
  SIGNAL Logical_Operator_out10113_out1            : std_logic;
  SIGNAL Logical_Operator_out10114_out1            : std_logic;
  SIGNAL Logical_Operator_out10115_out1            : std_logic;
  SIGNAL Logical_Operator_out10116_out1            : std_logic;
  SIGNAL Logical_Operator_out10117_out1            : std_logic;
  SIGNAL Logical_Operator_out10118_out1            : std_logic;
  SIGNAL Logical_Operator_out10119_out1            : std_logic;
  SIGNAL Logical_Operator_out10120_out1            : std_logic;
  SIGNAL Logical_Operator_out10121_out1            : std_logic;
  SIGNAL Logical_Operator_out10122_out1            : std_logic;
  SIGNAL Logical_Operator_out10123_out1            : std_logic;
  SIGNAL Logical_Operator_out10124_out1            : std_logic;
  SIGNAL Logical_Operator_out10125_out1            : std_logic;
  SIGNAL Logical_Operator_out10126_out1            : std_logic;
  SIGNAL Logical_Operator_out10127_out1            : std_logic;
  SIGNAL Logical_Operator_out10128_out1            : std_logic;
  SIGNAL Logical_Operator_out10129_out1            : std_logic;
  SIGNAL Logical_Operator_out10130_out1            : std_logic;
  SIGNAL Logical_Operator_out10131_out1            : std_logic;
  SIGNAL Logical_Operator_out10132_out1            : std_logic;
  SIGNAL Logical_Operator_out10133_out1            : std_logic;
  SIGNAL Logical_Operator_out10134_out1            : std_logic;
  SIGNAL Logical_Operator_out10135_out1            : std_logic;
  SIGNAL Logical_Operator_out10136_out1            : std_logic;
  SIGNAL Logical_Operator_out10137_out1            : std_logic;
  SIGNAL Logical_Operator_out10138_out1            : std_logic;
  SIGNAL Logical_Operator_out10139_out1            : std_logic;
  SIGNAL Logical_Operator_out10140_out1            : std_logic;
  SIGNAL Logical_Operator_out10141_out1            : std_logic;
  SIGNAL Logical_Operator_out10142_out1            : std_logic;
  SIGNAL Logical_Operator_out10143_out1            : std_logic;
  SIGNAL Logical_Operator_out10144_out1            : std_logic;
  SIGNAL Logical_Operator_out10145_out1            : std_logic;
  SIGNAL Logical_Operator_out10146_out1            : std_logic;
  SIGNAL Logical_Operator_out10147_out1            : std_logic;
  SIGNAL Logical_Operator_out10148_out1            : std_logic;
  SIGNAL Logical_Operator_out10149_out1            : std_logic;
  SIGNAL Logical_Operator_out10150_out1            : std_logic;
  SIGNAL Logical_Operator_out10151_out1            : std_logic;
  SIGNAL Logical_Operator_out10152_out1            : std_logic;
  SIGNAL Logical_Operator_out10153_out1            : std_logic;
  SIGNAL Logical_Operator_out10154_out1            : std_logic;
  SIGNAL Logical_Operator_out10155_out1            : std_logic;
  SIGNAL Logical_Operator_out10156_out1            : std_logic;
  SIGNAL Logical_Operator_out10157_out1            : std_logic;
  SIGNAL Logical_Operator_out10158_out1            : std_logic;
  SIGNAL Logical_Operator_out10159_out1            : std_logic;
  SIGNAL Logical_Operator_out10160_out1            : std_logic;
  SIGNAL Logical_Operator_out10161_out1            : std_logic;
  SIGNAL Logical_Operator_out10162_out1            : std_logic;
  SIGNAL Logical_Operator_out10163_out1            : std_logic;
  SIGNAL Logical_Operator_out10164_out1            : std_logic;
  SIGNAL Logical_Operator_out10165_out1            : std_logic;
  SIGNAL Logical_Operator_out10166_out1            : std_logic;
  SIGNAL Logical_Operator_out10167_out1            : std_logic;
  SIGNAL Logical_Operator_out10168_out1            : std_logic;
  SIGNAL Logical_Operator_out10169_out1            : std_logic;
  SIGNAL Logical_Operator_out10170_out1            : std_logic;
  SIGNAL Logical_Operator_out10171_out1            : std_logic;
  SIGNAL Logical_Operator_out10172_out1            : std_logic;
  SIGNAL Logical_Operator_out10173_out1            : std_logic;
  SIGNAL Logical_Operator_out10174_out1            : std_logic;
  SIGNAL Logical_Operator_out10175_out1            : std_logic;
  SIGNAL Logical_Operator_out10176_out1            : std_logic;
  SIGNAL Logical_Operator_out10177_out1            : std_logic;
  SIGNAL Logical_Operator_out10178_out1            : std_logic;
  SIGNAL Logical_Operator_out10179_out1            : std_logic;
  SIGNAL Logical_Operator_out10180_out1            : std_logic;
  SIGNAL Logical_Operator_out10181_out1            : std_logic;
  SIGNAL Logical_Operator_out10182_out1            : std_logic;
  SIGNAL Logical_Operator_out10183_out1            : std_logic;
  SIGNAL Logical_Operator_out10184_out1            : std_logic;
  SIGNAL Logical_Operator_out10185_out1            : std_logic;
  SIGNAL Logical_Operator_out10186_out1            : std_logic;
  SIGNAL Logical_Operator_out10187_out1            : std_logic;
  SIGNAL Logical_Operator_out10188_out1            : std_logic;
  SIGNAL Logical_Operator_out10189_out1            : std_logic;
  SIGNAL Logical_Operator_out10190_out1            : std_logic;
  SIGNAL Logical_Operator_out10191_out1            : std_logic;
  SIGNAL Logical_Operator_out10192_out1            : std_logic;
  SIGNAL Logical_Operator_out10193_out1            : std_logic;
  SIGNAL Logical_Operator_out10194_out1            : std_logic;
  SIGNAL Logical_Operator_out10195_out1            : std_logic;
  SIGNAL Logical_Operator_out10196_out1            : std_logic;
  SIGNAL Logical_Operator_out10197_out1            : std_logic;
  SIGNAL Logical_Operator_out10198_out1            : std_logic;
  SIGNAL Logical_Operator_out10199_out1            : std_logic;
  SIGNAL Logical_Operator_out10200_out1            : std_logic;
  SIGNAL Logical_Operator_out10201_out1            : std_logic;
  SIGNAL Logical_Operator_out10202_out1            : std_logic;
  SIGNAL Logical_Operator_out10203_out1            : std_logic;
  SIGNAL Logical_Operator_out10204_out1            : std_logic;
  SIGNAL Logical_Operator_out10205_out1            : std_logic;
  SIGNAL Logical_Operator_out10206_out1            : std_logic;
  SIGNAL Logical_Operator_out10207_out1            : std_logic;
  SIGNAL Logical_Operator_out10208_out1            : std_logic;
  SIGNAL Logical_Operator_out10209_out1            : std_logic;
  SIGNAL Logical_Operator_out10210_out1            : std_logic;
  SIGNAL Logical_Operator_out10211_out1            : std_logic;
  SIGNAL Logical_Operator_out10212_out1            : std_logic;
  SIGNAL Logical_Operator_out10213_out1            : std_logic;
  SIGNAL Logical_Operator_out10214_out1            : std_logic;
  SIGNAL Logical_Operator_out10215_out1            : std_logic;
  SIGNAL Logical_Operator_out10216_out1            : std_logic;
  SIGNAL Logical_Operator_out10217_out1            : std_logic;
  SIGNAL Logical_Operator_out10218_out1            : std_logic;
  SIGNAL Logical_Operator_out10219_out1            : std_logic;
  SIGNAL Logical_Operator_out10220_out1            : std_logic;
  SIGNAL Logical_Operator_out10221_out1            : std_logic;
  SIGNAL Logical_Operator_out10222_out1            : std_logic;
  SIGNAL Logical_Operator_out10223_out1            : std_logic;
  SIGNAL Logical_Operator_out10224_out1            : std_logic;
  SIGNAL Logical_Operator_out10225_out1            : std_logic;
  SIGNAL Logical_Operator_out10226_out1            : std_logic;
  SIGNAL Logical_Operator_out10227_out1            : std_logic;
  SIGNAL Logical_Operator_out10228_out1            : std_logic;
  SIGNAL Logical_Operator_out10229_out1            : std_logic;
  SIGNAL Logical_Operator_out10230_out1            : std_logic;
  SIGNAL Logical_Operator_out10231_out1            : std_logic;
  SIGNAL Logical_Operator_out10232_out1            : std_logic;
  SIGNAL Logical_Operator_out10233_out1            : std_logic;
  SIGNAL Logical_Operator_out10234_out1            : std_logic;
  SIGNAL Logical_Operator_out10235_out1            : std_logic;
  SIGNAL Logical_Operator_out10236_out1            : std_logic;
  SIGNAL Logical_Operator_out10237_out1            : std_logic;
  SIGNAL Logical_Operator_out10238_out1            : std_logic;
  SIGNAL Logical_Operator_out10239_out1            : std_logic;
  SIGNAL Logical_Operator_out10240_out1            : std_logic;
  SIGNAL Logical_Operator_out10241_out1            : std_logic;
  SIGNAL Logical_Operator_out10242_out1            : std_logic;
  SIGNAL Logical_Operator_out10243_out1            : std_logic;
  SIGNAL Logical_Operator_out10244_out1            : std_logic;
  SIGNAL Logical_Operator_out10245_out1            : std_logic;
  SIGNAL Logical_Operator_out10246_out1            : std_logic;
  SIGNAL Logical_Operator_out10247_out1            : std_logic;
  SIGNAL Logical_Operator_out10248_out1            : std_logic;
  SIGNAL Logical_Operator_out10249_out1            : std_logic;
  SIGNAL Logical_Operator_out10250_out1            : std_logic;
  SIGNAL Logical_Operator_out10251_out1            : std_logic;
  SIGNAL Logical_Operator_out10252_out1            : std_logic;
  SIGNAL Logical_Operator_out10253_out1            : std_logic;
  SIGNAL Logical_Operator_out10254_out1            : std_logic;
  SIGNAL Logical_Operator_out10255_out1            : std_logic;
  SIGNAL Logical_Operator_out10256_out1            : std_logic;
  SIGNAL Logical_Operator_out10257_out1            : std_logic;
  SIGNAL Logical_Operator_out10258_out1            : std_logic;
  SIGNAL Logical_Operator_out10259_out1            : std_logic;
  SIGNAL Logical_Operator_out10260_out1            : std_logic;
  SIGNAL Logical_Operator_out10261_out1            : std_logic;
  SIGNAL Logical_Operator_out10262_out1            : std_logic;
  SIGNAL Logical_Operator_out10263_out1            : std_logic;
  SIGNAL Logical_Operator_out10264_out1            : std_logic;
  SIGNAL Logical_Operator_out10265_out1            : std_logic;
  SIGNAL Logical_Operator_out10266_out1            : std_logic;
  SIGNAL Logical_Operator_out10267_out1            : std_logic;
  SIGNAL Logical_Operator_out10268_out1            : std_logic;
  SIGNAL Logical_Operator_out10269_out1            : std_logic;
  SIGNAL Logical_Operator_out10270_out1            : std_logic;
  SIGNAL Logical_Operator_out10271_out1            : std_logic;
  SIGNAL Logical_Operator_out10272_out1            : std_logic;
  SIGNAL Logical_Operator_out10273_out1            : std_logic;
  SIGNAL Logical_Operator_out10274_out1            : std_logic;
  SIGNAL Logical_Operator_out10275_out1            : std_logic;
  SIGNAL Logical_Operator_out10276_out1            : std_logic;
  SIGNAL Logical_Operator_out10277_out1            : std_logic;
  SIGNAL Logical_Operator_out10278_out1            : std_logic;
  SIGNAL Logical_Operator_out10279_out1            : std_logic;
  SIGNAL Logical_Operator_out10280_out1            : std_logic;
  SIGNAL Logical_Operator_out10281_out1            : std_logic;
  SIGNAL Logical_Operator_out10282_out1            : std_logic;
  SIGNAL Logical_Operator_out10283_out1            : std_logic;
  SIGNAL Logical_Operator_out10284_out1            : std_logic;
  SIGNAL Logical_Operator_out10285_out1            : std_logic;
  SIGNAL Logical_Operator_out10286_out1            : std_logic;
  SIGNAL Logical_Operator_out10287_out1            : std_logic;
  SIGNAL Logical_Operator_out10288_out1            : std_logic;
  SIGNAL Logical_Operator_out10289_out1            : std_logic;
  SIGNAL Logical_Operator_out10290_out1            : std_logic;
  SIGNAL Logical_Operator_out10291_out1            : std_logic;
  SIGNAL Logical_Operator_out10292_out1            : std_logic;
  SIGNAL Logical_Operator_out10293_out1            : std_logic;
  SIGNAL Logical_Operator_out10294_out1            : std_logic;
  SIGNAL Logical_Operator_out10295_out1            : std_logic;
  SIGNAL Logical_Operator_out10296_out1            : std_logic;
  SIGNAL Logical_Operator_out10297_out1            : std_logic;
  SIGNAL Logical_Operator_out10298_out1            : std_logic;
  SIGNAL Logical_Operator_out10299_out1            : std_logic;
  SIGNAL Logical_Operator_out10300_out1            : std_logic;
  SIGNAL Logical_Operator_out10301_out1            : std_logic;
  SIGNAL Logical_Operator_out10302_out1            : std_logic;
  SIGNAL Logical_Operator_out10303_out1            : std_logic;
  SIGNAL Logical_Operator_out10304_out1            : std_logic;
  SIGNAL Logical_Operator_out10305_out1            : std_logic;
  SIGNAL Logical_Operator_out10306_out1            : std_logic;
  SIGNAL Logical_Operator_out10307_out1            : std_logic;
  SIGNAL Logical_Operator_out10308_out1            : std_logic;
  SIGNAL Logical_Operator_out10309_out1            : std_logic;
  SIGNAL Logical_Operator_out10310_out1            : std_logic;
  SIGNAL Logical_Operator_out10311_out1            : std_logic;
  SIGNAL Logical_Operator_out10312_out1            : std_logic;
  SIGNAL Logical_Operator_out10313_out1            : std_logic;
  SIGNAL Logical_Operator_out10314_out1            : std_logic;
  SIGNAL Logical_Operator_out10315_out1            : std_logic;
  SIGNAL Logical_Operator_out10316_out1            : std_logic;
  SIGNAL Logical_Operator_out10317_out1            : std_logic;
  SIGNAL Logical_Operator_out10318_out1            : std_logic;
  SIGNAL Logical_Operator_out10319_out1            : std_logic;
  SIGNAL Logical_Operator_out10320_out1            : std_logic;
  SIGNAL Logical_Operator_out10321_out1            : std_logic;
  SIGNAL Logical_Operator_out10322_out1            : std_logic;
  SIGNAL Logical_Operator_out10323_out1            : std_logic;
  SIGNAL Logical_Operator_out10324_out1            : std_logic;
  SIGNAL Logical_Operator_out10325_out1            : std_logic;
  SIGNAL Logical_Operator_out10326_out1            : std_logic;
  SIGNAL Logical_Operator_out10327_out1            : std_logic;
  SIGNAL Logical_Operator_out10328_out1            : std_logic;
  SIGNAL Logical_Operator_out10329_out1            : std_logic;
  SIGNAL Logical_Operator_out10330_out1            : std_logic;
  SIGNAL Logical_Operator_out10331_out1            : std_logic;
  SIGNAL Logical_Operator_out10332_out1            : std_logic;
  SIGNAL Logical_Operator_out10333_out1            : std_logic;
  SIGNAL Logical_Operator_out10334_out1            : std_logic;
  SIGNAL Logical_Operator_out10335_out1            : std_logic;
  SIGNAL Logical_Operator_out10336_out1            : std_logic;
  SIGNAL Logical_Operator_out10337_out1            : std_logic;
  SIGNAL Logical_Operator_out10338_out1            : std_logic;
  SIGNAL Logical_Operator_out10339_out1            : std_logic;
  SIGNAL Logical_Operator_out10340_out1            : std_logic;
  SIGNAL Logical_Operator_out10341_out1            : std_logic;
  SIGNAL Logical_Operator_out10342_out1            : std_logic;
  SIGNAL Logical_Operator_out10343_out1            : std_logic;
  SIGNAL Logical_Operator_out10344_out1            : std_logic;
  SIGNAL Logical_Operator_out10345_out1            : std_logic;
  SIGNAL Logical_Operator_out10346_out1            : std_logic;
  SIGNAL Logical_Operator_out10347_out1            : std_logic;
  SIGNAL Logical_Operator_out10348_out1            : std_logic;
  SIGNAL Logical_Operator_out10349_out1            : std_logic;
  SIGNAL Logical_Operator_out10350_out1            : std_logic;
  SIGNAL Logical_Operator_out10351_out1            : std_logic;
  SIGNAL Logical_Operator_out10352_out1            : std_logic;
  SIGNAL Logical_Operator_out10353_out1            : std_logic;
  SIGNAL Logical_Operator_out10354_out1            : std_logic;
  SIGNAL Logical_Operator_out10355_out1            : std_logic;
  SIGNAL Logical_Operator_out10356_out1            : std_logic;
  SIGNAL Logical_Operator_out10357_out1            : std_logic;
  SIGNAL Logical_Operator_out10358_out1            : std_logic;
  SIGNAL Logical_Operator_out10359_out1            : std_logic;
  SIGNAL Logical_Operator_out10360_out1            : std_logic;
  SIGNAL Logical_Operator_out10361_out1            : std_logic;
  SIGNAL Logical_Operator_out10362_out1            : std_logic;
  SIGNAL Logical_Operator_out10363_out1            : std_logic;
  SIGNAL Logical_Operator_out10364_out1            : std_logic;
  SIGNAL Logical_Operator_out10365_out1            : std_logic;
  SIGNAL Logical_Operator_out10366_out1            : std_logic;
  SIGNAL Logical_Operator_out10367_out1            : std_logic;
  SIGNAL Logical_Operator_out10368_out1            : std_logic;
  SIGNAL Logical_Operator_out10369_out1            : std_logic;
  SIGNAL Logical_Operator_out10370_out1            : std_logic;
  SIGNAL Logical_Operator_out10371_out1            : std_logic;
  SIGNAL Logical_Operator_out10372_out1            : std_logic;
  SIGNAL Logical_Operator_out10373_out1            : std_logic;
  SIGNAL Logical_Operator_out10374_out1            : std_logic;
  SIGNAL Logical_Operator_out10375_out1            : std_logic;
  SIGNAL Logical_Operator_out10376_out1            : std_logic;
  SIGNAL Logical_Operator_out10377_out1            : std_logic;
  SIGNAL Logical_Operator_out10378_out1            : std_logic;
  SIGNAL Logical_Operator_out10379_out1            : std_logic;
  SIGNAL Logical_Operator_out10380_out1            : std_logic;
  SIGNAL Logical_Operator_out10381_out1            : std_logic;
  SIGNAL Logical_Operator_out10382_out1            : std_logic;
  SIGNAL Logical_Operator_out10383_out1            : std_logic;
  SIGNAL Logical_Operator_out10384_out1            : std_logic;
  SIGNAL Logical_Operator_out10385_out1            : std_logic;
  SIGNAL Logical_Operator_out10386_out1            : std_logic;
  SIGNAL Logical_Operator_out10387_out1            : std_logic;
  SIGNAL Logical_Operator_out10388_out1            : std_logic;
  SIGNAL Logical_Operator_out10389_out1            : std_logic;
  SIGNAL Logical_Operator_out10390_out1            : std_logic;
  SIGNAL Logical_Operator_out10391_out1            : std_logic;
  SIGNAL Logical_Operator_out10392_out1            : std_logic;
  SIGNAL Logical_Operator_out10393_out1            : std_logic;
  SIGNAL Logical_Operator_out10394_out1            : std_logic;
  SIGNAL Logical_Operator_out10395_out1            : std_logic;
  SIGNAL Logical_Operator_out10396_out1            : std_logic;
  SIGNAL Logical_Operator_out10397_out1            : std_logic;
  SIGNAL Logical_Operator_out10398_out1            : std_logic;
  SIGNAL Logical_Operator_out10399_out1            : std_logic;
  SIGNAL Logical_Operator_out10400_out1            : std_logic;
  SIGNAL Logical_Operator_out10401_out1            : std_logic;
  SIGNAL Logical_Operator_out10402_out1            : std_logic;
  SIGNAL Logical_Operator_out10403_out1            : std_logic;
  SIGNAL Logical_Operator_out10404_out1            : std_logic;
  SIGNAL Logical_Operator_out10405_out1            : std_logic;
  SIGNAL Logical_Operator_out10406_out1            : std_logic;
  SIGNAL Logical_Operator_out10407_out1            : std_logic;
  SIGNAL Logical_Operator_out10408_out1            : std_logic;
  SIGNAL Logical_Operator_out10409_out1            : std_logic;
  SIGNAL Logical_Operator_out10410_out1            : std_logic;
  SIGNAL Logical_Operator_out10411_out1            : std_logic;
  SIGNAL Logical_Operator_out10412_out1            : std_logic;
  SIGNAL Logical_Operator_out10413_out1            : std_logic;
  SIGNAL Logical_Operator_out10414_out1            : std_logic;
  SIGNAL Logical_Operator_out10415_out1            : std_logic;
  SIGNAL Logical_Operator_out10416_out1            : std_logic;
  SIGNAL Logical_Operator_out10417_out1            : std_logic;
  SIGNAL Logical_Operator_out10418_out1            : std_logic;
  SIGNAL Logical_Operator_out10419_out1            : std_logic;
  SIGNAL Logical_Operator_out10420_out1            : std_logic;
  SIGNAL Logical_Operator_out10421_out1            : std_logic;
  SIGNAL Logical_Operator_out10422_out1            : std_logic;
  SIGNAL Logical_Operator_out10423_out1            : std_logic;
  SIGNAL Logical_Operator_out10424_out1            : std_logic;
  SIGNAL Logical_Operator_out10425_out1            : std_logic;
  SIGNAL Logical_Operator_out10426_out1            : std_logic;
  SIGNAL Logical_Operator_out10427_out1            : std_logic;
  SIGNAL Logical_Operator_out10428_out1            : std_logic;
  SIGNAL Logical_Operator_out10429_out1            : std_logic;
  SIGNAL Logical_Operator_out10430_out1            : std_logic;
  SIGNAL Logical_Operator_out10431_out1            : std_logic;
  SIGNAL Logical_Operator_out10432_out1            : std_logic;
  SIGNAL Logical_Operator_out10433_out1            : std_logic;
  SIGNAL Logical_Operator_out10434_out1            : std_logic;
  SIGNAL Logical_Operator_out10435_out1            : std_logic;
  SIGNAL Logical_Operator_out10436_out1            : std_logic;
  SIGNAL Logical_Operator_out10437_out1            : std_logic;
  SIGNAL Logical_Operator_out10438_out1            : std_logic;
  SIGNAL Logical_Operator_out10439_out1            : std_logic;
  SIGNAL Logical_Operator_out10440_out1            : std_logic;
  SIGNAL Logical_Operator_out10441_out1            : std_logic;
  SIGNAL Logical_Operator_out10442_out1            : std_logic;
  SIGNAL Logical_Operator_out10443_out1            : std_logic;
  SIGNAL Logical_Operator_out10444_out1            : std_logic;
  SIGNAL Logical_Operator_out10445_out1            : std_logic;
  SIGNAL Logical_Operator_out10446_out1            : std_logic;
  SIGNAL Logical_Operator_out10447_out1            : std_logic;
  SIGNAL Logical_Operator_out10448_out1            : std_logic;
  SIGNAL Logical_Operator_out10449_out1            : std_logic;
  SIGNAL Logical_Operator_out10450_out1            : std_logic;
  SIGNAL Logical_Operator_out10451_out1            : std_logic;
  SIGNAL Logical_Operator_out10452_out1            : std_logic;
  SIGNAL Logical_Operator_out10453_out1            : std_logic;
  SIGNAL Logical_Operator_out10454_out1            : std_logic;
  SIGNAL Logical_Operator_out10455_out1            : std_logic;
  SIGNAL Logical_Operator_out10456_out1            : std_logic;
  SIGNAL Logical_Operator_out10457_out1            : std_logic;
  SIGNAL Logical_Operator_out10458_out1            : std_logic;
  SIGNAL Logical_Operator_out10459_out1            : std_logic;
  SIGNAL Logical_Operator_out10460_out1            : std_logic;
  SIGNAL Logical_Operator_out10461_out1            : std_logic;
  SIGNAL Logical_Operator_out10462_out1            : std_logic;
  SIGNAL Logical_Operator_out10463_out1            : std_logic;
  SIGNAL Logical_Operator_out10464_out1            : std_logic;
  SIGNAL Logical_Operator_out10465_out1            : std_logic;
  SIGNAL Logical_Operator_out10466_out1            : std_logic;
  SIGNAL Logical_Operator_out10467_out1            : std_logic;
  SIGNAL Logical_Operator_out10468_out1            : std_logic;
  SIGNAL Logical_Operator_out10469_out1            : std_logic;
  SIGNAL Logical_Operator_out10470_out1            : std_logic;
  SIGNAL Logical_Operator_out10471_out1            : std_logic;
  SIGNAL Logical_Operator_out10472_out1            : std_logic;
  SIGNAL Logical_Operator_out10473_out1            : std_logic;
  SIGNAL Logical_Operator_out10474_out1            : std_logic;
  SIGNAL Logical_Operator_out10475_out1            : std_logic;
  SIGNAL Logical_Operator_out10476_out1            : std_logic;
  SIGNAL Logical_Operator_out10477_out1            : std_logic;
  SIGNAL Logical_Operator_out10478_out1            : std_logic;
  SIGNAL Logical_Operator_out10479_out1            : std_logic;
  SIGNAL Logical_Operator_out10480_out1            : std_logic;
  SIGNAL Logical_Operator_out10481_out1            : std_logic;
  SIGNAL Logical_Operator_out10482_out1            : std_logic;
  SIGNAL Logical_Operator_out10483_out1            : std_logic;
  SIGNAL Logical_Operator_out10484_out1            : std_logic;
  SIGNAL Logical_Operator_out10485_out1            : std_logic;
  SIGNAL Logical_Operator_out10486_out1            : std_logic;
  SIGNAL Logical_Operator_out10487_out1            : std_logic;
  SIGNAL Logical_Operator_out10488_out1            : std_logic;
  SIGNAL Logical_Operator_out10489_out1            : std_logic;
  SIGNAL Logical_Operator_out10490_out1            : std_logic;
  SIGNAL Logical_Operator_out10491_out1            : std_logic;
  SIGNAL Logical_Operator_out10492_out1            : std_logic;
  SIGNAL Logical_Operator_out10493_out1            : std_logic;
  SIGNAL Logical_Operator_out10494_out1            : std_logic;
  SIGNAL Logical_Operator_out10495_out1            : std_logic;
  SIGNAL Logical_Operator_out10496_out1            : std_logic;
  SIGNAL Logical_Operator_out10497_out1            : std_logic;
  SIGNAL Logical_Operator_out10498_out1            : std_logic;
  SIGNAL Logical_Operator_out10499_out1            : std_logic;
  SIGNAL Logical_Operator_out10500_out1            : std_logic;
  SIGNAL Logical_Operator_out10501_out1            : std_logic;
  SIGNAL Logical_Operator_out10502_out1            : std_logic;
  SIGNAL Logical_Operator_out10503_out1            : std_logic;
  SIGNAL Logical_Operator_out10504_out1            : std_logic;
  SIGNAL Logical_Operator_out10505_out1            : std_logic;
  SIGNAL Logical_Operator_out10506_out1            : std_logic;
  SIGNAL Logical_Operator_out10507_out1            : std_logic;
  SIGNAL Logical_Operator_out10508_out1            : std_logic;
  SIGNAL Logical_Operator_out10509_out1            : std_logic;
  SIGNAL Logical_Operator_out10510_out1            : std_logic;
  SIGNAL Logical_Operator_out10511_out1            : std_logic;
  SIGNAL Logical_Operator_out10512_out1            : std_logic;
  SIGNAL Logical_Operator_out10513_out1            : std_logic;
  SIGNAL Logical_Operator_out10514_out1            : std_logic;
  SIGNAL Logical_Operator_out10515_out1            : std_logic;
  SIGNAL Logical_Operator_out10516_out1            : std_logic;
  SIGNAL Logical_Operator_out10517_out1            : std_logic;
  SIGNAL Logical_Operator_out10518_out1            : std_logic;
  SIGNAL Logical_Operator_out10519_out1            : std_logic;
  SIGNAL Logical_Operator_out10520_out1            : std_logic;
  SIGNAL Logical_Operator_out10521_out1            : std_logic;
  SIGNAL Logical_Operator_out10522_out1            : std_logic;
  SIGNAL Logical_Operator_out10523_out1            : std_logic;
  SIGNAL Logical_Operator_out10524_out1            : std_logic;
  SIGNAL Logical_Operator_out10525_out1            : std_logic;
  SIGNAL Logical_Operator_out10526_out1            : std_logic;
  SIGNAL Logical_Operator_out10527_out1            : std_logic;
  SIGNAL Logical_Operator_out10528_out1            : std_logic;
  SIGNAL Logical_Operator_out10529_out1            : std_logic;
  SIGNAL Logical_Operator_out10530_out1            : std_logic;
  SIGNAL Logical_Operator_out10531_out1            : std_logic;
  SIGNAL Logical_Operator_out10532_out1            : std_logic;
  SIGNAL Logical_Operator_out10533_out1            : std_logic;
  SIGNAL Logical_Operator_out10534_out1            : std_logic;
  SIGNAL Logical_Operator_out10535_out1            : std_logic;
  SIGNAL Logical_Operator_out10536_out1            : std_logic;
  SIGNAL Logical_Operator_out10537_out1            : std_logic;
  SIGNAL Logical_Operator_out10538_out1            : std_logic;
  SIGNAL Logical_Operator_out10539_out1            : std_logic;
  SIGNAL Logical_Operator_out10540_out1            : std_logic;
  SIGNAL Logical_Operator_out10541_out1            : std_logic;
  SIGNAL Logical_Operator_out10542_out1            : std_logic;
  SIGNAL Logical_Operator_out10543_out1            : std_logic;
  SIGNAL Logical_Operator_out10544_out1            : std_logic;
  SIGNAL Logical_Operator_out10545_out1            : std_logic;
  SIGNAL Logical_Operator_out10546_out1            : std_logic;
  SIGNAL Logical_Operator_out10547_out1            : std_logic;
  SIGNAL Logical_Operator_out10548_out1            : std_logic;
  SIGNAL Logical_Operator_out10549_out1            : std_logic;
  SIGNAL Logical_Operator_out10550_out1            : std_logic;
  SIGNAL Logical_Operator_out10551_out1            : std_logic;
  SIGNAL Logical_Operator_out10552_out1            : std_logic;
  SIGNAL Logical_Operator_out10553_out1            : std_logic;
  SIGNAL Logical_Operator_out10554_out1            : std_logic;
  SIGNAL Logical_Operator_out10555_out1            : std_logic;
  SIGNAL Logical_Operator_out10556_out1            : std_logic;
  SIGNAL Logical_Operator_out10557_out1            : std_logic;
  SIGNAL Logical_Operator_out10558_out1            : std_logic;
  SIGNAL Logical_Operator_out10559_out1            : std_logic;
  SIGNAL Logical_Operator_out10560_out1            : std_logic;
  SIGNAL Logical_Operator_out10561_out1            : std_logic;
  SIGNAL Logical_Operator_out10562_out1            : std_logic;
  SIGNAL Logical_Operator_out10563_out1            : std_logic;
  SIGNAL Logical_Operator_out10564_out1            : std_logic;
  SIGNAL Logical_Operator_out10565_out1            : std_logic;
  SIGNAL Logical_Operator_out10566_out1            : std_logic;
  SIGNAL Logical_Operator_out10567_out1            : std_logic;
  SIGNAL Logical_Operator_out10568_out1            : std_logic;
  SIGNAL Logical_Operator_out10569_out1            : std_logic;
  SIGNAL Logical_Operator_out10570_out1            : std_logic;
  SIGNAL Logical_Operator_out10571_out1            : std_logic;
  SIGNAL Logical_Operator_out10572_out1            : std_logic;
  SIGNAL Logical_Operator_out10573_out1            : std_logic;
  SIGNAL Logical_Operator_out10574_out1            : std_logic;
  SIGNAL Logical_Operator_out10575_out1            : std_logic;
  SIGNAL Logical_Operator_out10576_out1            : std_logic;
  SIGNAL Logical_Operator_out10577_out1            : std_logic;
  SIGNAL Logical_Operator_out10578_out1            : std_logic;
  SIGNAL Logical_Operator_out10579_out1            : std_logic;
  SIGNAL Logical_Operator_out10580_out1            : std_logic;
  SIGNAL Logical_Operator_out10581_out1            : std_logic;
  SIGNAL Logical_Operator_out10582_out1            : std_logic;
  SIGNAL Logical_Operator_out10583_out1            : std_logic;
  SIGNAL Logical_Operator_out10584_out1            : std_logic;
  SIGNAL Logical_Operator_out10585_out1            : std_logic;
  SIGNAL Logical_Operator_out10586_out1            : std_logic;
  SIGNAL Logical_Operator_out10587_out1            : std_logic;
  SIGNAL Logical_Operator_out10588_out1            : std_logic;
  SIGNAL Logical_Operator_out10589_out1            : std_logic;
  SIGNAL Logical_Operator_out10590_out1            : std_logic;
  SIGNAL Logical_Operator_out10591_out1            : std_logic;
  SIGNAL Logical_Operator_out10592_out1            : std_logic;
  SIGNAL Logical_Operator_out10593_out1            : std_logic;
  SIGNAL Logical_Operator_out10594_out1            : std_logic;
  SIGNAL Logical_Operator_out10595_out1            : std_logic;
  SIGNAL Logical_Operator_out10596_out1            : std_logic;
  SIGNAL Logical_Operator_out10597_out1            : std_logic;
  SIGNAL Logical_Operator_out10598_out1            : std_logic;
  SIGNAL Logical_Operator_out10599_out1            : std_logic;
  SIGNAL Logical_Operator_out10600_out1            : std_logic;
  SIGNAL Logical_Operator_out10601_out1            : std_logic;
  SIGNAL Logical_Operator_out10602_out1            : std_logic;
  SIGNAL Logical_Operator_out10603_out1            : std_logic;
  SIGNAL Logical_Operator_out10604_out1            : std_logic;
  SIGNAL Logical_Operator_out10605_out1            : std_logic;
  SIGNAL Logical_Operator_out10606_out1            : std_logic;
  SIGNAL Logical_Operator_out10607_out1            : std_logic;
  SIGNAL Logical_Operator_out10608_out1            : std_logic;
  SIGNAL Logical_Operator_out10609_out1            : std_logic;
  SIGNAL Logical_Operator_out10610_out1            : std_logic;
  SIGNAL Logical_Operator_out10611_out1            : std_logic;
  SIGNAL Logical_Operator_out10612_out1            : std_logic;
  SIGNAL Logical_Operator_out10613_out1            : std_logic;
  SIGNAL Logical_Operator_out10614_out1            : std_logic;
  SIGNAL Logical_Operator_out10615_out1            : std_logic;
  SIGNAL Logical_Operator_out10616_out1            : std_logic;
  SIGNAL Logical_Operator_out10617_out1            : std_logic;
  SIGNAL Logical_Operator_out10618_out1            : std_logic;
  SIGNAL Logical_Operator_out10619_out1            : std_logic;
  SIGNAL Logical_Operator_out10620_out1            : std_logic;
  SIGNAL Logical_Operator_out10621_out1            : std_logic;
  SIGNAL Logical_Operator_out10622_out1            : std_logic;
  SIGNAL Logical_Operator_out10623_out1            : std_logic;
  SIGNAL Logical_Operator_out10624_out1            : std_logic;
  SIGNAL Logical_Operator_out10625_out1            : std_logic;
  SIGNAL Logical_Operator_out10626_out1            : std_logic;
  SIGNAL Logical_Operator_out10627_out1            : std_logic;
  SIGNAL Logical_Operator_out10628_out1            : std_logic;
  SIGNAL Logical_Operator_out10629_out1            : std_logic;
  SIGNAL Logical_Operator_out10630_out1            : std_logic;
  SIGNAL Logical_Operator_out10631_out1            : std_logic;
  SIGNAL Logical_Operator_out10632_out1            : std_logic;
  SIGNAL Logical_Operator_out10633_out1            : std_logic;
  SIGNAL Logical_Operator_out10634_out1            : std_logic;
  SIGNAL Logical_Operator_out10635_out1            : std_logic;
  SIGNAL Logical_Operator_out10636_out1            : std_logic;
  SIGNAL Logical_Operator_out10637_out1            : std_logic;
  SIGNAL Logical_Operator_out10638_out1            : std_logic;
  SIGNAL Logical_Operator_out10639_out1            : std_logic;
  SIGNAL Logical_Operator_out10640_out1            : std_logic;
  SIGNAL Logical_Operator_out10641_out1            : std_logic;
  SIGNAL Logical_Operator_out10642_out1            : std_logic;
  SIGNAL Logical_Operator_out10643_out1            : std_logic;
  SIGNAL Logical_Operator_out10644_out1            : std_logic;
  SIGNAL Logical_Operator_out10645_out1            : std_logic;
  SIGNAL Logical_Operator_out10646_out1            : std_logic;
  SIGNAL Logical_Operator_out10647_out1            : std_logic;
  SIGNAL Logical_Operator_out10648_out1            : std_logic;
  SIGNAL Logical_Operator_out10649_out1            : std_logic;
  SIGNAL Logical_Operator_out10650_out1            : std_logic;
  SIGNAL Logical_Operator_out10651_out1            : std_logic;
  SIGNAL Logical_Operator_out10652_out1            : std_logic;
  SIGNAL Logical_Operator_out10653_out1            : std_logic;
  SIGNAL Logical_Operator_out10654_out1            : std_logic;
  SIGNAL Logical_Operator_out10655_out1            : std_logic;
  SIGNAL Logical_Operator_out10656_out1            : std_logic;
  SIGNAL Logical_Operator_out10657_out1            : std_logic;
  SIGNAL Logical_Operator_out10658_out1            : std_logic;
  SIGNAL Logical_Operator_out10659_out1            : std_logic;
  SIGNAL Logical_Operator_out10660_out1            : std_logic;
  SIGNAL Logical_Operator_out10661_out1            : std_logic;
  SIGNAL Logical_Operator_out10662_out1            : std_logic;
  SIGNAL Logical_Operator_out10663_out1            : std_logic;
  SIGNAL Logical_Operator_out10664_out1            : std_logic;
  SIGNAL Logical_Operator_out10665_out1            : std_logic;
  SIGNAL Logical_Operator_out10666_out1            : std_logic;
  SIGNAL Logical_Operator_out10667_out1            : std_logic;
  SIGNAL Logical_Operator_out10668_out1            : std_logic;
  SIGNAL Logical_Operator_out10669_out1            : std_logic;
  SIGNAL Logical_Operator_out10670_out1            : std_logic;
  SIGNAL Logical_Operator_out10671_out1            : std_logic;
  SIGNAL Logical_Operator_out10672_out1            : std_logic;
  SIGNAL Logical_Operator_out10673_out1            : std_logic;
  SIGNAL Logical_Operator_out10674_out1            : std_logic;
  SIGNAL Logical_Operator_out10675_out1            : std_logic;
  SIGNAL Logical_Operator_out10676_out1            : std_logic;
  SIGNAL Logical_Operator_out10677_out1            : std_logic;
  SIGNAL Logical_Operator_out10678_out1            : std_logic;
  SIGNAL Logical_Operator_out10679_out1            : std_logic;
  SIGNAL Logical_Operator_out10680_out1            : std_logic;
  SIGNAL Logical_Operator_out10681_out1            : std_logic;
  SIGNAL Logical_Operator_out10682_out1            : std_logic;
  SIGNAL Logical_Operator_out10683_out1            : std_logic;
  SIGNAL Logical_Operator_out10684_out1            : std_logic;
  SIGNAL Logical_Operator_out10685_out1            : std_logic;
  SIGNAL Logical_Operator_out10686_out1            : std_logic;
  SIGNAL Logical_Operator_out10687_out1            : std_logic;
  SIGNAL Logical_Operator_out10688_out1            : std_logic;
  SIGNAL Logical_Operator_out10689_out1            : std_logic;
  SIGNAL Logical_Operator_out10690_out1            : std_logic;
  SIGNAL Logical_Operator_out10691_out1            : std_logic;
  SIGNAL Logical_Operator_out10692_out1            : std_logic;
  SIGNAL Logical_Operator_out10693_out1            : std_logic;
  SIGNAL Logical_Operator_out10694_out1            : std_logic;
  SIGNAL Logical_Operator_out10695_out1            : std_logic;
  SIGNAL Logical_Operator_out10696_out1            : std_logic;
  SIGNAL Logical_Operator_out10697_out1            : std_logic;
  SIGNAL Logical_Operator_out10698_out1            : std_logic;
  SIGNAL Logical_Operator_out10699_out1            : std_logic;
  SIGNAL Logical_Operator_out10700_out1            : std_logic;
  SIGNAL Logical_Operator_out10701_out1            : std_logic;
  SIGNAL Logical_Operator_out10702_out1            : std_logic;
  SIGNAL Logical_Operator_out10703_out1            : std_logic;
  SIGNAL Logical_Operator_out10704_out1            : std_logic;
  SIGNAL Logical_Operator_out10705_out1            : std_logic;
  SIGNAL Logical_Operator_out10706_out1            : std_logic;
  SIGNAL Logical_Operator_out10707_out1            : std_logic;
  SIGNAL Logical_Operator_out10708_out1            : std_logic;
  SIGNAL Logical_Operator_out10709_out1            : std_logic;
  SIGNAL Logical_Operator_out10710_out1            : std_logic;
  SIGNAL Logical_Operator_out10711_out1            : std_logic;
  SIGNAL Logical_Operator_out10712_out1            : std_logic;
  SIGNAL Logical_Operator_out10713_out1            : std_logic;
  SIGNAL Logical_Operator_out10714_out1            : std_logic;
  SIGNAL Logical_Operator_out10715_out1            : std_logic;
  SIGNAL Logical_Operator_out10716_out1            : std_logic;
  SIGNAL Logical_Operator_out10717_out1            : std_logic;
  SIGNAL Logical_Operator_out10718_out1            : std_logic;
  SIGNAL Logical_Operator_out10719_out1            : std_logic;
  SIGNAL Logical_Operator_out10720_out1            : std_logic;
  SIGNAL Logical_Operator_out10721_out1            : std_logic;
  SIGNAL Logical_Operator_out10722_out1            : std_logic;
  SIGNAL Logical_Operator_out10723_out1            : std_logic;
  SIGNAL Logical_Operator_out10724_out1            : std_logic;
  SIGNAL Logical_Operator_out10725_out1            : std_logic;
  SIGNAL Logical_Operator_out10726_out1            : std_logic;
  SIGNAL Logical_Operator_out10727_out1            : std_logic;
  SIGNAL Logical_Operator_out10728_out1            : std_logic;
  SIGNAL Logical_Operator_out10729_out1            : std_logic;
  SIGNAL Logical_Operator_out10730_out1            : std_logic;
  SIGNAL Logical_Operator_out10731_out1            : std_logic;
  SIGNAL Logical_Operator_out10732_out1            : std_logic;
  SIGNAL Logical_Operator_out10733_out1            : std_logic;
  SIGNAL Logical_Operator_out10734_out1            : std_logic;
  SIGNAL Logical_Operator_out10735_out1            : std_logic;
  SIGNAL Logical_Operator_out10736_out1            : std_logic;
  SIGNAL Logical_Operator_out10737_out1            : std_logic;
  SIGNAL Logical_Operator_out10738_out1            : std_logic;
  SIGNAL Logical_Operator_out10739_out1            : std_logic;
  SIGNAL Logical_Operator_out10740_out1            : std_logic;
  SIGNAL Logical_Operator_out10741_out1            : std_logic;
  SIGNAL Logical_Operator_out10742_out1            : std_logic;
  SIGNAL Logical_Operator_out10743_out1            : std_logic;
  SIGNAL Logical_Operator_out10744_out1            : std_logic;
  SIGNAL Logical_Operator_out10745_out1            : std_logic;
  SIGNAL Logical_Operator_out10746_out1            : std_logic;
  SIGNAL Logical_Operator_out10747_out1            : std_logic;
  SIGNAL Logical_Operator_out10748_out1            : std_logic;
  SIGNAL Logical_Operator_out10749_out1            : std_logic;
  SIGNAL Logical_Operator_out10750_out1            : std_logic;
  SIGNAL Logical_Operator_out10751_out1            : std_logic;
  SIGNAL Logical_Operator_out10752_out1            : std_logic;
  SIGNAL Logical_Operator_out10753_out1            : std_logic;
  SIGNAL Logical_Operator_out10754_out1            : std_logic;
  SIGNAL Logical_Operator_out10755_out1            : std_logic;
  SIGNAL Logical_Operator_out10756_out1            : std_logic;
  SIGNAL Logical_Operator_out10757_out1            : std_logic;
  SIGNAL Logical_Operator_out10758_out1            : std_logic;
  SIGNAL Logical_Operator_out10759_out1            : std_logic;
  SIGNAL Logical_Operator_out10760_out1            : std_logic;
  SIGNAL Logical_Operator_out10761_out1            : std_logic;
  SIGNAL Logical_Operator_out10762_out1            : std_logic;
  SIGNAL Logical_Operator_out10763_out1            : std_logic;
  SIGNAL Logical_Operator_out10764_out1            : std_logic;
  SIGNAL Logical_Operator_out10765_out1            : std_logic;
  SIGNAL Logical_Operator_out10766_out1            : std_logic;
  SIGNAL Logical_Operator_out10767_out1            : std_logic;
  SIGNAL Logical_Operator_out10768_out1            : std_logic;
  SIGNAL Logical_Operator_out10769_out1            : std_logic;
  SIGNAL Logical_Operator_out10770_out1            : std_logic;
  SIGNAL Logical_Operator_out10771_out1            : std_logic;
  SIGNAL Logical_Operator_out10772_out1            : std_logic;
  SIGNAL Logical_Operator_out10773_out1            : std_logic;
  SIGNAL Logical_Operator_out10774_out1            : std_logic;
  SIGNAL Logical_Operator_out10775_out1            : std_logic;
  SIGNAL Logical_Operator_out10776_out1            : std_logic;
  SIGNAL Logical_Operator_out10777_out1            : std_logic;
  SIGNAL Logical_Operator_out10778_out1            : std_logic;
  SIGNAL Logical_Operator_out10779_out1            : std_logic;
  SIGNAL Logical_Operator_out10780_out1            : std_logic;
  SIGNAL Logical_Operator_out10781_out1            : std_logic;
  SIGNAL Logical_Operator_out10782_out1            : std_logic;
  SIGNAL Logical_Operator_out10783_out1            : std_logic;
  SIGNAL Logical_Operator_out10784_out1            : std_logic;
  SIGNAL Logical_Operator_out10785_out1            : std_logic;
  SIGNAL Logical_Operator_out10786_out1            : std_logic;
  SIGNAL Logical_Operator_out10787_out1            : std_logic;
  SIGNAL Logical_Operator_out10788_out1            : std_logic;
  SIGNAL Logical_Operator_out10789_out1            : std_logic;
  SIGNAL Logical_Operator_out10790_out1            : std_logic;
  SIGNAL Logical_Operator_out10791_out1            : std_logic;
  SIGNAL Logical_Operator_out10792_out1            : std_logic;
  SIGNAL Logical_Operator_out10793_out1            : std_logic;
  SIGNAL Logical_Operator_out10794_out1            : std_logic;
  SIGNAL Logical_Operator_out10795_out1            : std_logic;
  SIGNAL Logical_Operator_out10796_out1            : std_logic;
  SIGNAL Logical_Operator_out10797_out1            : std_logic;
  SIGNAL Logical_Operator_out10798_out1            : std_logic;
  SIGNAL Logical_Operator_out10799_out1            : std_logic;
  SIGNAL Logical_Operator_out10800_out1            : std_logic;
  SIGNAL Logical_Operator_out10801_out1            : std_logic;
  SIGNAL Logical_Operator_out10802_out1            : std_logic;
  SIGNAL Logical_Operator_out10803_out1            : std_logic;
  SIGNAL Logical_Operator_out10804_out1            : std_logic;
  SIGNAL Logical_Operator_out10805_out1            : std_logic;
  SIGNAL Logical_Operator_out10806_out1            : std_logic;
  SIGNAL Logical_Operator_out10807_out1            : std_logic;
  SIGNAL Logical_Operator_out10808_out1            : std_logic;
  SIGNAL Logical_Operator_out10809_out1            : std_logic;
  SIGNAL Logical_Operator_out10810_out1            : std_logic;
  SIGNAL Logical_Operator_out10811_out1            : std_logic;
  SIGNAL Logical_Operator_out10812_out1            : std_logic;
  SIGNAL Logical_Operator_out10813_out1            : std_logic;
  SIGNAL Logical_Operator_out10814_out1            : std_logic;
  SIGNAL Logical_Operator_out10815_out1            : std_logic;
  SIGNAL Logical_Operator_out10816_out1            : std_logic;
  SIGNAL Logical_Operator_out10817_out1            : std_logic;
  SIGNAL Logical_Operator_out10818_out1            : std_logic;
  SIGNAL Logical_Operator_out10819_out1            : std_logic;
  SIGNAL Logical_Operator_out10820_out1            : std_logic;
  SIGNAL Logical_Operator_out10821_out1            : std_logic;
  SIGNAL Logical_Operator_out10822_out1            : std_logic;
  SIGNAL Logical_Operator_out10823_out1            : std_logic;
  SIGNAL Logical_Operator_out10824_out1            : std_logic;
  SIGNAL Logical_Operator_out10825_out1            : std_logic;
  SIGNAL Logical_Operator_out10826_out1            : std_logic;
  SIGNAL Logical_Operator_out10827_out1            : std_logic;
  SIGNAL Logical_Operator_out10828_out1            : std_logic;
  SIGNAL Logical_Operator_out10829_out1            : std_logic;
  SIGNAL Logical_Operator_out10830_out1            : std_logic;
  SIGNAL Logical_Operator_out10831_out1            : std_logic;
  SIGNAL Logical_Operator_out10832_out1            : std_logic;
  SIGNAL Logical_Operator_out10833_out1            : std_logic;
  SIGNAL Logical_Operator_out10834_out1            : std_logic;
  SIGNAL Logical_Operator_out10835_out1            : std_logic;
  SIGNAL Logical_Operator_out10836_out1            : std_logic;
  SIGNAL Logical_Operator_out10837_out1            : std_logic;
  SIGNAL Logical_Operator_out10838_out1            : std_logic;
  SIGNAL Logical_Operator_out10839_out1            : std_logic;
  SIGNAL Logical_Operator_out10840_out1            : std_logic;
  SIGNAL Logical_Operator_out10841_out1            : std_logic;
  SIGNAL Logical_Operator_out10842_out1            : std_logic;
  SIGNAL Logical_Operator_out10843_out1            : std_logic;
  SIGNAL Logical_Operator_out10844_out1            : std_logic;
  SIGNAL Logical_Operator_out10845_out1            : std_logic;
  SIGNAL Logical_Operator_out10846_out1            : std_logic;
  SIGNAL Logical_Operator_out10847_out1            : std_logic;
  SIGNAL Logical_Operator_out10848_out1            : std_logic;
  SIGNAL Logical_Operator_out10849_out1            : std_logic;
  SIGNAL Logical_Operator_out10850_out1            : std_logic;
  SIGNAL Logical_Operator_out10851_out1            : std_logic;
  SIGNAL Logical_Operator_out10852_out1            : std_logic;
  SIGNAL Logical_Operator_out10853_out1            : std_logic;
  SIGNAL Logical_Operator_out10854_out1            : std_logic;
  SIGNAL Logical_Operator_out10855_out1            : std_logic;
  SIGNAL Logical_Operator_out10856_out1            : std_logic;
  SIGNAL Logical_Operator_out10857_out1            : std_logic;
  SIGNAL Logical_Operator_out10858_out1            : std_logic;
  SIGNAL Logical_Operator_out10859_out1            : std_logic;
  SIGNAL Logical_Operator_out10860_out1            : std_logic;
  SIGNAL Logical_Operator_out10861_out1            : std_logic;
  SIGNAL Logical_Operator_out10862_out1            : std_logic;
  SIGNAL Logical_Operator_out10863_out1            : std_logic;
  SIGNAL Logical_Operator_out10864_out1            : std_logic;
  SIGNAL Logical_Operator_out10865_out1            : std_logic;
  SIGNAL Logical_Operator_out10866_out1            : std_logic;
  SIGNAL Logical_Operator_out10867_out1            : std_logic;
  SIGNAL Logical_Operator_out10868_out1            : std_logic;
  SIGNAL Logical_Operator_out10869_out1            : std_logic;
  SIGNAL Logical_Operator_out10870_out1            : std_logic;
  SIGNAL Logical_Operator_out10871_out1            : std_logic;
  SIGNAL Logical_Operator_out10872_out1            : std_logic;
  SIGNAL Logical_Operator_out10873_out1            : std_logic;
  SIGNAL Logical_Operator_out10874_out1            : std_logic;
  SIGNAL Logical_Operator_out10875_out1            : std_logic;
  SIGNAL Logical_Operator_out10876_out1            : std_logic;
  SIGNAL Logical_Operator_out10877_out1            : std_logic;
  SIGNAL Logical_Operator_out10878_out1            : std_logic;
  SIGNAL Logical_Operator_out10879_out1            : std_logic;
  SIGNAL Logical_Operator_out10880_out1            : std_logic;
  SIGNAL Logical_Operator_out10881_out1            : std_logic;
  SIGNAL Logical_Operator_out10882_out1            : std_logic;
  SIGNAL Logical_Operator_out10883_out1            : std_logic;
  SIGNAL Logical_Operator_out10884_out1            : std_logic;
  SIGNAL Logical_Operator_out10885_out1            : std_logic;
  SIGNAL Logical_Operator_out10886_out1            : std_logic;
  SIGNAL Logical_Operator_out10887_out1            : std_logic;
  SIGNAL Logical_Operator_out10888_out1            : std_logic;
  SIGNAL Logical_Operator_out10889_out1            : std_logic;
  SIGNAL Logical_Operator_out10890_out1            : std_logic;
  SIGNAL Logical_Operator_out10891_out1            : std_logic;
  SIGNAL Logical_Operator_out10892_out1            : std_logic;
  SIGNAL Logical_Operator_out10893_out1            : std_logic;
  SIGNAL Logical_Operator_out10894_out1            : std_logic;
  SIGNAL Logical_Operator_out10895_out1            : std_logic;
  SIGNAL Logical_Operator_out10896_out1            : std_logic;
  SIGNAL Logical_Operator_out10897_out1            : std_logic;
  SIGNAL Logical_Operator_out10898_out1            : std_logic;
  SIGNAL Logical_Operator_out10899_out1            : std_logic;
  SIGNAL Logical_Operator_out10900_out1            : std_logic;
  SIGNAL Logical_Operator_out10901_out1            : std_logic;
  SIGNAL Logical_Operator_out10902_out1            : std_logic;
  SIGNAL Logical_Operator_out10903_out1            : std_logic;
  SIGNAL Logical_Operator_out10904_out1            : std_logic;
  SIGNAL Logical_Operator_out10905_out1            : std_logic;
  SIGNAL Logical_Operator_out10906_out1            : std_logic;
  SIGNAL Logical_Operator_out10907_out1            : std_logic;
  SIGNAL Logical_Operator_out10908_out1            : std_logic;
  SIGNAL Logical_Operator_out10909_out1            : std_logic;
  SIGNAL Logical_Operator_out10910_out1            : std_logic;
  SIGNAL Logical_Operator_out10911_out1            : std_logic;
  SIGNAL Logical_Operator_out10912_out1            : std_logic;
  SIGNAL Logical_Operator_out10913_out1            : std_logic;
  SIGNAL Logical_Operator_out10914_out1            : std_logic;
  SIGNAL Logical_Operator_out10915_out1            : std_logic;
  SIGNAL Logical_Operator_out10916_out1            : std_logic;
  SIGNAL Logical_Operator_out10917_out1            : std_logic;
  SIGNAL Logical_Operator_out10918_out1            : std_logic;
  SIGNAL Logical_Operator_out10919_out1            : std_logic;
  SIGNAL Logical_Operator_out10920_out1            : std_logic;
  SIGNAL Logical_Operator_out10921_out1            : std_logic;
  SIGNAL Logical_Operator_out10922_out1            : std_logic;
  SIGNAL Logical_Operator_out10923_out1            : std_logic;
  SIGNAL Logical_Operator_out10924_out1            : std_logic;
  SIGNAL Logical_Operator_out10925_out1            : std_logic;
  SIGNAL Logical_Operator_out10926_out1            : std_logic;
  SIGNAL Logical_Operator_out10927_out1            : std_logic;
  SIGNAL Logical_Operator_out10928_out1            : std_logic;
  SIGNAL Logical_Operator_out10929_out1            : std_logic;
  SIGNAL Logical_Operator_out10930_out1            : std_logic;
  SIGNAL Logical_Operator_out10931_out1            : std_logic;
  SIGNAL Logical_Operator_out10932_out1            : std_logic;
  SIGNAL Logical_Operator_out10933_out1            : std_logic;
  SIGNAL Logical_Operator_out10934_out1            : std_logic;
  SIGNAL Logical_Operator_out10935_out1            : std_logic;
  SIGNAL Logical_Operator_out10936_out1            : std_logic;
  SIGNAL Logical_Operator_out10937_out1            : std_logic;
  SIGNAL Logical_Operator_out10938_out1            : std_logic;
  SIGNAL Logical_Operator_out10939_out1            : std_logic;
  SIGNAL Logical_Operator_out10940_out1            : std_logic;
  SIGNAL Logical_Operator_out10941_out1            : std_logic;
  SIGNAL Logical_Operator_out10942_out1            : std_logic;
  SIGNAL Logical_Operator_out10943_out1            : std_logic;
  SIGNAL Logical_Operator_out10944_out1            : std_logic;
  SIGNAL Logical_Operator_out10945_out1            : std_logic;
  SIGNAL Logical_Operator_out10946_out1            : std_logic;
  SIGNAL Logical_Operator_out10947_out1            : std_logic;
  SIGNAL Logical_Operator_out10948_out1            : std_logic;
  SIGNAL Logical_Operator_out10949_out1            : std_logic;
  SIGNAL Logical_Operator_out10950_out1            : std_logic;
  SIGNAL Logical_Operator_out10951_out1            : std_logic;
  SIGNAL Logical_Operator_out10952_out1            : std_logic;
  SIGNAL Logical_Operator_out10953_out1            : std_logic;
  SIGNAL Logical_Operator_out10954_out1            : std_logic;
  SIGNAL Logical_Operator_out10955_out1            : std_logic;
  SIGNAL Logical_Operator_out10956_out1            : std_logic;
  SIGNAL Logical_Operator_out10957_out1            : std_logic;
  SIGNAL Logical_Operator_out10958_out1            : std_logic;
  SIGNAL Logical_Operator_out10959_out1            : std_logic;
  SIGNAL Logical_Operator_out10960_out1            : std_logic;
  SIGNAL Logical_Operator_out10961_out1            : std_logic;
  SIGNAL Logical_Operator_out10962_out1            : std_logic;
  SIGNAL Logical_Operator_out10963_out1            : std_logic;
  SIGNAL Logical_Operator_out10964_out1            : std_logic;
  SIGNAL Logical_Operator_out10965_out1            : std_logic;
  SIGNAL Logical_Operator_out10966_out1            : std_logic;
  SIGNAL Logical_Operator_out10967_out1            : std_logic;
  SIGNAL Logical_Operator_out10968_out1            : std_logic;
  SIGNAL Logical_Operator_out10969_out1            : std_logic;
  SIGNAL Logical_Operator_out10970_out1            : std_logic;
  SIGNAL Logical_Operator_out10971_out1            : std_logic;
  SIGNAL Logical_Operator_out10972_out1            : std_logic;
  SIGNAL Logical_Operator_out10973_out1            : std_logic;
  SIGNAL Logical_Operator_out10974_out1            : std_logic;
  SIGNAL Logical_Operator_out10975_out1            : std_logic;
  SIGNAL Logical_Operator_out10976_out1            : std_logic;
  SIGNAL Logical_Operator_out10977_out1            : std_logic;
  SIGNAL Logical_Operator_out10978_out1            : std_logic;
  SIGNAL Logical_Operator_out10979_out1            : std_logic;
  SIGNAL Logical_Operator_out10980_out1            : std_logic;
  SIGNAL Logical_Operator_out10981_out1            : std_logic;
  SIGNAL Logical_Operator_out10982_out1            : std_logic;
  SIGNAL Logical_Operator_out10983_out1            : std_logic;
  SIGNAL Logical_Operator_out10984_out1            : std_logic;
  SIGNAL Logical_Operator_out10985_out1            : std_logic;
  SIGNAL Logical_Operator_out10986_out1            : std_logic;
  SIGNAL Logical_Operator_out10987_out1            : std_logic;
  SIGNAL Logical_Operator_out10988_out1            : std_logic;
  SIGNAL Logical_Operator_out10989_out1            : std_logic;
  SIGNAL Logical_Operator_out10990_out1            : std_logic;
  SIGNAL Logical_Operator_out10991_out1            : std_logic;
  SIGNAL Logical_Operator_out10992_out1            : std_logic;
  SIGNAL Logical_Operator_out10993_out1            : std_logic;
  SIGNAL Logical_Operator_out10994_out1            : std_logic;
  SIGNAL Logical_Operator_out10995_out1            : std_logic;
  SIGNAL Logical_Operator_out10996_out1            : std_logic;
  SIGNAL Logical_Operator_out10997_out1            : std_logic;
  SIGNAL Logical_Operator_out10998_out1            : std_logic;
  SIGNAL Logical_Operator_out10999_out1            : std_logic;
  SIGNAL Logical_Operator_out11000_out1            : std_logic;
  SIGNAL Logical_Operator_out11001_out1            : std_logic;
  SIGNAL Logical_Operator_out11002_out1            : std_logic;
  SIGNAL Logical_Operator_out11003_out1            : std_logic;
  SIGNAL Logical_Operator_out11004_out1            : std_logic;
  SIGNAL Logical_Operator_out11005_out1            : std_logic;
  SIGNAL Logical_Operator_out11006_out1            : std_logic;
  SIGNAL Logical_Operator_out11007_out1            : std_logic;
  SIGNAL Logical_Operator_out11008_out1            : std_logic;
  SIGNAL Logical_Operator_out11009_out1            : std_logic;
  SIGNAL Logical_Operator_out11010_out1            : std_logic;
  SIGNAL Logical_Operator_out11011_out1            : std_logic;
  SIGNAL Logical_Operator_out11012_out1            : std_logic;
  SIGNAL Logical_Operator_out11013_out1            : std_logic;
  SIGNAL Logical_Operator_out11014_out1            : std_logic;
  SIGNAL Logical_Operator_out11015_out1            : std_logic;
  SIGNAL Logical_Operator_out11016_out1            : std_logic;
  SIGNAL Logical_Operator_out11017_out1            : std_logic;
  SIGNAL Logical_Operator_out11018_out1            : std_logic;
  SIGNAL Logical_Operator_out11019_out1            : std_logic;
  SIGNAL Logical_Operator_out11020_out1            : std_logic;
  SIGNAL Logical_Operator_out11021_out1            : std_logic;
  SIGNAL Logical_Operator_out11022_out1            : std_logic;
  SIGNAL Logical_Operator_out11023_out1            : std_logic;
  SIGNAL Logical_Operator_out11024_out1            : std_logic;
  SIGNAL Logical_Operator_out11025_out1            : std_logic;
  SIGNAL Logical_Operator_out11026_out1            : std_logic;
  SIGNAL Logical_Operator_out11027_out1            : std_logic;
  SIGNAL Logical_Operator_out11028_out1            : std_logic;
  SIGNAL Logical_Operator_out11029_out1            : std_logic;
  SIGNAL Logical_Operator_out11030_out1            : std_logic;
  SIGNAL Logical_Operator_out11031_out1            : std_logic;
  SIGNAL Logical_Operator_out11032_out1            : std_logic;
  SIGNAL Logical_Operator_out11033_out1            : std_logic;
  SIGNAL Logical_Operator_out11034_out1            : std_logic;
  SIGNAL Logical_Operator_out11035_out1            : std_logic;
  SIGNAL Logical_Operator_out11036_out1            : std_logic;
  SIGNAL Logical_Operator_out11037_out1            : std_logic;
  SIGNAL Logical_Operator_out11038_out1            : std_logic;
  SIGNAL Logical_Operator_out11039_out1            : std_logic;
  SIGNAL Logical_Operator_out11040_out1            : std_logic;
  SIGNAL Logical_Operator_out11041_out1            : std_logic;
  SIGNAL Logical_Operator_out11042_out1            : std_logic;
  SIGNAL Logical_Operator_out11043_out1            : std_logic;
  SIGNAL Logical_Operator_out11044_out1            : std_logic;
  SIGNAL Logical_Operator_out11045_out1            : std_logic;
  SIGNAL Logical_Operator_out11046_out1            : std_logic;
  SIGNAL Logical_Operator_out11047_out1            : std_logic;
  SIGNAL Logical_Operator_out11048_out1            : std_logic;
  SIGNAL Logical_Operator_out11049_out1            : std_logic;
  SIGNAL Logical_Operator_out11050_out1            : std_logic;
  SIGNAL Logical_Operator_out11051_out1            : std_logic;
  SIGNAL Logical_Operator_out11052_out1            : std_logic;
  SIGNAL Logical_Operator_out11053_out1            : std_logic;
  SIGNAL Logical_Operator_out11054_out1            : std_logic;
  SIGNAL Logical_Operator_out11055_out1            : std_logic;
  SIGNAL Logical_Operator_out11056_out1            : std_logic;
  SIGNAL Logical_Operator_out11057_out1            : std_logic;
  SIGNAL Logical_Operator_out11058_out1            : std_logic;
  SIGNAL Logical_Operator_out11059_out1            : std_logic;
  SIGNAL Logical_Operator_out11060_out1            : std_logic;
  SIGNAL Logical_Operator_out11061_out1            : std_logic;
  SIGNAL Logical_Operator_out11062_out1            : std_logic;
  SIGNAL Logical_Operator_out11063_out1            : std_logic;
  SIGNAL Logical_Operator_out11064_out1            : std_logic;
  SIGNAL Logical_Operator_out11065_out1            : std_logic;
  SIGNAL Logical_Operator_out11066_out1            : std_logic;
  SIGNAL Logical_Operator_out11067_out1            : std_logic;
  SIGNAL Logical_Operator_out11068_out1            : std_logic;
  SIGNAL Logical_Operator_out11069_out1            : std_logic;
  SIGNAL Logical_Operator_out11070_out1            : std_logic;
  SIGNAL Logical_Operator_out11071_out1            : std_logic;
  SIGNAL Logical_Operator_out11072_out1            : std_logic;
  SIGNAL Logical_Operator_out11073_out1            : std_logic;
  SIGNAL Logical_Operator_out11074_out1            : std_logic;
  SIGNAL Logical_Operator_out11075_out1            : std_logic;
  SIGNAL Logical_Operator_out11076_out1            : std_logic;
  SIGNAL Logical_Operator_out11077_out1            : std_logic;
  SIGNAL Logical_Operator_out11078_out1            : std_logic;
  SIGNAL Logical_Operator_out11079_out1            : std_logic;
  SIGNAL Logical_Operator_out11080_out1            : std_logic;
  SIGNAL Logical_Operator_out11081_out1            : std_logic;
  SIGNAL Logical_Operator_out11082_out1            : std_logic;
  SIGNAL Logical_Operator_out11083_out1            : std_logic;
  SIGNAL Logical_Operator_out11084_out1            : std_logic;
  SIGNAL Logical_Operator_out11085_out1            : std_logic;
  SIGNAL Logical_Operator_out11086_out1            : std_logic;
  SIGNAL Logical_Operator_out11087_out1            : std_logic;
  SIGNAL Logical_Operator_out11088_out1            : std_logic;
  SIGNAL Logical_Operator_out11089_out1            : std_logic;
  SIGNAL Logical_Operator_out11090_out1            : std_logic;
  SIGNAL Logical_Operator_out11091_out1            : std_logic;
  SIGNAL Logical_Operator_out11092_out1            : std_logic;
  SIGNAL Logical_Operator_out11093_out1            : std_logic;
  SIGNAL Logical_Operator_out11094_out1            : std_logic;
  SIGNAL Logical_Operator_out11095_out1            : std_logic;
  SIGNAL Logical_Operator_out11096_out1            : std_logic;
  SIGNAL Logical_Operator_out11097_out1            : std_logic;
  SIGNAL Logical_Operator_out11098_out1            : std_logic;
  SIGNAL Logical_Operator_out11099_out1            : std_logic;
  SIGNAL Logical_Operator_out11100_out1            : std_logic;
  SIGNAL Logical_Operator_out11101_out1            : std_logic;
  SIGNAL Logical_Operator_out11102_out1            : std_logic;
  SIGNAL Logical_Operator_out11103_out1            : std_logic;
  SIGNAL Logical_Operator_out11104_out1            : std_logic;
  SIGNAL Logical_Operator_out11105_out1            : std_logic;
  SIGNAL Logical_Operator_out11106_out1            : std_logic;
  SIGNAL Logical_Operator_out11107_out1            : std_logic;
  SIGNAL Logical_Operator_out11108_out1            : std_logic;
  SIGNAL Logical_Operator_out11109_out1            : std_logic;
  SIGNAL Logical_Operator_out11110_out1            : std_logic;
  SIGNAL Logical_Operator_out11111_out1            : std_logic;
  SIGNAL Logical_Operator_out11112_out1            : std_logic;
  SIGNAL Logical_Operator_out11113_out1            : std_logic;
  SIGNAL Logical_Operator_out11114_out1            : std_logic;
  SIGNAL Logical_Operator_out11115_out1            : std_logic;
  SIGNAL Logical_Operator_out11116_out1            : std_logic;
  SIGNAL Logical_Operator_out11117_out1            : std_logic;
  SIGNAL Logical_Operator_out11118_out1            : std_logic;
  SIGNAL Logical_Operator_out11119_out1            : std_logic;
  SIGNAL Logical_Operator_out11120_out1            : std_logic;
  SIGNAL Logical_Operator_out11121_out1            : std_logic;
  SIGNAL Logical_Operator_out11122_out1            : std_logic;
  SIGNAL Logical_Operator_out11123_out1            : std_logic;
  SIGNAL Logical_Operator_out11124_out1            : std_logic;
  SIGNAL Logical_Operator_out11125_out1            : std_logic;
  SIGNAL Logical_Operator_out11126_out1            : std_logic;
  SIGNAL Logical_Operator_out11127_out1            : std_logic;
  SIGNAL Logical_Operator_out11128_out1            : std_logic;
  SIGNAL Logical_Operator_out11129_out1            : std_logic;
  SIGNAL Logical_Operator_out11130_out1            : std_logic;
  SIGNAL Logical_Operator_out11131_out1            : std_logic;
  SIGNAL Logical_Operator_out11132_out1            : std_logic;
  SIGNAL Logical_Operator_out11133_out1            : std_logic;
  SIGNAL Logical_Operator_out11134_out1            : std_logic;
  SIGNAL Logical_Operator_out11135_out1            : std_logic;
  SIGNAL Logical_Operator_out11136_out1            : std_logic;
  SIGNAL Logical_Operator_out11137_out1            : std_logic;
  SIGNAL Logical_Operator_out11138_out1            : std_logic;
  SIGNAL Logical_Operator_out11139_out1            : std_logic;
  SIGNAL Logical_Operator_out11140_out1            : std_logic;
  SIGNAL Logical_Operator_out11141_out1            : std_logic;
  SIGNAL Logical_Operator_out11142_out1            : std_logic;
  SIGNAL Logical_Operator_out11143_out1            : std_logic;
  SIGNAL Logical_Operator_out11144_out1            : std_logic;
  SIGNAL Logical_Operator_out11145_out1            : std_logic;
  SIGNAL Logical_Operator_out11146_out1            : std_logic;
  SIGNAL Logical_Operator_out11147_out1            : std_logic;
  SIGNAL Logical_Operator_out11148_out1            : std_logic;
  SIGNAL Logical_Operator_out11149_out1            : std_logic;
  SIGNAL Logical_Operator_out11150_out1            : std_logic;
  SIGNAL Logical_Operator_out11151_out1            : std_logic;
  SIGNAL Logical_Operator_out11152_out1            : std_logic;
  SIGNAL Logical_Operator_out11153_out1            : std_logic;
  SIGNAL Logical_Operator_out11154_out1            : std_logic;
  SIGNAL Logical_Operator_out11155_out1            : std_logic;
  SIGNAL Logical_Operator_out11156_out1            : std_logic;
  SIGNAL Logical_Operator_out11157_out1            : std_logic;
  SIGNAL Logical_Operator_out11158_out1            : std_logic;
  SIGNAL Logical_Operator_out11159_out1            : std_logic;
  SIGNAL Logical_Operator_out11160_out1            : std_logic;
  SIGNAL Logical_Operator_out11161_out1            : std_logic;
  SIGNAL Logical_Operator_out11162_out1            : std_logic;
  SIGNAL Logical_Operator_out11163_out1            : std_logic;
  SIGNAL Logical_Operator_out11164_out1            : std_logic;
  SIGNAL Logical_Operator_out11165_out1            : std_logic;
  SIGNAL Logical_Operator_out11166_out1            : std_logic;
  SIGNAL Logical_Operator_out11167_out1            : std_logic;
  SIGNAL Logical_Operator_out11168_out1            : std_logic;
  SIGNAL Logical_Operator_out11169_out1            : std_logic;
  SIGNAL Logical_Operator_out11170_out1            : std_logic;
  SIGNAL Logical_Operator_out11171_out1            : std_logic;
  SIGNAL Logical_Operator_out11172_out1            : std_logic;
  SIGNAL Logical_Operator_out11173_out1            : std_logic;
  SIGNAL Logical_Operator_out11174_out1            : std_logic;
  SIGNAL Logical_Operator_out11175_out1            : std_logic;
  SIGNAL Logical_Operator_out11176_out1            : std_logic;
  SIGNAL Logical_Operator_out11177_out1            : std_logic;
  SIGNAL Logical_Operator_out11178_out1            : std_logic;
  SIGNAL Logical_Operator_out11179_out1            : std_logic;
  SIGNAL Logical_Operator_out11180_out1            : std_logic;
  SIGNAL Logical_Operator_out11181_out1            : std_logic;
  SIGNAL Logical_Operator_out11182_out1            : std_logic;
  SIGNAL Logical_Operator_out11183_out1            : std_logic;
  SIGNAL Logical_Operator_out11184_out1            : std_logic;
  SIGNAL Logical_Operator_out11185_out1            : std_logic;
  SIGNAL Logical_Operator_out11186_out1            : std_logic;
  SIGNAL Logical_Operator_out11187_out1            : std_logic;
  SIGNAL Logical_Operator_out11188_out1            : std_logic;
  SIGNAL Logical_Operator_out11189_out1            : std_logic;
  SIGNAL Logical_Operator_out11190_out1            : std_logic;
  SIGNAL Logical_Operator_out11191_out1            : std_logic;
  SIGNAL Logical_Operator_out11192_out1            : std_logic;
  SIGNAL Logical_Operator_out11193_out1            : std_logic;
  SIGNAL Logical_Operator_out11194_out1            : std_logic;
  SIGNAL Logical_Operator_out11195_out1            : std_logic;
  SIGNAL Logical_Operator_out11196_out1            : std_logic;
  SIGNAL Logical_Operator_out11197_out1            : std_logic;
  SIGNAL Logical_Operator_out11198_out1            : std_logic;
  SIGNAL Logical_Operator_out11199_out1            : std_logic;
  SIGNAL Logical_Operator_out11200_out1            : std_logic;
  SIGNAL Logical_Operator_out11201_out1            : std_logic;
  SIGNAL Logical_Operator_out11202_out1            : std_logic;
  SIGNAL Logical_Operator_out11203_out1            : std_logic;
  SIGNAL Logical_Operator_out11204_out1            : std_logic;
  SIGNAL Logical_Operator_out11205_out1            : std_logic;
  SIGNAL Logical_Operator_out11206_out1            : std_logic;
  SIGNAL Logical_Operator_out11207_out1            : std_logic;
  SIGNAL Logical_Operator_out11208_out1            : std_logic;
  SIGNAL Logical_Operator_out11209_out1            : std_logic;
  SIGNAL Logical_Operator_out11210_out1            : std_logic;
  SIGNAL Logical_Operator_out11211_out1            : std_logic;
  SIGNAL Logical_Operator_out11212_out1            : std_logic;
  SIGNAL Logical_Operator_out11213_out1            : std_logic;
  SIGNAL Logical_Operator_out11214_out1            : std_logic;
  SIGNAL Logical_Operator_out11215_out1            : std_logic;
  SIGNAL Logical_Operator_out11216_out1            : std_logic;
  SIGNAL Logical_Operator_out11217_out1            : std_logic;
  SIGNAL Logical_Operator_out11218_out1            : std_logic;
  SIGNAL Logical_Operator_out11219_out1            : std_logic;
  SIGNAL Logical_Operator_out11220_out1            : std_logic;
  SIGNAL Logical_Operator_out11221_out1            : std_logic;
  SIGNAL Logical_Operator_out11222_out1            : std_logic;
  SIGNAL Logical_Operator_out11223_out1            : std_logic;
  SIGNAL Logical_Operator_out11224_out1            : std_logic;
  SIGNAL Logical_Operator_out11225_out1            : std_logic;
  SIGNAL Logical_Operator_out11226_out1            : std_logic;
  SIGNAL Logical_Operator_out11227_out1            : std_logic;
  SIGNAL Logical_Operator_out11228_out1            : std_logic;
  SIGNAL Logical_Operator_out11229_out1            : std_logic;
  SIGNAL Logical_Operator_out11230_out1            : std_logic;
  SIGNAL Logical_Operator_out11231_out1            : std_logic;
  SIGNAL Logical_Operator_out11232_out1            : std_logic;
  SIGNAL Logical_Operator_out11233_out1            : std_logic;
  SIGNAL Logical_Operator_out11234_out1            : std_logic;
  SIGNAL Logical_Operator_out11235_out1            : std_logic;
  SIGNAL Logical_Operator_out11236_out1            : std_logic;
  SIGNAL Logical_Operator_out11237_out1            : std_logic;
  SIGNAL Logical_Operator_out11238_out1            : std_logic;
  SIGNAL Logical_Operator_out11239_out1            : std_logic;
  SIGNAL Logical_Operator_out11240_out1            : std_logic;
  SIGNAL Logical_Operator_out11241_out1            : std_logic;
  SIGNAL Logical_Operator_out11242_out1            : std_logic;
  SIGNAL Logical_Operator_out11243_out1            : std_logic;
  SIGNAL Logical_Operator_out11244_out1            : std_logic;
  SIGNAL Logical_Operator_out11245_out1            : std_logic;
  SIGNAL Logical_Operator_out11246_out1            : std_logic;
  SIGNAL Logical_Operator_out11247_out1            : std_logic;
  SIGNAL Logical_Operator_out11248_out1            : std_logic;
  SIGNAL Logical_Operator_out11249_out1            : std_logic;
  SIGNAL Logical_Operator_out11250_out1            : std_logic;
  SIGNAL Logical_Operator_out11251_out1            : std_logic;
  SIGNAL Logical_Operator_out11252_out1            : std_logic;
  SIGNAL Logical_Operator_out11253_out1            : std_logic;
  SIGNAL Logical_Operator_out11254_out1            : std_logic;
  SIGNAL Logical_Operator_out11255_out1            : std_logic;
  SIGNAL Logical_Operator_out11256_out1            : std_logic;
  SIGNAL Logical_Operator_out11257_out1            : std_logic;
  SIGNAL Logical_Operator_out11258_out1            : std_logic;
  SIGNAL Logical_Operator_out11259_out1            : std_logic;
  SIGNAL Logical_Operator_out11260_out1            : std_logic;
  SIGNAL Logical_Operator_out11261_out1            : std_logic;
  SIGNAL Logical_Operator_out11262_out1            : std_logic;
  SIGNAL Logical_Operator_out11263_out1            : std_logic;
  SIGNAL Logical_Operator_out11264_out1            : std_logic;

BEGIN

  Logical_Operator_out1_out1 <= in1 XOR in2;

  Logical_Operator_out2_out1 <= in3 XOR in4;

  Logical_Operator_out3_out1 <= in5 XOR in6;

  Logical_Operator_out4_out1 <= in7 XOR in8;

  Logical_Operator_out5_out1 <= in9 XOR in10;

  Logical_Operator_out6_out1 <= in11 XOR in12;

  Logical_Operator_out7_out1 <= in13 XOR in14;

  Logical_Operator_out8_out1 <= in15 XOR in16;

  Logical_Operator_out9_out1 <= in17 XOR in18;

  Logical_Operator_out10_out1 <= in19 XOR in20;

  Logical_Operator_out11_out1 <= in21 XOR in22;

  Logical_Operator_out12_out1 <= in23 XOR in24;

  Logical_Operator_out13_out1 <= in25 XOR in26;

  Logical_Operator_out14_out1 <= in27 XOR in28;

  Logical_Operator_out15_out1 <= in29 XOR in30;

  Logical_Operator_out16_out1 <= in31 XOR in32;

  Logical_Operator_out17_out1 <= in33 XOR in34;

  Logical_Operator_out18_out1 <= in35 XOR in36;

  Logical_Operator_out19_out1 <= in37 XOR in38;

  Logical_Operator_out20_out1 <= in39 XOR in40;

  Logical_Operator_out21_out1 <= in41 XOR in42;

  Logical_Operator_out22_out1 <= in43 XOR in44;

  Logical_Operator_out23_out1 <= in45 XOR in46;

  Logical_Operator_out24_out1 <= in47 XOR in48;

  Logical_Operator_out25_out1 <= in49 XOR in50;

  Logical_Operator_out26_out1 <= in51 XOR in52;

  Logical_Operator_out27_out1 <= in53 XOR in54;

  Logical_Operator_out28_out1 <= in55 XOR in56;

  Logical_Operator_out29_out1 <= in57 XOR in58;

  Logical_Operator_out30_out1 <= in59 XOR in60;

  Logical_Operator_out31_out1 <= in61 XOR in62;

  Logical_Operator_out32_out1 <= in63 XOR in64;

  Logical_Operator_out33_out1 <= in65 XOR in66;

  Logical_Operator_out34_out1 <= in67 XOR in68;

  Logical_Operator_out35_out1 <= in69 XOR in70;

  Logical_Operator_out36_out1 <= in71 XOR in72;

  Logical_Operator_out37_out1 <= in73 XOR in74;

  Logical_Operator_out38_out1 <= in75 XOR in76;

  Logical_Operator_out39_out1 <= in77 XOR in78;

  Logical_Operator_out40_out1 <= in79 XOR in80;

  Logical_Operator_out41_out1 <= in81 XOR in82;

  Logical_Operator_out42_out1 <= in83 XOR in84;

  Logical_Operator_out43_out1 <= in85 XOR in86;

  Logical_Operator_out44_out1 <= in87 XOR in88;

  Logical_Operator_out45_out1 <= in89 XOR in90;

  Logical_Operator_out46_out1 <= in91 XOR in92;

  Logical_Operator_out47_out1 <= in93 XOR in94;

  Logical_Operator_out48_out1 <= in95 XOR in96;

  Logical_Operator_out49_out1 <= in97 XOR in98;

  Logical_Operator_out50_out1 <= in99 XOR in100;

  Logical_Operator_out51_out1 <= in101 XOR in102;

  Logical_Operator_out52_out1 <= in103 XOR in104;

  Logical_Operator_out53_out1 <= in105 XOR in106;

  Logical_Operator_out54_out1 <= in107 XOR in108;

  Logical_Operator_out55_out1 <= in109 XOR in110;

  Logical_Operator_out56_out1 <= in111 XOR in112;

  Logical_Operator_out57_out1 <= in113 XOR in114;

  Logical_Operator_out58_out1 <= in115 XOR in116;

  Logical_Operator_out59_out1 <= in117 XOR in118;

  Logical_Operator_out60_out1 <= in119 XOR in120;

  Logical_Operator_out61_out1 <= in121 XOR in122;

  Logical_Operator_out62_out1 <= in123 XOR in124;

  Logical_Operator_out63_out1 <= in125 XOR in126;

  Logical_Operator_out64_out1 <= in127 XOR in128;

  Logical_Operator_out65_out1 <= in129 XOR in130;

  Logical_Operator_out66_out1 <= in131 XOR in132;

  Logical_Operator_out67_out1 <= in133 XOR in134;

  Logical_Operator_out68_out1 <= in135 XOR in136;

  Logical_Operator_out69_out1 <= in137 XOR in138;

  Logical_Operator_out70_out1 <= in139 XOR in140;

  Logical_Operator_out71_out1 <= in141 XOR in142;

  Logical_Operator_out72_out1 <= in143 XOR in144;

  Logical_Operator_out73_out1 <= in145 XOR in146;

  Logical_Operator_out74_out1 <= in147 XOR in148;

  Logical_Operator_out75_out1 <= in149 XOR in150;

  Logical_Operator_out76_out1 <= in151 XOR in152;

  Logical_Operator_out77_out1 <= in153 XOR in154;

  Logical_Operator_out78_out1 <= in155 XOR in156;

  Logical_Operator_out79_out1 <= in157 XOR in158;

  Logical_Operator_out80_out1 <= in159 XOR in160;

  Logical_Operator_out81_out1 <= in161 XOR in162;

  Logical_Operator_out82_out1 <= in163 XOR in164;

  Logical_Operator_out83_out1 <= in165 XOR in166;

  Logical_Operator_out84_out1 <= in167 XOR in168;

  Logical_Operator_out85_out1 <= in169 XOR in170;

  Logical_Operator_out86_out1 <= in171 XOR in172;

  Logical_Operator_out87_out1 <= in173 XOR in174;

  Logical_Operator_out88_out1 <= in175 XOR in176;

  Logical_Operator_out89_out1 <= in177 XOR in178;

  Logical_Operator_out90_out1 <= in179 XOR in180;

  Logical_Operator_out91_out1 <= in181 XOR in182;

  Logical_Operator_out92_out1 <= in183 XOR in184;

  Logical_Operator_out93_out1 <= in185 XOR in186;

  Logical_Operator_out94_out1 <= in187 XOR in188;

  Logical_Operator_out95_out1 <= in189 XOR in190;

  Logical_Operator_out96_out1 <= in191 XOR in192;

  Logical_Operator_out97_out1 <= in193 XOR in194;

  Logical_Operator_out98_out1 <= in195 XOR in196;

  Logical_Operator_out99_out1 <= in197 XOR in198;

  Logical_Operator_out100_out1 <= in199 XOR in200;

  Logical_Operator_out101_out1 <= in201 XOR in202;

  Logical_Operator_out102_out1 <= in203 XOR in204;

  Logical_Operator_out103_out1 <= in205 XOR in206;

  Logical_Operator_out104_out1 <= in207 XOR in208;

  Logical_Operator_out105_out1 <= in209 XOR in210;

  Logical_Operator_out106_out1 <= in211 XOR in212;

  Logical_Operator_out107_out1 <= in213 XOR in214;

  Logical_Operator_out108_out1 <= in215 XOR in216;

  Logical_Operator_out109_out1 <= in217 XOR in218;

  Logical_Operator_out110_out1 <= in219 XOR in220;

  Logical_Operator_out111_out1 <= in221 XOR in222;

  Logical_Operator_out112_out1 <= in223 XOR in224;

  Logical_Operator_out113_out1 <= in225 XOR in226;

  Logical_Operator_out114_out1 <= in227 XOR in228;

  Logical_Operator_out115_out1 <= in229 XOR in230;

  Logical_Operator_out116_out1 <= in231 XOR in232;

  Logical_Operator_out117_out1 <= in233 XOR in234;

  Logical_Operator_out118_out1 <= in235 XOR in236;

  Logical_Operator_out119_out1 <= in237 XOR in238;

  Logical_Operator_out120_out1 <= in239 XOR in240;

  Logical_Operator_out121_out1 <= in241 XOR in242;

  Logical_Operator_out122_out1 <= in243 XOR in244;

  Logical_Operator_out123_out1 <= in245 XOR in246;

  Logical_Operator_out124_out1 <= in247 XOR in248;

  Logical_Operator_out125_out1 <= in249 XOR in250;

  Logical_Operator_out126_out1 <= in251 XOR in252;

  Logical_Operator_out127_out1 <= in253 XOR in254;

  Logical_Operator_out128_out1 <= in255 XOR in256;

  Logical_Operator_out129_out1 <= in257 XOR in258;

  Logical_Operator_out130_out1 <= in259 XOR in260;

  Logical_Operator_out131_out1 <= in261 XOR in262;

  Logical_Operator_out132_out1 <= in263 XOR in264;

  Logical_Operator_out133_out1 <= in265 XOR in266;

  Logical_Operator_out134_out1 <= in267 XOR in268;

  Logical_Operator_out135_out1 <= in269 XOR in270;

  Logical_Operator_out136_out1 <= in271 XOR in272;

  Logical_Operator_out137_out1 <= in273 XOR in274;

  Logical_Operator_out138_out1 <= in275 XOR in276;

  Logical_Operator_out139_out1 <= in277 XOR in278;

  Logical_Operator_out140_out1 <= in279 XOR in280;

  Logical_Operator_out141_out1 <= in281 XOR in282;

  Logical_Operator_out142_out1 <= in283 XOR in284;

  Logical_Operator_out143_out1 <= in285 XOR in286;

  Logical_Operator_out144_out1 <= in287 XOR in288;

  Logical_Operator_out145_out1 <= in289 XOR in290;

  Logical_Operator_out146_out1 <= in291 XOR in292;

  Logical_Operator_out147_out1 <= in293 XOR in294;

  Logical_Operator_out148_out1 <= in295 XOR in296;

  Logical_Operator_out149_out1 <= in297 XOR in298;

  Logical_Operator_out150_out1 <= in299 XOR in300;

  Logical_Operator_out151_out1 <= in301 XOR in302;

  Logical_Operator_out152_out1 <= in303 XOR in304;

  Logical_Operator_out153_out1 <= in305 XOR in306;

  Logical_Operator_out154_out1 <= in307 XOR in308;

  Logical_Operator_out155_out1 <= in309 XOR in310;

  Logical_Operator_out156_out1 <= in311 XOR in312;

  Logical_Operator_out157_out1 <= in313 XOR in314;

  Logical_Operator_out158_out1 <= in315 XOR in316;

  Logical_Operator_out159_out1 <= in317 XOR in318;

  Logical_Operator_out160_out1 <= in319 XOR in320;

  Logical_Operator_out161_out1 <= in321 XOR in322;

  Logical_Operator_out162_out1 <= in323 XOR in324;

  Logical_Operator_out163_out1 <= in325 XOR in326;

  Logical_Operator_out164_out1 <= in327 XOR in328;

  Logical_Operator_out165_out1 <= in329 XOR in330;

  Logical_Operator_out166_out1 <= in331 XOR in332;

  Logical_Operator_out167_out1 <= in333 XOR in334;

  Logical_Operator_out168_out1 <= in335 XOR in336;

  Logical_Operator_out169_out1 <= in337 XOR in338;

  Logical_Operator_out170_out1 <= in339 XOR in340;

  Logical_Operator_out171_out1 <= in341 XOR in342;

  Logical_Operator_out172_out1 <= in343 XOR in344;

  Logical_Operator_out173_out1 <= in345 XOR in346;

  Logical_Operator_out174_out1 <= in347 XOR in348;

  Logical_Operator_out175_out1 <= in349 XOR in350;

  Logical_Operator_out176_out1 <= in351 XOR in352;

  Logical_Operator_out177_out1 <= in353 XOR in354;

  Logical_Operator_out178_out1 <= in355 XOR in356;

  Logical_Operator_out179_out1 <= in357 XOR in358;

  Logical_Operator_out180_out1 <= in359 XOR in360;

  Logical_Operator_out181_out1 <= in361 XOR in362;

  Logical_Operator_out182_out1 <= in363 XOR in364;

  Logical_Operator_out183_out1 <= in365 XOR in366;

  Logical_Operator_out184_out1 <= in367 XOR in368;

  Logical_Operator_out185_out1 <= in369 XOR in370;

  Logical_Operator_out186_out1 <= in371 XOR in372;

  Logical_Operator_out187_out1 <= in373 XOR in374;

  Logical_Operator_out188_out1 <= in375 XOR in376;

  Logical_Operator_out189_out1 <= in377 XOR in378;

  Logical_Operator_out190_out1 <= in379 XOR in380;

  Logical_Operator_out191_out1 <= in381 XOR in382;

  Logical_Operator_out192_out1 <= in383 XOR in384;

  Logical_Operator_out193_out1 <= in385 XOR in386;

  Logical_Operator_out194_out1 <= in387 XOR in388;

  Logical_Operator_out195_out1 <= in389 XOR in390;

  Logical_Operator_out196_out1 <= in391 XOR in392;

  Logical_Operator_out197_out1 <= in393 XOR in394;

  Logical_Operator_out198_out1 <= in395 XOR in396;

  Logical_Operator_out199_out1 <= in397 XOR in398;

  Logical_Operator_out200_out1 <= in399 XOR in400;

  Logical_Operator_out201_out1 <= in401 XOR in402;

  Logical_Operator_out202_out1 <= in403 XOR in404;

  Logical_Operator_out203_out1 <= in405 XOR in406;

  Logical_Operator_out204_out1 <= in407 XOR in408;

  Logical_Operator_out205_out1 <= in409 XOR in410;

  Logical_Operator_out206_out1 <= in411 XOR in412;

  Logical_Operator_out207_out1 <= in413 XOR in414;

  Logical_Operator_out208_out1 <= in415 XOR in416;

  Logical_Operator_out209_out1 <= in417 XOR in418;

  Logical_Operator_out210_out1 <= in419 XOR in420;

  Logical_Operator_out211_out1 <= in421 XOR in422;

  Logical_Operator_out212_out1 <= in423 XOR in424;

  Logical_Operator_out213_out1 <= in425 XOR in426;

  Logical_Operator_out214_out1 <= in427 XOR in428;

  Logical_Operator_out215_out1 <= in429 XOR in430;

  Logical_Operator_out216_out1 <= in431 XOR in432;

  Logical_Operator_out217_out1 <= in433 XOR in434;

  Logical_Operator_out218_out1 <= in435 XOR in436;

  Logical_Operator_out219_out1 <= in437 XOR in438;

  Logical_Operator_out220_out1 <= in439 XOR in440;

  Logical_Operator_out221_out1 <= in441 XOR in442;

  Logical_Operator_out222_out1 <= in443 XOR in444;

  Logical_Operator_out223_out1 <= in445 XOR in446;

  Logical_Operator_out224_out1 <= in447 XOR in448;

  Logical_Operator_out225_out1 <= in449 XOR in450;

  Logical_Operator_out226_out1 <= in451 XOR in452;

  Logical_Operator_out227_out1 <= in453 XOR in454;

  Logical_Operator_out228_out1 <= in455 XOR in456;

  Logical_Operator_out229_out1 <= in457 XOR in458;

  Logical_Operator_out230_out1 <= in459 XOR in460;

  Logical_Operator_out231_out1 <= in461 XOR in462;

  Logical_Operator_out232_out1 <= in463 XOR in464;

  Logical_Operator_out233_out1 <= in465 XOR in466;

  Logical_Operator_out234_out1 <= in467 XOR in468;

  Logical_Operator_out235_out1 <= in469 XOR in470;

  Logical_Operator_out236_out1 <= in471 XOR in472;

  Logical_Operator_out237_out1 <= in473 XOR in474;

  Logical_Operator_out238_out1 <= in475 XOR in476;

  Logical_Operator_out239_out1 <= in477 XOR in478;

  Logical_Operator_out240_out1 <= in479 XOR in480;

  Logical_Operator_out241_out1 <= in481 XOR in482;

  Logical_Operator_out242_out1 <= in483 XOR in484;

  Logical_Operator_out243_out1 <= in485 XOR in486;

  Logical_Operator_out244_out1 <= in487 XOR in488;

  Logical_Operator_out245_out1 <= in489 XOR in490;

  Logical_Operator_out246_out1 <= in491 XOR in492;

  Logical_Operator_out247_out1 <= in493 XOR in494;

  Logical_Operator_out248_out1 <= in495 XOR in496;

  Logical_Operator_out249_out1 <= in497 XOR in498;

  Logical_Operator_out250_out1 <= in499 XOR in500;

  Logical_Operator_out251_out1 <= in501 XOR in502;

  Logical_Operator_out252_out1 <= in503 XOR in504;

  Logical_Operator_out253_out1 <= in505 XOR in506;

  Logical_Operator_out254_out1 <= in507 XOR in508;

  Logical_Operator_out255_out1 <= in509 XOR in510;

  Logical_Operator_out256_out1 <= in511 XOR in512;

  Logical_Operator_out257_out1 <= in513 XOR in514;

  Logical_Operator_out258_out1 <= in515 XOR in516;

  Logical_Operator_out259_out1 <= in517 XOR in518;

  Logical_Operator_out260_out1 <= in519 XOR in520;

  Logical_Operator_out261_out1 <= in521 XOR in522;

  Logical_Operator_out262_out1 <= in523 XOR in524;

  Logical_Operator_out263_out1 <= in525 XOR in526;

  Logical_Operator_out264_out1 <= in527 XOR in528;

  Logical_Operator_out265_out1 <= in529 XOR in530;

  Logical_Operator_out266_out1 <= in531 XOR in532;

  Logical_Operator_out267_out1 <= in533 XOR in534;

  Logical_Operator_out268_out1 <= in535 XOR in536;

  Logical_Operator_out269_out1 <= in537 XOR in538;

  Logical_Operator_out270_out1 <= in539 XOR in540;

  Logical_Operator_out271_out1 <= in541 XOR in542;

  Logical_Operator_out272_out1 <= in543 XOR in544;

  Logical_Operator_out273_out1 <= in545 XOR in546;

  Logical_Operator_out274_out1 <= in547 XOR in548;

  Logical_Operator_out275_out1 <= in549 XOR in550;

  Logical_Operator_out276_out1 <= in551 XOR in552;

  Logical_Operator_out277_out1 <= in553 XOR in554;

  Logical_Operator_out278_out1 <= in555 XOR in556;

  Logical_Operator_out279_out1 <= in557 XOR in558;

  Logical_Operator_out280_out1 <= in559 XOR in560;

  Logical_Operator_out281_out1 <= in561 XOR in562;

  Logical_Operator_out282_out1 <= in563 XOR in564;

  Logical_Operator_out283_out1 <= in565 XOR in566;

  Logical_Operator_out284_out1 <= in567 XOR in568;

  Logical_Operator_out285_out1 <= in569 XOR in570;

  Logical_Operator_out286_out1 <= in571 XOR in572;

  Logical_Operator_out287_out1 <= in573 XOR in574;

  Logical_Operator_out288_out1 <= in575 XOR in576;

  Logical_Operator_out289_out1 <= in577 XOR in578;

  Logical_Operator_out290_out1 <= in579 XOR in580;

  Logical_Operator_out291_out1 <= in581 XOR in582;

  Logical_Operator_out292_out1 <= in583 XOR in584;

  Logical_Operator_out293_out1 <= in585 XOR in586;

  Logical_Operator_out294_out1 <= in587 XOR in588;

  Logical_Operator_out295_out1 <= in589 XOR in590;

  Logical_Operator_out296_out1 <= in591 XOR in592;

  Logical_Operator_out297_out1 <= in593 XOR in594;

  Logical_Operator_out298_out1 <= in595 XOR in596;

  Logical_Operator_out299_out1 <= in597 XOR in598;

  Logical_Operator_out300_out1 <= in599 XOR in600;

  Logical_Operator_out301_out1 <= in601 XOR in602;

  Logical_Operator_out302_out1 <= in603 XOR in604;

  Logical_Operator_out303_out1 <= in605 XOR in606;

  Logical_Operator_out304_out1 <= in607 XOR in608;

  Logical_Operator_out305_out1 <= in609 XOR in610;

  Logical_Operator_out306_out1 <= in611 XOR in612;

  Logical_Operator_out307_out1 <= in613 XOR in614;

  Logical_Operator_out308_out1 <= in615 XOR in616;

  Logical_Operator_out309_out1 <= in617 XOR in618;

  Logical_Operator_out310_out1 <= in619 XOR in620;

  Logical_Operator_out311_out1 <= in621 XOR in622;

  Logical_Operator_out312_out1 <= in623 XOR in624;

  Logical_Operator_out313_out1 <= in625 XOR in626;

  Logical_Operator_out314_out1 <= in627 XOR in628;

  Logical_Operator_out315_out1 <= in629 XOR in630;

  Logical_Operator_out316_out1 <= in631 XOR in632;

  Logical_Operator_out317_out1 <= in633 XOR in634;

  Logical_Operator_out318_out1 <= in635 XOR in636;

  Logical_Operator_out319_out1 <= in637 XOR in638;

  Logical_Operator_out320_out1 <= in639 XOR in640;

  Logical_Operator_out321_out1 <= in641 XOR in642;

  Logical_Operator_out322_out1 <= in643 XOR in644;

  Logical_Operator_out323_out1 <= in645 XOR in646;

  Logical_Operator_out324_out1 <= in647 XOR in648;

  Logical_Operator_out325_out1 <= in649 XOR in650;

  Logical_Operator_out326_out1 <= in651 XOR in652;

  Logical_Operator_out327_out1 <= in653 XOR in654;

  Logical_Operator_out328_out1 <= in655 XOR in656;

  Logical_Operator_out329_out1 <= in657 XOR in658;

  Logical_Operator_out330_out1 <= in659 XOR in660;

  Logical_Operator_out331_out1 <= in661 XOR in662;

  Logical_Operator_out332_out1 <= in663 XOR in664;

  Logical_Operator_out333_out1 <= in665 XOR in666;

  Logical_Operator_out334_out1 <= in667 XOR in668;

  Logical_Operator_out335_out1 <= in669 XOR in670;

  Logical_Operator_out336_out1 <= in671 XOR in672;

  Logical_Operator_out337_out1 <= in673 XOR in674;

  Logical_Operator_out338_out1 <= in675 XOR in676;

  Logical_Operator_out339_out1 <= in677 XOR in678;

  Logical_Operator_out340_out1 <= in679 XOR in680;

  Logical_Operator_out341_out1 <= in681 XOR in682;

  Logical_Operator_out342_out1 <= in683 XOR in684;

  Logical_Operator_out343_out1 <= in685 XOR in686;

  Logical_Operator_out344_out1 <= in687 XOR in688;

  Logical_Operator_out345_out1 <= in689 XOR in690;

  Logical_Operator_out346_out1 <= in691 XOR in692;

  Logical_Operator_out347_out1 <= in693 XOR in694;

  Logical_Operator_out348_out1 <= in695 XOR in696;

  Logical_Operator_out349_out1 <= in697 XOR in698;

  Logical_Operator_out350_out1 <= in699 XOR in700;

  Logical_Operator_out351_out1 <= in701 XOR in702;

  Logical_Operator_out352_out1 <= in703 XOR in704;

  Logical_Operator_out353_out1 <= in705 XOR in706;

  Logical_Operator_out354_out1 <= in707 XOR in708;

  Logical_Operator_out355_out1 <= in709 XOR in710;

  Logical_Operator_out356_out1 <= in711 XOR in712;

  Logical_Operator_out357_out1 <= in713 XOR in714;

  Logical_Operator_out358_out1 <= in715 XOR in716;

  Logical_Operator_out359_out1 <= in717 XOR in718;

  Logical_Operator_out360_out1 <= in719 XOR in720;

  Logical_Operator_out361_out1 <= in721 XOR in722;

  Logical_Operator_out362_out1 <= in723 XOR in724;

  Logical_Operator_out363_out1 <= in725 XOR in726;

  Logical_Operator_out364_out1 <= in727 XOR in728;

  Logical_Operator_out365_out1 <= in729 XOR in730;

  Logical_Operator_out366_out1 <= in731 XOR in732;

  Logical_Operator_out367_out1 <= in733 XOR in734;

  Logical_Operator_out368_out1 <= in735 XOR in736;

  Logical_Operator_out369_out1 <= in737 XOR in738;

  Logical_Operator_out370_out1 <= in739 XOR in740;

  Logical_Operator_out371_out1 <= in741 XOR in742;

  Logical_Operator_out372_out1 <= in743 XOR in744;

  Logical_Operator_out373_out1 <= in745 XOR in746;

  Logical_Operator_out374_out1 <= in747 XOR in748;

  Logical_Operator_out375_out1 <= in749 XOR in750;

  Logical_Operator_out376_out1 <= in751 XOR in752;

  Logical_Operator_out377_out1 <= in753 XOR in754;

  Logical_Operator_out378_out1 <= in755 XOR in756;

  Logical_Operator_out379_out1 <= in757 XOR in758;

  Logical_Operator_out380_out1 <= in759 XOR in760;

  Logical_Operator_out381_out1 <= in761 XOR in762;

  Logical_Operator_out382_out1 <= in763 XOR in764;

  Logical_Operator_out383_out1 <= in765 XOR in766;

  Logical_Operator_out384_out1 <= in767 XOR in768;

  Logical_Operator_out385_out1 <= in769 XOR in770;

  Logical_Operator_out386_out1 <= in771 XOR in772;

  Logical_Operator_out387_out1 <= in773 XOR in774;

  Logical_Operator_out388_out1 <= in775 XOR in776;

  Logical_Operator_out389_out1 <= in777 XOR in778;

  Logical_Operator_out390_out1 <= in779 XOR in780;

  Logical_Operator_out391_out1 <= in781 XOR in782;

  Logical_Operator_out392_out1 <= in783 XOR in784;

  Logical_Operator_out393_out1 <= in785 XOR in786;

  Logical_Operator_out394_out1 <= in787 XOR in788;

  Logical_Operator_out395_out1 <= in789 XOR in790;

  Logical_Operator_out396_out1 <= in791 XOR in792;

  Logical_Operator_out397_out1 <= in793 XOR in794;

  Logical_Operator_out398_out1 <= in795 XOR in796;

  Logical_Operator_out399_out1 <= in797 XOR in798;

  Logical_Operator_out400_out1 <= in799 XOR in800;

  Logical_Operator_out401_out1 <= in801 XOR in802;

  Logical_Operator_out402_out1 <= in803 XOR in804;

  Logical_Operator_out403_out1 <= in805 XOR in806;

  Logical_Operator_out404_out1 <= in807 XOR in808;

  Logical_Operator_out405_out1 <= in809 XOR in810;

  Logical_Operator_out406_out1 <= in811 XOR in812;

  Logical_Operator_out407_out1 <= in813 XOR in814;

  Logical_Operator_out408_out1 <= in815 XOR in816;

  Logical_Operator_out409_out1 <= in817 XOR in818;

  Logical_Operator_out410_out1 <= in819 XOR in820;

  Logical_Operator_out411_out1 <= in821 XOR in822;

  Logical_Operator_out412_out1 <= in823 XOR in824;

  Logical_Operator_out413_out1 <= in825 XOR in826;

  Logical_Operator_out414_out1 <= in827 XOR in828;

  Logical_Operator_out415_out1 <= in829 XOR in830;

  Logical_Operator_out416_out1 <= in831 XOR in832;

  Logical_Operator_out417_out1 <= in833 XOR in834;

  Logical_Operator_out418_out1 <= in835 XOR in836;

  Logical_Operator_out419_out1 <= in837 XOR in838;

  Logical_Operator_out420_out1 <= in839 XOR in840;

  Logical_Operator_out421_out1 <= in841 XOR in842;

  Logical_Operator_out422_out1 <= in843 XOR in844;

  Logical_Operator_out423_out1 <= in845 XOR in846;

  Logical_Operator_out424_out1 <= in847 XOR in848;

  Logical_Operator_out425_out1 <= in849 XOR in850;

  Logical_Operator_out426_out1 <= in851 XOR in852;

  Logical_Operator_out427_out1 <= in853 XOR in854;

  Logical_Operator_out428_out1 <= in855 XOR in856;

  Logical_Operator_out429_out1 <= in857 XOR in858;

  Logical_Operator_out430_out1 <= in859 XOR in860;

  Logical_Operator_out431_out1 <= in861 XOR in862;

  Logical_Operator_out432_out1 <= in863 XOR in864;

  Logical_Operator_out433_out1 <= in865 XOR in866;

  Logical_Operator_out434_out1 <= in867 XOR in868;

  Logical_Operator_out435_out1 <= in869 XOR in870;

  Logical_Operator_out436_out1 <= in871 XOR in872;

  Logical_Operator_out437_out1 <= in873 XOR in874;

  Logical_Operator_out438_out1 <= in875 XOR in876;

  Logical_Operator_out439_out1 <= in877 XOR in878;

  Logical_Operator_out440_out1 <= in879 XOR in880;

  Logical_Operator_out441_out1 <= in881 XOR in882;

  Logical_Operator_out442_out1 <= in883 XOR in884;

  Logical_Operator_out443_out1 <= in885 XOR in886;

  Logical_Operator_out444_out1 <= in887 XOR in888;

  Logical_Operator_out445_out1 <= in889 XOR in890;

  Logical_Operator_out446_out1 <= in891 XOR in892;

  Logical_Operator_out447_out1 <= in893 XOR in894;

  Logical_Operator_out448_out1 <= in895 XOR in896;

  Logical_Operator_out449_out1 <= in897 XOR in898;

  Logical_Operator_out450_out1 <= in899 XOR in900;

  Logical_Operator_out451_out1 <= in901 XOR in902;

  Logical_Operator_out452_out1 <= in903 XOR in904;

  Logical_Operator_out453_out1 <= in905 XOR in906;

  Logical_Operator_out454_out1 <= in907 XOR in908;

  Logical_Operator_out455_out1 <= in909 XOR in910;

  Logical_Operator_out456_out1 <= in911 XOR in912;

  Logical_Operator_out457_out1 <= in913 XOR in914;

  Logical_Operator_out458_out1 <= in915 XOR in916;

  Logical_Operator_out459_out1 <= in917 XOR in918;

  Logical_Operator_out460_out1 <= in919 XOR in920;

  Logical_Operator_out461_out1 <= in921 XOR in922;

  Logical_Operator_out462_out1 <= in923 XOR in924;

  Logical_Operator_out463_out1 <= in925 XOR in926;

  Logical_Operator_out464_out1 <= in927 XOR in928;

  Logical_Operator_out465_out1 <= in929 XOR in930;

  Logical_Operator_out466_out1 <= in931 XOR in932;

  Logical_Operator_out467_out1 <= in933 XOR in934;

  Logical_Operator_out468_out1 <= in935 XOR in936;

  Logical_Operator_out469_out1 <= in937 XOR in938;

  Logical_Operator_out470_out1 <= in939 XOR in940;

  Logical_Operator_out471_out1 <= in941 XOR in942;

  Logical_Operator_out472_out1 <= in943 XOR in944;

  Logical_Operator_out473_out1 <= in945 XOR in946;

  Logical_Operator_out474_out1 <= in947 XOR in948;

  Logical_Operator_out475_out1 <= in949 XOR in950;

  Logical_Operator_out476_out1 <= in951 XOR in952;

  Logical_Operator_out477_out1 <= in953 XOR in954;

  Logical_Operator_out478_out1 <= in955 XOR in956;

  Logical_Operator_out479_out1 <= in957 XOR in958;

  Logical_Operator_out480_out1 <= in959 XOR in960;

  Logical_Operator_out481_out1 <= in961 XOR in962;

  Logical_Operator_out482_out1 <= in963 XOR in964;

  Logical_Operator_out483_out1 <= in965 XOR in966;

  Logical_Operator_out484_out1 <= in967 XOR in968;

  Logical_Operator_out485_out1 <= in969 XOR in970;

  Logical_Operator_out486_out1 <= in971 XOR in972;

  Logical_Operator_out487_out1 <= in973 XOR in974;

  Logical_Operator_out488_out1 <= in975 XOR in976;

  Logical_Operator_out489_out1 <= in977 XOR in978;

  Logical_Operator_out490_out1 <= in979 XOR in980;

  Logical_Operator_out491_out1 <= in981 XOR in982;

  Logical_Operator_out492_out1 <= in983 XOR in984;

  Logical_Operator_out493_out1 <= in985 XOR in986;

  Logical_Operator_out494_out1 <= in987 XOR in988;

  Logical_Operator_out495_out1 <= in989 XOR in990;

  Logical_Operator_out496_out1 <= in991 XOR in992;

  Logical_Operator_out497_out1 <= in993 XOR in994;

  Logical_Operator_out498_out1 <= in995 XOR in996;

  Logical_Operator_out499_out1 <= in997 XOR in998;

  Logical_Operator_out500_out1 <= in999 XOR in1000;

  Logical_Operator_out501_out1 <= in1001 XOR in1002;

  Logical_Operator_out502_out1 <= in1003 XOR in1004;

  Logical_Operator_out503_out1 <= in1005 XOR in1006;

  Logical_Operator_out504_out1 <= in1007 XOR in1008;

  Logical_Operator_out505_out1 <= in1009 XOR in1010;

  Logical_Operator_out506_out1 <= in1011 XOR in1012;

  Logical_Operator_out507_out1 <= in1013 XOR in1014;

  Logical_Operator_out508_out1 <= in1015 XOR in1016;

  Logical_Operator_out509_out1 <= in1017 XOR in1018;

  Logical_Operator_out510_out1 <= in1019 XOR in1020;

  Logical_Operator_out511_out1 <= in1021 XOR in1022;

  Logical_Operator_out512_out1 <= in1023 XOR in1024;

  Logical_Operator_out513_out1 <= in1025 XOR in1026;

  Logical_Operator_out514_out1 <= in1027 XOR in1028;

  Logical_Operator_out515_out1 <= in1029 XOR in1030;

  Logical_Operator_out516_out1 <= in1031 XOR in1032;

  Logical_Operator_out517_out1 <= in1033 XOR in1034;

  Logical_Operator_out518_out1 <= in1035 XOR in1036;

  Logical_Operator_out519_out1 <= in1037 XOR in1038;

  Logical_Operator_out520_out1 <= in1039 XOR in1040;

  Logical_Operator_out521_out1 <= in1041 XOR in1042;

  Logical_Operator_out522_out1 <= in1043 XOR in1044;

  Logical_Operator_out523_out1 <= in1045 XOR in1046;

  Logical_Operator_out524_out1 <= in1047 XOR in1048;

  Logical_Operator_out525_out1 <= in1049 XOR in1050;

  Logical_Operator_out526_out1 <= in1051 XOR in1052;

  Logical_Operator_out527_out1 <= in1053 XOR in1054;

  Logical_Operator_out528_out1 <= in1055 XOR in1056;

  Logical_Operator_out529_out1 <= in1057 XOR in1058;

  Logical_Operator_out530_out1 <= in1059 XOR in1060;

  Logical_Operator_out531_out1 <= in1061 XOR in1062;

  Logical_Operator_out532_out1 <= in1063 XOR in1064;

  Logical_Operator_out533_out1 <= in1065 XOR in1066;

  Logical_Operator_out534_out1 <= in1067 XOR in1068;

  Logical_Operator_out535_out1 <= in1069 XOR in1070;

  Logical_Operator_out536_out1 <= in1071 XOR in1072;

  Logical_Operator_out537_out1 <= in1073 XOR in1074;

  Logical_Operator_out538_out1 <= in1075 XOR in1076;

  Logical_Operator_out539_out1 <= in1077 XOR in1078;

  Logical_Operator_out540_out1 <= in1079 XOR in1080;

  Logical_Operator_out541_out1 <= in1081 XOR in1082;

  Logical_Operator_out542_out1 <= in1083 XOR in1084;

  Logical_Operator_out543_out1 <= in1085 XOR in1086;

  Logical_Operator_out544_out1 <= in1087 XOR in1088;

  Logical_Operator_out545_out1 <= in1089 XOR in1090;

  Logical_Operator_out546_out1 <= in1091 XOR in1092;

  Logical_Operator_out547_out1 <= in1093 XOR in1094;

  Logical_Operator_out548_out1 <= in1095 XOR in1096;

  Logical_Operator_out549_out1 <= in1097 XOR in1098;

  Logical_Operator_out550_out1 <= in1099 XOR in1100;

  Logical_Operator_out551_out1 <= in1101 XOR in1102;

  Logical_Operator_out552_out1 <= in1103 XOR in1104;

  Logical_Operator_out553_out1 <= in1105 XOR in1106;

  Logical_Operator_out554_out1 <= in1107 XOR in1108;

  Logical_Operator_out555_out1 <= in1109 XOR in1110;

  Logical_Operator_out556_out1 <= in1111 XOR in1112;

  Logical_Operator_out557_out1 <= in1113 XOR in1114;

  Logical_Operator_out558_out1 <= in1115 XOR in1116;

  Logical_Operator_out559_out1 <= in1117 XOR in1118;

  Logical_Operator_out560_out1 <= in1119 XOR in1120;

  Logical_Operator_out561_out1 <= in1121 XOR in1122;

  Logical_Operator_out562_out1 <= in1123 XOR in1124;

  Logical_Operator_out563_out1 <= in1125 XOR in1126;

  Logical_Operator_out564_out1 <= in1127 XOR in1128;

  Logical_Operator_out565_out1 <= in1129 XOR in1130;

  Logical_Operator_out566_out1 <= in1131 XOR in1132;

  Logical_Operator_out567_out1 <= in1133 XOR in1134;

  Logical_Operator_out568_out1 <= in1135 XOR in1136;

  Logical_Operator_out569_out1 <= in1137 XOR in1138;

  Logical_Operator_out570_out1 <= in1139 XOR in1140;

  Logical_Operator_out571_out1 <= in1141 XOR in1142;

  Logical_Operator_out572_out1 <= in1143 XOR in1144;

  Logical_Operator_out573_out1 <= in1145 XOR in1146;

  Logical_Operator_out574_out1 <= in1147 XOR in1148;

  Logical_Operator_out575_out1 <= in1149 XOR in1150;

  Logical_Operator_out576_out1 <= in1151 XOR in1152;

  Logical_Operator_out577_out1 <= in1153 XOR in1154;

  Logical_Operator_out578_out1 <= in1155 XOR in1156;

  Logical_Operator_out579_out1 <= in1157 XOR in1158;

  Logical_Operator_out580_out1 <= in1159 XOR in1160;

  Logical_Operator_out581_out1 <= in1161 XOR in1162;

  Logical_Operator_out582_out1 <= in1163 XOR in1164;

  Logical_Operator_out583_out1 <= in1165 XOR in1166;

  Logical_Operator_out584_out1 <= in1167 XOR in1168;

  Logical_Operator_out585_out1 <= in1169 XOR in1170;

  Logical_Operator_out586_out1 <= in1171 XOR in1172;

  Logical_Operator_out587_out1 <= in1173 XOR in1174;

  Logical_Operator_out588_out1 <= in1175 XOR in1176;

  Logical_Operator_out589_out1 <= in1177 XOR in1178;

  Logical_Operator_out590_out1 <= in1179 XOR in1180;

  Logical_Operator_out591_out1 <= in1181 XOR in1182;

  Logical_Operator_out592_out1 <= in1183 XOR in1184;

  Logical_Operator_out593_out1 <= in1185 XOR in1186;

  Logical_Operator_out594_out1 <= in1187 XOR in1188;

  Logical_Operator_out595_out1 <= in1189 XOR in1190;

  Logical_Operator_out596_out1 <= in1191 XOR in1192;

  Logical_Operator_out597_out1 <= in1193 XOR in1194;

  Logical_Operator_out598_out1 <= in1195 XOR in1196;

  Logical_Operator_out599_out1 <= in1197 XOR in1198;

  Logical_Operator_out600_out1 <= in1199 XOR in1200;

  Logical_Operator_out601_out1 <= in1201 XOR in1202;

  Logical_Operator_out602_out1 <= in1203 XOR in1204;

  Logical_Operator_out603_out1 <= in1205 XOR in1206;

  Logical_Operator_out604_out1 <= in1207 XOR in1208;

  Logical_Operator_out605_out1 <= in1209 XOR in1210;

  Logical_Operator_out606_out1 <= in1211 XOR in1212;

  Logical_Operator_out607_out1 <= in1213 XOR in1214;

  Logical_Operator_out608_out1 <= in1215 XOR in1216;

  Logical_Operator_out609_out1 <= in1217 XOR in1218;

  Logical_Operator_out610_out1 <= in1219 XOR in1220;

  Logical_Operator_out611_out1 <= in1221 XOR in1222;

  Logical_Operator_out612_out1 <= in1223 XOR in1224;

  Logical_Operator_out613_out1 <= in1225 XOR in1226;

  Logical_Operator_out614_out1 <= in1227 XOR in1228;

  Logical_Operator_out615_out1 <= in1229 XOR in1230;

  Logical_Operator_out616_out1 <= in1231 XOR in1232;

  Logical_Operator_out617_out1 <= in1233 XOR in1234;

  Logical_Operator_out618_out1 <= in1235 XOR in1236;

  Logical_Operator_out619_out1 <= in1237 XOR in1238;

  Logical_Operator_out620_out1 <= in1239 XOR in1240;

  Logical_Operator_out621_out1 <= in1241 XOR in1242;

  Logical_Operator_out622_out1 <= in1243 XOR in1244;

  Logical_Operator_out623_out1 <= in1245 XOR in1246;

  Logical_Operator_out624_out1 <= in1247 XOR in1248;

  Logical_Operator_out625_out1 <= in1249 XOR in1250;

  Logical_Operator_out626_out1 <= in1251 XOR in1252;

  Logical_Operator_out627_out1 <= in1253 XOR in1254;

  Logical_Operator_out628_out1 <= in1255 XOR in1256;

  Logical_Operator_out629_out1 <= in1257 XOR in1258;

  Logical_Operator_out630_out1 <= in1259 XOR in1260;

  Logical_Operator_out631_out1 <= in1261 XOR in1262;

  Logical_Operator_out632_out1 <= in1263 XOR in1264;

  Logical_Operator_out633_out1 <= in1265 XOR in1266;

  Logical_Operator_out634_out1 <= in1267 XOR in1268;

  Logical_Operator_out635_out1 <= in1269 XOR in1270;

  Logical_Operator_out636_out1 <= in1271 XOR in1272;

  Logical_Operator_out637_out1 <= in1273 XOR in1274;

  Logical_Operator_out638_out1 <= in1275 XOR in1276;

  Logical_Operator_out639_out1 <= in1277 XOR in1278;

  Logical_Operator_out640_out1 <= in1279 XOR in1280;

  Logical_Operator_out641_out1 <= in1281 XOR in1282;

  Logical_Operator_out642_out1 <= in1283 XOR in1284;

  Logical_Operator_out643_out1 <= in1285 XOR in1286;

  Logical_Operator_out644_out1 <= in1287 XOR in1288;

  Logical_Operator_out645_out1 <= in1289 XOR in1290;

  Logical_Operator_out646_out1 <= in1291 XOR in1292;

  Logical_Operator_out647_out1 <= in1293 XOR in1294;

  Logical_Operator_out648_out1 <= in1295 XOR in1296;

  Logical_Operator_out649_out1 <= in1297 XOR in1298;

  Logical_Operator_out650_out1 <= in1299 XOR in1300;

  Logical_Operator_out651_out1 <= in1301 XOR in1302;

  Logical_Operator_out652_out1 <= in1303 XOR in1304;

  Logical_Operator_out653_out1 <= in1305 XOR in1306;

  Logical_Operator_out654_out1 <= in1307 XOR in1308;

  Logical_Operator_out655_out1 <= in1309 XOR in1310;

  Logical_Operator_out656_out1 <= in1311 XOR in1312;

  Logical_Operator_out657_out1 <= in1313 XOR in1314;

  Logical_Operator_out658_out1 <= in1315 XOR in1316;

  Logical_Operator_out659_out1 <= in1317 XOR in1318;

  Logical_Operator_out660_out1 <= in1319 XOR in1320;

  Logical_Operator_out661_out1 <= in1321 XOR in1322;

  Logical_Operator_out662_out1 <= in1323 XOR in1324;

  Logical_Operator_out663_out1 <= in1325 XOR in1326;

  Logical_Operator_out664_out1 <= in1327 XOR in1328;

  Logical_Operator_out665_out1 <= in1329 XOR in1330;

  Logical_Operator_out666_out1 <= in1331 XOR in1332;

  Logical_Operator_out667_out1 <= in1333 XOR in1334;

  Logical_Operator_out668_out1 <= in1335 XOR in1336;

  Logical_Operator_out669_out1 <= in1337 XOR in1338;

  Logical_Operator_out670_out1 <= in1339 XOR in1340;

  Logical_Operator_out671_out1 <= in1341 XOR in1342;

  Logical_Operator_out672_out1 <= in1343 XOR in1344;

  Logical_Operator_out673_out1 <= in1345 XOR in1346;

  Logical_Operator_out674_out1 <= in1347 XOR in1348;

  Logical_Operator_out675_out1 <= in1349 XOR in1350;

  Logical_Operator_out676_out1 <= in1351 XOR in1352;

  Logical_Operator_out677_out1 <= in1353 XOR in1354;

  Logical_Operator_out678_out1 <= in1355 XOR in1356;

  Logical_Operator_out679_out1 <= in1357 XOR in1358;

  Logical_Operator_out680_out1 <= in1359 XOR in1360;

  Logical_Operator_out681_out1 <= in1361 XOR in1362;

  Logical_Operator_out682_out1 <= in1363 XOR in1364;

  Logical_Operator_out683_out1 <= in1365 XOR in1366;

  Logical_Operator_out684_out1 <= in1367 XOR in1368;

  Logical_Operator_out685_out1 <= in1369 XOR in1370;

  Logical_Operator_out686_out1 <= in1371 XOR in1372;

  Logical_Operator_out687_out1 <= in1373 XOR in1374;

  Logical_Operator_out688_out1 <= in1375 XOR in1376;

  Logical_Operator_out689_out1 <= in1377 XOR in1378;

  Logical_Operator_out690_out1 <= in1379 XOR in1380;

  Logical_Operator_out691_out1 <= in1381 XOR in1382;

  Logical_Operator_out692_out1 <= in1383 XOR in1384;

  Logical_Operator_out693_out1 <= in1385 XOR in1386;

  Logical_Operator_out694_out1 <= in1387 XOR in1388;

  Logical_Operator_out695_out1 <= in1389 XOR in1390;

  Logical_Operator_out696_out1 <= in1391 XOR in1392;

  Logical_Operator_out697_out1 <= in1393 XOR in1394;

  Logical_Operator_out698_out1 <= in1395 XOR in1396;

  Logical_Operator_out699_out1 <= in1397 XOR in1398;

  Logical_Operator_out700_out1 <= in1399 XOR in1400;

  Logical_Operator_out701_out1 <= in1401 XOR in1402;

  Logical_Operator_out702_out1 <= in1403 XOR in1404;

  Logical_Operator_out703_out1 <= in1405 XOR in1406;

  Logical_Operator_out704_out1 <= in1407 XOR in1408;

  Logical_Operator_out705_out1 <= in1409 XOR in1410;

  Logical_Operator_out706_out1 <= in1411 XOR in1412;

  Logical_Operator_out707_out1 <= in1413 XOR in1414;

  Logical_Operator_out708_out1 <= in1415 XOR in1416;

  Logical_Operator_out709_out1 <= in1417 XOR in1418;

  Logical_Operator_out710_out1 <= in1419 XOR in1420;

  Logical_Operator_out711_out1 <= in1421 XOR in1422;

  Logical_Operator_out712_out1 <= in1423 XOR in1424;

  Logical_Operator_out713_out1 <= in1425 XOR in1426;

  Logical_Operator_out714_out1 <= in1427 XOR in1428;

  Logical_Operator_out715_out1 <= in1429 XOR in1430;

  Logical_Operator_out716_out1 <= in1431 XOR in1432;

  Logical_Operator_out717_out1 <= in1433 XOR in1434;

  Logical_Operator_out718_out1 <= in1435 XOR in1436;

  Logical_Operator_out719_out1 <= in1437 XOR in1438;

  Logical_Operator_out720_out1 <= in1439 XOR in1440;

  Logical_Operator_out721_out1 <= in1441 XOR in1442;

  Logical_Operator_out722_out1 <= in1443 XOR in1444;

  Logical_Operator_out723_out1 <= in1445 XOR in1446;

  Logical_Operator_out724_out1 <= in1447 XOR in1448;

  Logical_Operator_out725_out1 <= in1449 XOR in1450;

  Logical_Operator_out726_out1 <= in1451 XOR in1452;

  Logical_Operator_out727_out1 <= in1453 XOR in1454;

  Logical_Operator_out728_out1 <= in1455 XOR in1456;

  Logical_Operator_out729_out1 <= in1457 XOR in1458;

  Logical_Operator_out730_out1 <= in1459 XOR in1460;

  Logical_Operator_out731_out1 <= in1461 XOR in1462;

  Logical_Operator_out732_out1 <= in1463 XOR in1464;

  Logical_Operator_out733_out1 <= in1465 XOR in1466;

  Logical_Operator_out734_out1 <= in1467 XOR in1468;

  Logical_Operator_out735_out1 <= in1469 XOR in1470;

  Logical_Operator_out736_out1 <= in1471 XOR in1472;

  Logical_Operator_out737_out1 <= in1473 XOR in1474;

  Logical_Operator_out738_out1 <= in1475 XOR in1476;

  Logical_Operator_out739_out1 <= in1477 XOR in1478;

  Logical_Operator_out740_out1 <= in1479 XOR in1480;

  Logical_Operator_out741_out1 <= in1481 XOR in1482;

  Logical_Operator_out742_out1 <= in1483 XOR in1484;

  Logical_Operator_out743_out1 <= in1485 XOR in1486;

  Logical_Operator_out744_out1 <= in1487 XOR in1488;

  Logical_Operator_out745_out1 <= in1489 XOR in1490;

  Logical_Operator_out746_out1 <= in1491 XOR in1492;

  Logical_Operator_out747_out1 <= in1493 XOR in1494;

  Logical_Operator_out748_out1 <= in1495 XOR in1496;

  Logical_Operator_out749_out1 <= in1497 XOR in1498;

  Logical_Operator_out750_out1 <= in1499 XOR in1500;

  Logical_Operator_out751_out1 <= in1501 XOR in1502;

  Logical_Operator_out752_out1 <= in1503 XOR in1504;

  Logical_Operator_out753_out1 <= in1505 XOR in1506;

  Logical_Operator_out754_out1 <= in1507 XOR in1508;

  Logical_Operator_out755_out1 <= in1509 XOR in1510;

  Logical_Operator_out756_out1 <= in1511 XOR in1512;

  Logical_Operator_out757_out1 <= in1513 XOR in1514;

  Logical_Operator_out758_out1 <= in1515 XOR in1516;

  Logical_Operator_out759_out1 <= in1517 XOR in1518;

  Logical_Operator_out760_out1 <= in1519 XOR in1520;

  Logical_Operator_out761_out1 <= in1521 XOR in1522;

  Logical_Operator_out762_out1 <= in1523 XOR in1524;

  Logical_Operator_out763_out1 <= in1525 XOR in1526;

  Logical_Operator_out764_out1 <= in1527 XOR in1528;

  Logical_Operator_out765_out1 <= in1529 XOR in1530;

  Logical_Operator_out766_out1 <= in1531 XOR in1532;

  Logical_Operator_out767_out1 <= in1533 XOR in1534;

  Logical_Operator_out768_out1 <= in1535 XOR in1536;

  Logical_Operator_out769_out1 <= in1537 XOR in1538;

  Logical_Operator_out770_out1 <= in1539 XOR in1540;

  Logical_Operator_out771_out1 <= in1541 XOR in1542;

  Logical_Operator_out772_out1 <= in1543 XOR in1544;

  Logical_Operator_out773_out1 <= in1545 XOR in1546;

  Logical_Operator_out774_out1 <= in1547 XOR in1548;

  Logical_Operator_out775_out1 <= in1549 XOR in1550;

  Logical_Operator_out776_out1 <= in1551 XOR in1552;

  Logical_Operator_out777_out1 <= in1553 XOR in1554;

  Logical_Operator_out778_out1 <= in1555 XOR in1556;

  Logical_Operator_out779_out1 <= in1557 XOR in1558;

  Logical_Operator_out780_out1 <= in1559 XOR in1560;

  Logical_Operator_out781_out1 <= in1561 XOR in1562;

  Logical_Operator_out782_out1 <= in1563 XOR in1564;

  Logical_Operator_out783_out1 <= in1565 XOR in1566;

  Logical_Operator_out784_out1 <= in1567 XOR in1568;

  Logical_Operator_out785_out1 <= in1569 XOR in1570;

  Logical_Operator_out786_out1 <= in1571 XOR in1572;

  Logical_Operator_out787_out1 <= in1573 XOR in1574;

  Logical_Operator_out788_out1 <= in1575 XOR in1576;

  Logical_Operator_out789_out1 <= in1577 XOR in1578;

  Logical_Operator_out790_out1 <= in1579 XOR in1580;

  Logical_Operator_out791_out1 <= in1581 XOR in1582;

  Logical_Operator_out792_out1 <= in1583 XOR in1584;

  Logical_Operator_out793_out1 <= in1585 XOR in1586;

  Logical_Operator_out794_out1 <= in1587 XOR in1588;

  Logical_Operator_out795_out1 <= in1589 XOR in1590;

  Logical_Operator_out796_out1 <= in1591 XOR in1592;

  Logical_Operator_out797_out1 <= in1593 XOR in1594;

  Logical_Operator_out798_out1 <= in1595 XOR in1596;

  Logical_Operator_out799_out1 <= in1597 XOR in1598;

  Logical_Operator_out800_out1 <= in1599 XOR in1600;

  Logical_Operator_out801_out1 <= in1601 XOR in1602;

  Logical_Operator_out802_out1 <= in1603 XOR in1604;

  Logical_Operator_out803_out1 <= in1605 XOR in1606;

  Logical_Operator_out804_out1 <= in1607 XOR in1608;

  Logical_Operator_out805_out1 <= in1609 XOR in1610;

  Logical_Operator_out806_out1 <= in1611 XOR in1612;

  Logical_Operator_out807_out1 <= in1613 XOR in1614;

  Logical_Operator_out808_out1 <= in1615 XOR in1616;

  Logical_Operator_out809_out1 <= in1617 XOR in1618;

  Logical_Operator_out810_out1 <= in1619 XOR in1620;

  Logical_Operator_out811_out1 <= in1621 XOR in1622;

  Logical_Operator_out812_out1 <= in1623 XOR in1624;

  Logical_Operator_out813_out1 <= in1625 XOR in1626;

  Logical_Operator_out814_out1 <= in1627 XOR in1628;

  Logical_Operator_out815_out1 <= in1629 XOR in1630;

  Logical_Operator_out816_out1 <= in1631 XOR in1632;

  Logical_Operator_out817_out1 <= in1633 XOR in1634;

  Logical_Operator_out818_out1 <= in1635 XOR in1636;

  Logical_Operator_out819_out1 <= in1637 XOR in1638;

  Logical_Operator_out820_out1 <= in1639 XOR in1640;

  Logical_Operator_out821_out1 <= in1641 XOR in1642;

  Logical_Operator_out822_out1 <= in1643 XOR in1644;

  Logical_Operator_out823_out1 <= in1645 XOR in1646;

  Logical_Operator_out824_out1 <= in1647 XOR in1648;

  Logical_Operator_out825_out1 <= in1649 XOR in1650;

  Logical_Operator_out826_out1 <= in1651 XOR in1652;

  Logical_Operator_out827_out1 <= in1653 XOR in1654;

  Logical_Operator_out828_out1 <= in1655 XOR in1656;

  Logical_Operator_out829_out1 <= in1657 XOR in1658;

  Logical_Operator_out830_out1 <= in1659 XOR in1660;

  Logical_Operator_out831_out1 <= in1661 XOR in1662;

  Logical_Operator_out832_out1 <= in1663 XOR in1664;

  Logical_Operator_out833_out1 <= in1665 XOR in1666;

  Logical_Operator_out834_out1 <= in1667 XOR in1668;

  Logical_Operator_out835_out1 <= in1669 XOR in1670;

  Logical_Operator_out836_out1 <= in1671 XOR in1672;

  Logical_Operator_out837_out1 <= in1673 XOR in1674;

  Logical_Operator_out838_out1 <= in1675 XOR in1676;

  Logical_Operator_out839_out1 <= in1677 XOR in1678;

  Logical_Operator_out840_out1 <= in1679 XOR in1680;

  Logical_Operator_out841_out1 <= in1681 XOR in1682;

  Logical_Operator_out842_out1 <= in1683 XOR in1684;

  Logical_Operator_out843_out1 <= in1685 XOR in1686;

  Logical_Operator_out844_out1 <= in1687 XOR in1688;

  Logical_Operator_out845_out1 <= in1689 XOR in1690;

  Logical_Operator_out846_out1 <= in1691 XOR in1692;

  Logical_Operator_out847_out1 <= in1693 XOR in1694;

  Logical_Operator_out848_out1 <= in1695 XOR in1696;

  Logical_Operator_out849_out1 <= in1697 XOR in1698;

  Logical_Operator_out850_out1 <= in1699 XOR in1700;

  Logical_Operator_out851_out1 <= in1701 XOR in1702;

  Logical_Operator_out852_out1 <= in1703 XOR in1704;

  Logical_Operator_out853_out1 <= in1705 XOR in1706;

  Logical_Operator_out854_out1 <= in1707 XOR in1708;

  Logical_Operator_out855_out1 <= in1709 XOR in1710;

  Logical_Operator_out856_out1 <= in1711 XOR in1712;

  Logical_Operator_out857_out1 <= in1713 XOR in1714;

  Logical_Operator_out858_out1 <= in1715 XOR in1716;

  Logical_Operator_out859_out1 <= in1717 XOR in1718;

  Logical_Operator_out860_out1 <= in1719 XOR in1720;

  Logical_Operator_out861_out1 <= in1721 XOR in1722;

  Logical_Operator_out862_out1 <= in1723 XOR in1724;

  Logical_Operator_out863_out1 <= in1725 XOR in1726;

  Logical_Operator_out864_out1 <= in1727 XOR in1728;

  Logical_Operator_out865_out1 <= in1729 XOR in1730;

  Logical_Operator_out866_out1 <= in1731 XOR in1732;

  Logical_Operator_out867_out1 <= in1733 XOR in1734;

  Logical_Operator_out868_out1 <= in1735 XOR in1736;

  Logical_Operator_out869_out1 <= in1737 XOR in1738;

  Logical_Operator_out870_out1 <= in1739 XOR in1740;

  Logical_Operator_out871_out1 <= in1741 XOR in1742;

  Logical_Operator_out872_out1 <= in1743 XOR in1744;

  Logical_Operator_out873_out1 <= in1745 XOR in1746;

  Logical_Operator_out874_out1 <= in1747 XOR in1748;

  Logical_Operator_out875_out1 <= in1749 XOR in1750;

  Logical_Operator_out876_out1 <= in1751 XOR in1752;

  Logical_Operator_out877_out1 <= in1753 XOR in1754;

  Logical_Operator_out878_out1 <= in1755 XOR in1756;

  Logical_Operator_out879_out1 <= in1757 XOR in1758;

  Logical_Operator_out880_out1 <= in1759 XOR in1760;

  Logical_Operator_out881_out1 <= in1761 XOR in1762;

  Logical_Operator_out882_out1 <= in1763 XOR in1764;

  Logical_Operator_out883_out1 <= in1765 XOR in1766;

  Logical_Operator_out884_out1 <= in1767 XOR in1768;

  Logical_Operator_out885_out1 <= in1769 XOR in1770;

  Logical_Operator_out886_out1 <= in1771 XOR in1772;

  Logical_Operator_out887_out1 <= in1773 XOR in1774;

  Logical_Operator_out888_out1 <= in1775 XOR in1776;

  Logical_Operator_out889_out1 <= in1777 XOR in1778;

  Logical_Operator_out890_out1 <= in1779 XOR in1780;

  Logical_Operator_out891_out1 <= in1781 XOR in1782;

  Logical_Operator_out892_out1 <= in1783 XOR in1784;

  Logical_Operator_out893_out1 <= in1785 XOR in1786;

  Logical_Operator_out894_out1 <= in1787 XOR in1788;

  Logical_Operator_out895_out1 <= in1789 XOR in1790;

  Logical_Operator_out896_out1 <= in1791 XOR in1792;

  Logical_Operator_out897_out1 <= in1793 XOR in1794;

  Logical_Operator_out898_out1 <= in1795 XOR in1796;

  Logical_Operator_out899_out1 <= in1797 XOR in1798;

  Logical_Operator_out900_out1 <= in1799 XOR in1800;

  Logical_Operator_out901_out1 <= in1801 XOR in1802;

  Logical_Operator_out902_out1 <= in1803 XOR in1804;

  Logical_Operator_out903_out1 <= in1805 XOR in1806;

  Logical_Operator_out904_out1 <= in1807 XOR in1808;

  Logical_Operator_out905_out1 <= in1809 XOR in1810;

  Logical_Operator_out906_out1 <= in1811 XOR in1812;

  Logical_Operator_out907_out1 <= in1813 XOR in1814;

  Logical_Operator_out908_out1 <= in1815 XOR in1816;

  Logical_Operator_out909_out1 <= in1817 XOR in1818;

  Logical_Operator_out910_out1 <= in1819 XOR in1820;

  Logical_Operator_out911_out1 <= in1821 XOR in1822;

  Logical_Operator_out912_out1 <= in1823 XOR in1824;

  Logical_Operator_out913_out1 <= in1825 XOR in1826;

  Logical_Operator_out914_out1 <= in1827 XOR in1828;

  Logical_Operator_out915_out1 <= in1829 XOR in1830;

  Logical_Operator_out916_out1 <= in1831 XOR in1832;

  Logical_Operator_out917_out1 <= in1833 XOR in1834;

  Logical_Operator_out918_out1 <= in1835 XOR in1836;

  Logical_Operator_out919_out1 <= in1837 XOR in1838;

  Logical_Operator_out920_out1 <= in1839 XOR in1840;

  Logical_Operator_out921_out1 <= in1841 XOR in1842;

  Logical_Operator_out922_out1 <= in1843 XOR in1844;

  Logical_Operator_out923_out1 <= in1845 XOR in1846;

  Logical_Operator_out924_out1 <= in1847 XOR in1848;

  Logical_Operator_out925_out1 <= in1849 XOR in1850;

  Logical_Operator_out926_out1 <= in1851 XOR in1852;

  Logical_Operator_out927_out1 <= in1853 XOR in1854;

  Logical_Operator_out928_out1 <= in1855 XOR in1856;

  Logical_Operator_out929_out1 <= in1857 XOR in1858;

  Logical_Operator_out930_out1 <= in1859 XOR in1860;

  Logical_Operator_out931_out1 <= in1861 XOR in1862;

  Logical_Operator_out932_out1 <= in1863 XOR in1864;

  Logical_Operator_out933_out1 <= in1865 XOR in1866;

  Logical_Operator_out934_out1 <= in1867 XOR in1868;

  Logical_Operator_out935_out1 <= in1869 XOR in1870;

  Logical_Operator_out936_out1 <= in1871 XOR in1872;

  Logical_Operator_out937_out1 <= in1873 XOR in1874;

  Logical_Operator_out938_out1 <= in1875 XOR in1876;

  Logical_Operator_out939_out1 <= in1877 XOR in1878;

  Logical_Operator_out940_out1 <= in1879 XOR in1880;

  Logical_Operator_out941_out1 <= in1881 XOR in1882;

  Logical_Operator_out942_out1 <= in1883 XOR in1884;

  Logical_Operator_out943_out1 <= in1885 XOR in1886;

  Logical_Operator_out944_out1 <= in1887 XOR in1888;

  Logical_Operator_out945_out1 <= in1889 XOR in1890;

  Logical_Operator_out946_out1 <= in1891 XOR in1892;

  Logical_Operator_out947_out1 <= in1893 XOR in1894;

  Logical_Operator_out948_out1 <= in1895 XOR in1896;

  Logical_Operator_out949_out1 <= in1897 XOR in1898;

  Logical_Operator_out950_out1 <= in1899 XOR in1900;

  Logical_Operator_out951_out1 <= in1901 XOR in1902;

  Logical_Operator_out952_out1 <= in1903 XOR in1904;

  Logical_Operator_out953_out1 <= in1905 XOR in1906;

  Logical_Operator_out954_out1 <= in1907 XOR in1908;

  Logical_Operator_out955_out1 <= in1909 XOR in1910;

  Logical_Operator_out956_out1 <= in1911 XOR in1912;

  Logical_Operator_out957_out1 <= in1913 XOR in1914;

  Logical_Operator_out958_out1 <= in1915 XOR in1916;

  Logical_Operator_out959_out1 <= in1917 XOR in1918;

  Logical_Operator_out960_out1 <= in1919 XOR in1920;

  Logical_Operator_out961_out1 <= in1921 XOR in1922;

  Logical_Operator_out962_out1 <= in1923 XOR in1924;

  Logical_Operator_out963_out1 <= in1925 XOR in1926;

  Logical_Operator_out964_out1 <= in1927 XOR in1928;

  Logical_Operator_out965_out1 <= in1929 XOR in1930;

  Logical_Operator_out966_out1 <= in1931 XOR in1932;

  Logical_Operator_out967_out1 <= in1933 XOR in1934;

  Logical_Operator_out968_out1 <= in1935 XOR in1936;

  Logical_Operator_out969_out1 <= in1937 XOR in1938;

  Logical_Operator_out970_out1 <= in1939 XOR in1940;

  Logical_Operator_out971_out1 <= in1941 XOR in1942;

  Logical_Operator_out972_out1 <= in1943 XOR in1944;

  Logical_Operator_out973_out1 <= in1945 XOR in1946;

  Logical_Operator_out974_out1 <= in1947 XOR in1948;

  Logical_Operator_out975_out1 <= in1949 XOR in1950;

  Logical_Operator_out976_out1 <= in1951 XOR in1952;

  Logical_Operator_out977_out1 <= in1953 XOR in1954;

  Logical_Operator_out978_out1 <= in1955 XOR in1956;

  Logical_Operator_out979_out1 <= in1957 XOR in1958;

  Logical_Operator_out980_out1 <= in1959 XOR in1960;

  Logical_Operator_out981_out1 <= in1961 XOR in1962;

  Logical_Operator_out982_out1 <= in1963 XOR in1964;

  Logical_Operator_out983_out1 <= in1965 XOR in1966;

  Logical_Operator_out984_out1 <= in1967 XOR in1968;

  Logical_Operator_out985_out1 <= in1969 XOR in1970;

  Logical_Operator_out986_out1 <= in1971 XOR in1972;

  Logical_Operator_out987_out1 <= in1973 XOR in1974;

  Logical_Operator_out988_out1 <= in1975 XOR in1976;

  Logical_Operator_out989_out1 <= in1977 XOR in1978;

  Logical_Operator_out990_out1 <= in1979 XOR in1980;

  Logical_Operator_out991_out1 <= in1981 XOR in1982;

  Logical_Operator_out992_out1 <= in1983 XOR in1984;

  Logical_Operator_out993_out1 <= in1985 XOR in1986;

  Logical_Operator_out994_out1 <= in1987 XOR in1988;

  Logical_Operator_out995_out1 <= in1989 XOR in1990;

  Logical_Operator_out996_out1 <= in1991 XOR in1992;

  Logical_Operator_out997_out1 <= in1993 XOR in1994;

  Logical_Operator_out998_out1 <= in1995 XOR in1996;

  Logical_Operator_out999_out1 <= in1997 XOR in1998;

  Logical_Operator_out1000_out1 <= in1999 XOR in2000;

  Logical_Operator_out1001_out1 <= in2001 XOR in2002;

  Logical_Operator_out1002_out1 <= in2003 XOR in2004;

  Logical_Operator_out1003_out1 <= in2005 XOR in2006;

  Logical_Operator_out1004_out1 <= in2007 XOR in2008;

  Logical_Operator_out1005_out1 <= in2009 XOR in2010;

  Logical_Operator_out1006_out1 <= in2011 XOR in2012;

  Logical_Operator_out1007_out1 <= in2013 XOR in2014;

  Logical_Operator_out1008_out1 <= in2015 XOR in2016;

  Logical_Operator_out1009_out1 <= in2017 XOR in2018;

  Logical_Operator_out1010_out1 <= in2019 XOR in2020;

  Logical_Operator_out1011_out1 <= in2021 XOR in2022;

  Logical_Operator_out1012_out1 <= in2023 XOR in2024;

  Logical_Operator_out1013_out1 <= in2025 XOR in2026;

  Logical_Operator_out1014_out1 <= in2027 XOR in2028;

  Logical_Operator_out1015_out1 <= in2029 XOR in2030;

  Logical_Operator_out1016_out1 <= in2031 XOR in2032;

  Logical_Operator_out1017_out1 <= in2033 XOR in2034;

  Logical_Operator_out1018_out1 <= in2035 XOR in2036;

  Logical_Operator_out1019_out1 <= in2037 XOR in2038;

  Logical_Operator_out1020_out1 <= in2039 XOR in2040;

  Logical_Operator_out1021_out1 <= in2041 XOR in2042;

  Logical_Operator_out1022_out1 <= in2043 XOR in2044;

  Logical_Operator_out1023_out1 <= in2045 XOR in2046;

  Logical_Operator_out1024_out1 <= in2047 XOR in2048;

  Logical_Operator_out1025_out1 <= Logical_Operator_out1_out1 XOR Logical_Operator_out2_out1;

  Logical_Operator_out1026_out1 <= in2 XOR in4;

  Logical_Operator_out1027_out1 <= Logical_Operator_out3_out1 XOR Logical_Operator_out4_out1;

  Logical_Operator_out1028_out1 <= in6 XOR in8;

  Logical_Operator_out1029_out1 <= Logical_Operator_out5_out1 XOR Logical_Operator_out6_out1;

  Logical_Operator_out1030_out1 <= in10 XOR in12;

  Logical_Operator_out1031_out1 <= Logical_Operator_out7_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out1032_out1 <= in14 XOR in16;

  Logical_Operator_out1033_out1 <= Logical_Operator_out9_out1 XOR Logical_Operator_out10_out1;

  Logical_Operator_out1034_out1 <= in18 XOR in20;

  Logical_Operator_out1035_out1 <= Logical_Operator_out11_out1 XOR Logical_Operator_out12_out1;

  Logical_Operator_out1036_out1 <= in22 XOR in24;

  Logical_Operator_out1037_out1 <= Logical_Operator_out13_out1 XOR Logical_Operator_out14_out1;

  Logical_Operator_out1038_out1 <= in26 XOR in28;

  Logical_Operator_out1039_out1 <= Logical_Operator_out15_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out1040_out1 <= in30 XOR in32;

  Logical_Operator_out1041_out1 <= Logical_Operator_out17_out1 XOR Logical_Operator_out18_out1;

  Logical_Operator_out1042_out1 <= in34 XOR in36;

  Logical_Operator_out1043_out1 <= Logical_Operator_out19_out1 XOR Logical_Operator_out20_out1;

  Logical_Operator_out1044_out1 <= in38 XOR in40;

  Logical_Operator_out1045_out1 <= Logical_Operator_out21_out1 XOR Logical_Operator_out22_out1;

  Logical_Operator_out1046_out1 <= in42 XOR in44;

  Logical_Operator_out1047_out1 <= Logical_Operator_out23_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out1048_out1 <= in46 XOR in48;

  Logical_Operator_out1049_out1 <= Logical_Operator_out25_out1 XOR Logical_Operator_out26_out1;

  Logical_Operator_out1050_out1 <= in50 XOR in52;

  Logical_Operator_out1051_out1 <= Logical_Operator_out27_out1 XOR Logical_Operator_out28_out1;

  Logical_Operator_out1052_out1 <= in54 XOR in56;

  Logical_Operator_out1053_out1 <= Logical_Operator_out29_out1 XOR Logical_Operator_out30_out1;

  Logical_Operator_out1054_out1 <= in58 XOR in60;

  Logical_Operator_out1055_out1 <= Logical_Operator_out31_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out1056_out1 <= in62 XOR in64;

  Logical_Operator_out1057_out1 <= Logical_Operator_out33_out1 XOR Logical_Operator_out34_out1;

  Logical_Operator_out1058_out1 <= in66 XOR in68;

  Logical_Operator_out1059_out1 <= Logical_Operator_out35_out1 XOR Logical_Operator_out36_out1;

  Logical_Operator_out1060_out1 <= in70 XOR in72;

  Logical_Operator_out1061_out1 <= Logical_Operator_out37_out1 XOR Logical_Operator_out38_out1;

  Logical_Operator_out1062_out1 <= in74 XOR in76;

  Logical_Operator_out1063_out1 <= Logical_Operator_out39_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out1064_out1 <= in78 XOR in80;

  Logical_Operator_out1065_out1 <= Logical_Operator_out41_out1 XOR Logical_Operator_out42_out1;

  Logical_Operator_out1066_out1 <= in82 XOR in84;

  Logical_Operator_out1067_out1 <= Logical_Operator_out43_out1 XOR Logical_Operator_out44_out1;

  Logical_Operator_out1068_out1 <= in86 XOR in88;

  Logical_Operator_out1069_out1 <= Logical_Operator_out45_out1 XOR Logical_Operator_out46_out1;

  Logical_Operator_out1070_out1 <= in90 XOR in92;

  Logical_Operator_out1071_out1 <= Logical_Operator_out47_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out1072_out1 <= in94 XOR in96;

  Logical_Operator_out1073_out1 <= Logical_Operator_out49_out1 XOR Logical_Operator_out50_out1;

  Logical_Operator_out1074_out1 <= in98 XOR in100;

  Logical_Operator_out1075_out1 <= Logical_Operator_out51_out1 XOR Logical_Operator_out52_out1;

  Logical_Operator_out1076_out1 <= in102 XOR in104;

  Logical_Operator_out1077_out1 <= Logical_Operator_out53_out1 XOR Logical_Operator_out54_out1;

  Logical_Operator_out1078_out1 <= in106 XOR in108;

  Logical_Operator_out1079_out1 <= Logical_Operator_out55_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out1080_out1 <= in110 XOR in112;

  Logical_Operator_out1081_out1 <= Logical_Operator_out57_out1 XOR Logical_Operator_out58_out1;

  Logical_Operator_out1082_out1 <= in114 XOR in116;

  Logical_Operator_out1083_out1 <= Logical_Operator_out59_out1 XOR Logical_Operator_out60_out1;

  Logical_Operator_out1084_out1 <= in118 XOR in120;

  Logical_Operator_out1085_out1 <= Logical_Operator_out61_out1 XOR Logical_Operator_out62_out1;

  Logical_Operator_out1086_out1 <= in122 XOR in124;

  Logical_Operator_out1087_out1 <= Logical_Operator_out63_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out1088_out1 <= in126 XOR in128;

  Logical_Operator_out1089_out1 <= Logical_Operator_out65_out1 XOR Logical_Operator_out66_out1;

  Logical_Operator_out1090_out1 <= in130 XOR in132;

  Logical_Operator_out1091_out1 <= Logical_Operator_out67_out1 XOR Logical_Operator_out68_out1;

  Logical_Operator_out1092_out1 <= in134 XOR in136;

  Logical_Operator_out1093_out1 <= Logical_Operator_out69_out1 XOR Logical_Operator_out70_out1;

  Logical_Operator_out1094_out1 <= in138 XOR in140;

  Logical_Operator_out1095_out1 <= Logical_Operator_out71_out1 XOR Logical_Operator_out72_out1;

  Logical_Operator_out1096_out1 <= in142 XOR in144;

  Logical_Operator_out1097_out1 <= Logical_Operator_out73_out1 XOR Logical_Operator_out74_out1;

  Logical_Operator_out1098_out1 <= in146 XOR in148;

  Logical_Operator_out1099_out1 <= Logical_Operator_out75_out1 XOR Logical_Operator_out76_out1;

  Logical_Operator_out1100_out1 <= in150 XOR in152;

  Logical_Operator_out1101_out1 <= Logical_Operator_out77_out1 XOR Logical_Operator_out78_out1;

  Logical_Operator_out1102_out1 <= in154 XOR in156;

  Logical_Operator_out1103_out1 <= Logical_Operator_out79_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out1104_out1 <= in158 XOR in160;

  Logical_Operator_out1105_out1 <= Logical_Operator_out81_out1 XOR Logical_Operator_out82_out1;

  Logical_Operator_out1106_out1 <= in162 XOR in164;

  Logical_Operator_out1107_out1 <= Logical_Operator_out83_out1 XOR Logical_Operator_out84_out1;

  Logical_Operator_out1108_out1 <= in166 XOR in168;

  Logical_Operator_out1109_out1 <= Logical_Operator_out85_out1 XOR Logical_Operator_out86_out1;

  Logical_Operator_out1110_out1 <= in170 XOR in172;

  Logical_Operator_out1111_out1 <= Logical_Operator_out87_out1 XOR Logical_Operator_out88_out1;

  Logical_Operator_out1112_out1 <= in174 XOR in176;

  Logical_Operator_out1113_out1 <= Logical_Operator_out89_out1 XOR Logical_Operator_out90_out1;

  Logical_Operator_out1114_out1 <= in178 XOR in180;

  Logical_Operator_out1115_out1 <= Logical_Operator_out91_out1 XOR Logical_Operator_out92_out1;

  Logical_Operator_out1116_out1 <= in182 XOR in184;

  Logical_Operator_out1117_out1 <= Logical_Operator_out93_out1 XOR Logical_Operator_out94_out1;

  Logical_Operator_out1118_out1 <= in186 XOR in188;

  Logical_Operator_out1119_out1 <= Logical_Operator_out95_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out1120_out1 <= in190 XOR in192;

  Logical_Operator_out1121_out1 <= Logical_Operator_out97_out1 XOR Logical_Operator_out98_out1;

  Logical_Operator_out1122_out1 <= in194 XOR in196;

  Logical_Operator_out1123_out1 <= Logical_Operator_out99_out1 XOR Logical_Operator_out100_out1;

  Logical_Operator_out1124_out1 <= in198 XOR in200;

  Logical_Operator_out1125_out1 <= Logical_Operator_out101_out1 XOR Logical_Operator_out102_out1;

  Logical_Operator_out1126_out1 <= in202 XOR in204;

  Logical_Operator_out1127_out1 <= Logical_Operator_out103_out1 XOR Logical_Operator_out104_out1;

  Logical_Operator_out1128_out1 <= in206 XOR in208;

  Logical_Operator_out1129_out1 <= Logical_Operator_out105_out1 XOR Logical_Operator_out106_out1;

  Logical_Operator_out1130_out1 <= in210 XOR in212;

  Logical_Operator_out1131_out1 <= Logical_Operator_out107_out1 XOR Logical_Operator_out108_out1;

  Logical_Operator_out1132_out1 <= in214 XOR in216;

  Logical_Operator_out1133_out1 <= Logical_Operator_out109_out1 XOR Logical_Operator_out110_out1;

  Logical_Operator_out1134_out1 <= in218 XOR in220;

  Logical_Operator_out1135_out1 <= Logical_Operator_out111_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out1136_out1 <= in222 XOR in224;

  Logical_Operator_out1137_out1 <= Logical_Operator_out113_out1 XOR Logical_Operator_out114_out1;

  Logical_Operator_out1138_out1 <= in226 XOR in228;

  Logical_Operator_out1139_out1 <= Logical_Operator_out115_out1 XOR Logical_Operator_out116_out1;

  Logical_Operator_out1140_out1 <= in230 XOR in232;

  Logical_Operator_out1141_out1 <= Logical_Operator_out117_out1 XOR Logical_Operator_out118_out1;

  Logical_Operator_out1142_out1 <= in234 XOR in236;

  Logical_Operator_out1143_out1 <= Logical_Operator_out119_out1 XOR Logical_Operator_out120_out1;

  Logical_Operator_out1144_out1 <= in238 XOR in240;

  Logical_Operator_out1145_out1 <= Logical_Operator_out121_out1 XOR Logical_Operator_out122_out1;

  Logical_Operator_out1146_out1 <= in242 XOR in244;

  Logical_Operator_out1147_out1 <= Logical_Operator_out123_out1 XOR Logical_Operator_out124_out1;

  Logical_Operator_out1148_out1 <= in246 XOR in248;

  Logical_Operator_out1149_out1 <= Logical_Operator_out125_out1 XOR Logical_Operator_out126_out1;

  Logical_Operator_out1150_out1 <= in250 XOR in252;

  Logical_Operator_out1151_out1 <= Logical_Operator_out127_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out1152_out1 <= in254 XOR in256;

  Logical_Operator_out1153_out1 <= Logical_Operator_out129_out1 XOR Logical_Operator_out130_out1;

  Logical_Operator_out1154_out1 <= in258 XOR in260;

  Logical_Operator_out1155_out1 <= Logical_Operator_out131_out1 XOR Logical_Operator_out132_out1;

  Logical_Operator_out1156_out1 <= in262 XOR in264;

  Logical_Operator_out1157_out1 <= Logical_Operator_out133_out1 XOR Logical_Operator_out134_out1;

  Logical_Operator_out1158_out1 <= in266 XOR in268;

  Logical_Operator_out1159_out1 <= Logical_Operator_out135_out1 XOR Logical_Operator_out136_out1;

  Logical_Operator_out1160_out1 <= in270 XOR in272;

  Logical_Operator_out1161_out1 <= Logical_Operator_out137_out1 XOR Logical_Operator_out138_out1;

  Logical_Operator_out1162_out1 <= in274 XOR in276;

  Logical_Operator_out1163_out1 <= Logical_Operator_out139_out1 XOR Logical_Operator_out140_out1;

  Logical_Operator_out1164_out1 <= in278 XOR in280;

  Logical_Operator_out1165_out1 <= Logical_Operator_out141_out1 XOR Logical_Operator_out142_out1;

  Logical_Operator_out1166_out1 <= in282 XOR in284;

  Logical_Operator_out1167_out1 <= Logical_Operator_out143_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out1168_out1 <= in286 XOR in288;

  Logical_Operator_out1169_out1 <= Logical_Operator_out145_out1 XOR Logical_Operator_out146_out1;

  Logical_Operator_out1170_out1 <= in290 XOR in292;

  Logical_Operator_out1171_out1 <= Logical_Operator_out147_out1 XOR Logical_Operator_out148_out1;

  Logical_Operator_out1172_out1 <= in294 XOR in296;

  Logical_Operator_out1173_out1 <= Logical_Operator_out149_out1 XOR Logical_Operator_out150_out1;

  Logical_Operator_out1174_out1 <= in298 XOR in300;

  Logical_Operator_out1175_out1 <= Logical_Operator_out151_out1 XOR Logical_Operator_out152_out1;

  Logical_Operator_out1176_out1 <= in302 XOR in304;

  Logical_Operator_out1177_out1 <= Logical_Operator_out153_out1 XOR Logical_Operator_out154_out1;

  Logical_Operator_out1178_out1 <= in306 XOR in308;

  Logical_Operator_out1179_out1 <= Logical_Operator_out155_out1 XOR Logical_Operator_out156_out1;

  Logical_Operator_out1180_out1 <= in310 XOR in312;

  Logical_Operator_out1181_out1 <= Logical_Operator_out157_out1 XOR Logical_Operator_out158_out1;

  Logical_Operator_out1182_out1 <= in314 XOR in316;

  Logical_Operator_out1183_out1 <= Logical_Operator_out159_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out1184_out1 <= in318 XOR in320;

  Logical_Operator_out1185_out1 <= Logical_Operator_out161_out1 XOR Logical_Operator_out162_out1;

  Logical_Operator_out1186_out1 <= in322 XOR in324;

  Logical_Operator_out1187_out1 <= Logical_Operator_out163_out1 XOR Logical_Operator_out164_out1;

  Logical_Operator_out1188_out1 <= in326 XOR in328;

  Logical_Operator_out1189_out1 <= Logical_Operator_out165_out1 XOR Logical_Operator_out166_out1;

  Logical_Operator_out1190_out1 <= in330 XOR in332;

  Logical_Operator_out1191_out1 <= Logical_Operator_out167_out1 XOR Logical_Operator_out168_out1;

  Logical_Operator_out1192_out1 <= in334 XOR in336;

  Logical_Operator_out1193_out1 <= Logical_Operator_out169_out1 XOR Logical_Operator_out170_out1;

  Logical_Operator_out1194_out1 <= in338 XOR in340;

  Logical_Operator_out1195_out1 <= Logical_Operator_out171_out1 XOR Logical_Operator_out172_out1;

  Logical_Operator_out1196_out1 <= in342 XOR in344;

  Logical_Operator_out1197_out1 <= Logical_Operator_out173_out1 XOR Logical_Operator_out174_out1;

  Logical_Operator_out1198_out1 <= in346 XOR in348;

  Logical_Operator_out1199_out1 <= Logical_Operator_out175_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out1200_out1 <= in350 XOR in352;

  Logical_Operator_out1201_out1 <= Logical_Operator_out177_out1 XOR Logical_Operator_out178_out1;

  Logical_Operator_out1202_out1 <= in354 XOR in356;

  Logical_Operator_out1203_out1 <= Logical_Operator_out179_out1 XOR Logical_Operator_out180_out1;

  Logical_Operator_out1204_out1 <= in358 XOR in360;

  Logical_Operator_out1205_out1 <= Logical_Operator_out181_out1 XOR Logical_Operator_out182_out1;

  Logical_Operator_out1206_out1 <= in362 XOR in364;

  Logical_Operator_out1207_out1 <= Logical_Operator_out183_out1 XOR Logical_Operator_out184_out1;

  Logical_Operator_out1208_out1 <= in366 XOR in368;

  Logical_Operator_out1209_out1 <= Logical_Operator_out185_out1 XOR Logical_Operator_out186_out1;

  Logical_Operator_out1210_out1 <= in370 XOR in372;

  Logical_Operator_out1211_out1 <= Logical_Operator_out187_out1 XOR Logical_Operator_out188_out1;

  Logical_Operator_out1212_out1 <= in374 XOR in376;

  Logical_Operator_out1213_out1 <= Logical_Operator_out189_out1 XOR Logical_Operator_out190_out1;

  Logical_Operator_out1214_out1 <= in378 XOR in380;

  Logical_Operator_out1215_out1 <= Logical_Operator_out191_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out1216_out1 <= in382 XOR in384;

  Logical_Operator_out1217_out1 <= Logical_Operator_out193_out1 XOR Logical_Operator_out194_out1;

  Logical_Operator_out1218_out1 <= in386 XOR in388;

  Logical_Operator_out1219_out1 <= Logical_Operator_out195_out1 XOR Logical_Operator_out196_out1;

  Logical_Operator_out1220_out1 <= in390 XOR in392;

  Logical_Operator_out1221_out1 <= Logical_Operator_out197_out1 XOR Logical_Operator_out198_out1;

  Logical_Operator_out1222_out1 <= in394 XOR in396;

  Logical_Operator_out1223_out1 <= Logical_Operator_out199_out1 XOR Logical_Operator_out200_out1;

  Logical_Operator_out1224_out1 <= in398 XOR in400;

  Logical_Operator_out1225_out1 <= Logical_Operator_out201_out1 XOR Logical_Operator_out202_out1;

  Logical_Operator_out1226_out1 <= in402 XOR in404;

  Logical_Operator_out1227_out1 <= Logical_Operator_out203_out1 XOR Logical_Operator_out204_out1;

  Logical_Operator_out1228_out1 <= in406 XOR in408;

  Logical_Operator_out1229_out1 <= Logical_Operator_out205_out1 XOR Logical_Operator_out206_out1;

  Logical_Operator_out1230_out1 <= in410 XOR in412;

  Logical_Operator_out1231_out1 <= Logical_Operator_out207_out1 XOR Logical_Operator_out208_out1;

  Logical_Operator_out1232_out1 <= in414 XOR in416;

  Logical_Operator_out1233_out1 <= Logical_Operator_out209_out1 XOR Logical_Operator_out210_out1;

  Logical_Operator_out1234_out1 <= in418 XOR in420;

  Logical_Operator_out1235_out1 <= Logical_Operator_out211_out1 XOR Logical_Operator_out212_out1;

  Logical_Operator_out1236_out1 <= in422 XOR in424;

  Logical_Operator_out1237_out1 <= Logical_Operator_out213_out1 XOR Logical_Operator_out214_out1;

  Logical_Operator_out1238_out1 <= in426 XOR in428;

  Logical_Operator_out1239_out1 <= Logical_Operator_out215_out1 XOR Logical_Operator_out216_out1;

  Logical_Operator_out1240_out1 <= in430 XOR in432;

  Logical_Operator_out1241_out1 <= Logical_Operator_out217_out1 XOR Logical_Operator_out218_out1;

  Logical_Operator_out1242_out1 <= in434 XOR in436;

  Logical_Operator_out1243_out1 <= Logical_Operator_out219_out1 XOR Logical_Operator_out220_out1;

  Logical_Operator_out1244_out1 <= in438 XOR in440;

  Logical_Operator_out1245_out1 <= Logical_Operator_out221_out1 XOR Logical_Operator_out222_out1;

  Logical_Operator_out1246_out1 <= in442 XOR in444;

  Logical_Operator_out1247_out1 <= Logical_Operator_out223_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out1248_out1 <= in446 XOR in448;

  Logical_Operator_out1249_out1 <= Logical_Operator_out225_out1 XOR Logical_Operator_out226_out1;

  Logical_Operator_out1250_out1 <= in450 XOR in452;

  Logical_Operator_out1251_out1 <= Logical_Operator_out227_out1 XOR Logical_Operator_out228_out1;

  Logical_Operator_out1252_out1 <= in454 XOR in456;

  Logical_Operator_out1253_out1 <= Logical_Operator_out229_out1 XOR Logical_Operator_out230_out1;

  Logical_Operator_out1254_out1 <= in458 XOR in460;

  Logical_Operator_out1255_out1 <= Logical_Operator_out231_out1 XOR Logical_Operator_out232_out1;

  Logical_Operator_out1256_out1 <= in462 XOR in464;

  Logical_Operator_out1257_out1 <= Logical_Operator_out233_out1 XOR Logical_Operator_out234_out1;

  Logical_Operator_out1258_out1 <= in466 XOR in468;

  Logical_Operator_out1259_out1 <= Logical_Operator_out235_out1 XOR Logical_Operator_out236_out1;

  Logical_Operator_out1260_out1 <= in470 XOR in472;

  Logical_Operator_out1261_out1 <= Logical_Operator_out237_out1 XOR Logical_Operator_out238_out1;

  Logical_Operator_out1262_out1 <= in474 XOR in476;

  Logical_Operator_out1263_out1 <= Logical_Operator_out239_out1 XOR Logical_Operator_out240_out1;

  Logical_Operator_out1264_out1 <= in478 XOR in480;

  Logical_Operator_out1265_out1 <= Logical_Operator_out241_out1 XOR Logical_Operator_out242_out1;

  Logical_Operator_out1266_out1 <= in482 XOR in484;

  Logical_Operator_out1267_out1 <= Logical_Operator_out243_out1 XOR Logical_Operator_out244_out1;

  Logical_Operator_out1268_out1 <= in486 XOR in488;

  Logical_Operator_out1269_out1 <= Logical_Operator_out245_out1 XOR Logical_Operator_out246_out1;

  Logical_Operator_out1270_out1 <= in490 XOR in492;

  Logical_Operator_out1271_out1 <= Logical_Operator_out247_out1 XOR Logical_Operator_out248_out1;

  Logical_Operator_out1272_out1 <= in494 XOR in496;

  Logical_Operator_out1273_out1 <= Logical_Operator_out249_out1 XOR Logical_Operator_out250_out1;

  Logical_Operator_out1274_out1 <= in498 XOR in500;

  Logical_Operator_out1275_out1 <= Logical_Operator_out251_out1 XOR Logical_Operator_out252_out1;

  Logical_Operator_out1276_out1 <= in502 XOR in504;

  Logical_Operator_out1277_out1 <= Logical_Operator_out253_out1 XOR Logical_Operator_out254_out1;

  Logical_Operator_out1278_out1 <= in506 XOR in508;

  Logical_Operator_out1279_out1 <= Logical_Operator_out255_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out1280_out1 <= in510 XOR in512;

  Logical_Operator_out1281_out1 <= Logical_Operator_out257_out1 XOR Logical_Operator_out258_out1;

  Logical_Operator_out1282_out1 <= in514 XOR in516;

  Logical_Operator_out1283_out1 <= Logical_Operator_out259_out1 XOR Logical_Operator_out260_out1;

  Logical_Operator_out1284_out1 <= in518 XOR in520;

  Logical_Operator_out1285_out1 <= Logical_Operator_out261_out1 XOR Logical_Operator_out262_out1;

  Logical_Operator_out1286_out1 <= in522 XOR in524;

  Logical_Operator_out1287_out1 <= Logical_Operator_out263_out1 XOR Logical_Operator_out264_out1;

  Logical_Operator_out1288_out1 <= in526 XOR in528;

  Logical_Operator_out1289_out1 <= Logical_Operator_out265_out1 XOR Logical_Operator_out266_out1;

  Logical_Operator_out1290_out1 <= in530 XOR in532;

  Logical_Operator_out1291_out1 <= Logical_Operator_out267_out1 XOR Logical_Operator_out268_out1;

  Logical_Operator_out1292_out1 <= in534 XOR in536;

  Logical_Operator_out1293_out1 <= Logical_Operator_out269_out1 XOR Logical_Operator_out270_out1;

  Logical_Operator_out1294_out1 <= in538 XOR in540;

  Logical_Operator_out1295_out1 <= Logical_Operator_out271_out1 XOR Logical_Operator_out272_out1;

  Logical_Operator_out1296_out1 <= in542 XOR in544;

  Logical_Operator_out1297_out1 <= Logical_Operator_out273_out1 XOR Logical_Operator_out274_out1;

  Logical_Operator_out1298_out1 <= in546 XOR in548;

  Logical_Operator_out1299_out1 <= Logical_Operator_out275_out1 XOR Logical_Operator_out276_out1;

  Logical_Operator_out1300_out1 <= in550 XOR in552;

  Logical_Operator_out1301_out1 <= Logical_Operator_out277_out1 XOR Logical_Operator_out278_out1;

  Logical_Operator_out1302_out1 <= in554 XOR in556;

  Logical_Operator_out1303_out1 <= Logical_Operator_out279_out1 XOR Logical_Operator_out280_out1;

  Logical_Operator_out1304_out1 <= in558 XOR in560;

  Logical_Operator_out1305_out1 <= Logical_Operator_out281_out1 XOR Logical_Operator_out282_out1;

  Logical_Operator_out1306_out1 <= in562 XOR in564;

  Logical_Operator_out1307_out1 <= Logical_Operator_out283_out1 XOR Logical_Operator_out284_out1;

  Logical_Operator_out1308_out1 <= in566 XOR in568;

  Logical_Operator_out1309_out1 <= Logical_Operator_out285_out1 XOR Logical_Operator_out286_out1;

  Logical_Operator_out1310_out1 <= in570 XOR in572;

  Logical_Operator_out1311_out1 <= Logical_Operator_out287_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out1312_out1 <= in574 XOR in576;

  Logical_Operator_out1313_out1 <= Logical_Operator_out289_out1 XOR Logical_Operator_out290_out1;

  Logical_Operator_out1314_out1 <= in578 XOR in580;

  Logical_Operator_out1315_out1 <= Logical_Operator_out291_out1 XOR Logical_Operator_out292_out1;

  Logical_Operator_out1316_out1 <= in582 XOR in584;

  Logical_Operator_out1317_out1 <= Logical_Operator_out293_out1 XOR Logical_Operator_out294_out1;

  Logical_Operator_out1318_out1 <= in586 XOR in588;

  Logical_Operator_out1319_out1 <= Logical_Operator_out295_out1 XOR Logical_Operator_out296_out1;

  Logical_Operator_out1320_out1 <= in590 XOR in592;

  Logical_Operator_out1321_out1 <= Logical_Operator_out297_out1 XOR Logical_Operator_out298_out1;

  Logical_Operator_out1322_out1 <= in594 XOR in596;

  Logical_Operator_out1323_out1 <= Logical_Operator_out299_out1 XOR Logical_Operator_out300_out1;

  Logical_Operator_out1324_out1 <= in598 XOR in600;

  Logical_Operator_out1325_out1 <= Logical_Operator_out301_out1 XOR Logical_Operator_out302_out1;

  Logical_Operator_out1326_out1 <= in602 XOR in604;

  Logical_Operator_out1327_out1 <= Logical_Operator_out303_out1 XOR Logical_Operator_out304_out1;

  Logical_Operator_out1328_out1 <= in606 XOR in608;

  Logical_Operator_out1329_out1 <= Logical_Operator_out305_out1 XOR Logical_Operator_out306_out1;

  Logical_Operator_out1330_out1 <= in610 XOR in612;

  Logical_Operator_out1331_out1 <= Logical_Operator_out307_out1 XOR Logical_Operator_out308_out1;

  Logical_Operator_out1332_out1 <= in614 XOR in616;

  Logical_Operator_out1333_out1 <= Logical_Operator_out309_out1 XOR Logical_Operator_out310_out1;

  Logical_Operator_out1334_out1 <= in618 XOR in620;

  Logical_Operator_out1335_out1 <= Logical_Operator_out311_out1 XOR Logical_Operator_out312_out1;

  Logical_Operator_out1336_out1 <= in622 XOR in624;

  Logical_Operator_out1337_out1 <= Logical_Operator_out313_out1 XOR Logical_Operator_out314_out1;

  Logical_Operator_out1338_out1 <= in626 XOR in628;

  Logical_Operator_out1339_out1 <= Logical_Operator_out315_out1 XOR Logical_Operator_out316_out1;

  Logical_Operator_out1340_out1 <= in630 XOR in632;

  Logical_Operator_out1341_out1 <= Logical_Operator_out317_out1 XOR Logical_Operator_out318_out1;

  Logical_Operator_out1342_out1 <= in634 XOR in636;

  Logical_Operator_out1343_out1 <= Logical_Operator_out319_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out1344_out1 <= in638 XOR in640;

  Logical_Operator_out1345_out1 <= Logical_Operator_out321_out1 XOR Logical_Operator_out322_out1;

  Logical_Operator_out1346_out1 <= in642 XOR in644;

  Logical_Operator_out1347_out1 <= Logical_Operator_out323_out1 XOR Logical_Operator_out324_out1;

  Logical_Operator_out1348_out1 <= in646 XOR in648;

  Logical_Operator_out1349_out1 <= Logical_Operator_out325_out1 XOR Logical_Operator_out326_out1;

  Logical_Operator_out1350_out1 <= in650 XOR in652;

  Logical_Operator_out1351_out1 <= Logical_Operator_out327_out1 XOR Logical_Operator_out328_out1;

  Logical_Operator_out1352_out1 <= in654 XOR in656;

  Logical_Operator_out1353_out1 <= Logical_Operator_out329_out1 XOR Logical_Operator_out330_out1;

  Logical_Operator_out1354_out1 <= in658 XOR in660;

  Logical_Operator_out1355_out1 <= Logical_Operator_out331_out1 XOR Logical_Operator_out332_out1;

  Logical_Operator_out1356_out1 <= in662 XOR in664;

  Logical_Operator_out1357_out1 <= Logical_Operator_out333_out1 XOR Logical_Operator_out334_out1;

  Logical_Operator_out1358_out1 <= in666 XOR in668;

  Logical_Operator_out1359_out1 <= Logical_Operator_out335_out1 XOR Logical_Operator_out336_out1;

  Logical_Operator_out1360_out1 <= in670 XOR in672;

  Logical_Operator_out1361_out1 <= Logical_Operator_out337_out1 XOR Logical_Operator_out338_out1;

  Logical_Operator_out1362_out1 <= in674 XOR in676;

  Logical_Operator_out1363_out1 <= Logical_Operator_out339_out1 XOR Logical_Operator_out340_out1;

  Logical_Operator_out1364_out1 <= in678 XOR in680;

  Logical_Operator_out1365_out1 <= Logical_Operator_out341_out1 XOR Logical_Operator_out342_out1;

  Logical_Operator_out1366_out1 <= in682 XOR in684;

  Logical_Operator_out1367_out1 <= Logical_Operator_out343_out1 XOR Logical_Operator_out344_out1;

  Logical_Operator_out1368_out1 <= in686 XOR in688;

  Logical_Operator_out1369_out1 <= Logical_Operator_out345_out1 XOR Logical_Operator_out346_out1;

  Logical_Operator_out1370_out1 <= in690 XOR in692;

  Logical_Operator_out1371_out1 <= Logical_Operator_out347_out1 XOR Logical_Operator_out348_out1;

  Logical_Operator_out1372_out1 <= in694 XOR in696;

  Logical_Operator_out1373_out1 <= Logical_Operator_out349_out1 XOR Logical_Operator_out350_out1;

  Logical_Operator_out1374_out1 <= in698 XOR in700;

  Logical_Operator_out1375_out1 <= Logical_Operator_out351_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out1376_out1 <= in702 XOR in704;

  Logical_Operator_out1377_out1 <= Logical_Operator_out353_out1 XOR Logical_Operator_out354_out1;

  Logical_Operator_out1378_out1 <= in706 XOR in708;

  Logical_Operator_out1379_out1 <= Logical_Operator_out355_out1 XOR Logical_Operator_out356_out1;

  Logical_Operator_out1380_out1 <= in710 XOR in712;

  Logical_Operator_out1381_out1 <= Logical_Operator_out357_out1 XOR Logical_Operator_out358_out1;

  Logical_Operator_out1382_out1 <= in714 XOR in716;

  Logical_Operator_out1383_out1 <= Logical_Operator_out359_out1 XOR Logical_Operator_out360_out1;

  Logical_Operator_out1384_out1 <= in718 XOR in720;

  Logical_Operator_out1385_out1 <= Logical_Operator_out361_out1 XOR Logical_Operator_out362_out1;

  Logical_Operator_out1386_out1 <= in722 XOR in724;

  Logical_Operator_out1387_out1 <= Logical_Operator_out363_out1 XOR Logical_Operator_out364_out1;

  Logical_Operator_out1388_out1 <= in726 XOR in728;

  Logical_Operator_out1389_out1 <= Logical_Operator_out365_out1 XOR Logical_Operator_out366_out1;

  Logical_Operator_out1390_out1 <= in730 XOR in732;

  Logical_Operator_out1391_out1 <= Logical_Operator_out367_out1 XOR Logical_Operator_out368_out1;

  Logical_Operator_out1392_out1 <= in734 XOR in736;

  Logical_Operator_out1393_out1 <= Logical_Operator_out369_out1 XOR Logical_Operator_out370_out1;

  Logical_Operator_out1394_out1 <= in738 XOR in740;

  Logical_Operator_out1395_out1 <= Logical_Operator_out371_out1 XOR Logical_Operator_out372_out1;

  Logical_Operator_out1396_out1 <= in742 XOR in744;

  Logical_Operator_out1397_out1 <= Logical_Operator_out373_out1 XOR Logical_Operator_out374_out1;

  Logical_Operator_out1398_out1 <= in746 XOR in748;

  Logical_Operator_out1399_out1 <= Logical_Operator_out375_out1 XOR Logical_Operator_out376_out1;

  Logical_Operator_out1400_out1 <= in750 XOR in752;

  Logical_Operator_out1401_out1 <= Logical_Operator_out377_out1 XOR Logical_Operator_out378_out1;

  Logical_Operator_out1402_out1 <= in754 XOR in756;

  Logical_Operator_out1403_out1 <= Logical_Operator_out379_out1 XOR Logical_Operator_out380_out1;

  Logical_Operator_out1404_out1 <= in758 XOR in760;

  Logical_Operator_out1405_out1 <= Logical_Operator_out381_out1 XOR Logical_Operator_out382_out1;

  Logical_Operator_out1406_out1 <= in762 XOR in764;

  Logical_Operator_out1407_out1 <= Logical_Operator_out383_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out1408_out1 <= in766 XOR in768;

  Logical_Operator_out1409_out1 <= Logical_Operator_out385_out1 XOR Logical_Operator_out386_out1;

  Logical_Operator_out1410_out1 <= in770 XOR in772;

  Logical_Operator_out1411_out1 <= Logical_Operator_out387_out1 XOR Logical_Operator_out388_out1;

  Logical_Operator_out1412_out1 <= in774 XOR in776;

  Logical_Operator_out1413_out1 <= Logical_Operator_out389_out1 XOR Logical_Operator_out390_out1;

  Logical_Operator_out1414_out1 <= in778 XOR in780;

  Logical_Operator_out1415_out1 <= Logical_Operator_out391_out1 XOR Logical_Operator_out392_out1;

  Logical_Operator_out1416_out1 <= in782 XOR in784;

  Logical_Operator_out1417_out1 <= Logical_Operator_out393_out1 XOR Logical_Operator_out394_out1;

  Logical_Operator_out1418_out1 <= in786 XOR in788;

  Logical_Operator_out1419_out1 <= Logical_Operator_out395_out1 XOR Logical_Operator_out396_out1;

  Logical_Operator_out1420_out1 <= in790 XOR in792;

  Logical_Operator_out1421_out1 <= Logical_Operator_out397_out1 XOR Logical_Operator_out398_out1;

  Logical_Operator_out1422_out1 <= in794 XOR in796;

  Logical_Operator_out1423_out1 <= Logical_Operator_out399_out1 XOR Logical_Operator_out400_out1;

  Logical_Operator_out1424_out1 <= in798 XOR in800;

  Logical_Operator_out1425_out1 <= Logical_Operator_out401_out1 XOR Logical_Operator_out402_out1;

  Logical_Operator_out1426_out1 <= in802 XOR in804;

  Logical_Operator_out1427_out1 <= Logical_Operator_out403_out1 XOR Logical_Operator_out404_out1;

  Logical_Operator_out1428_out1 <= in806 XOR in808;

  Logical_Operator_out1429_out1 <= Logical_Operator_out405_out1 XOR Logical_Operator_out406_out1;

  Logical_Operator_out1430_out1 <= in810 XOR in812;

  Logical_Operator_out1431_out1 <= Logical_Operator_out407_out1 XOR Logical_Operator_out408_out1;

  Logical_Operator_out1432_out1 <= in814 XOR in816;

  Logical_Operator_out1433_out1 <= Logical_Operator_out409_out1 XOR Logical_Operator_out410_out1;

  Logical_Operator_out1434_out1 <= in818 XOR in820;

  Logical_Operator_out1435_out1 <= Logical_Operator_out411_out1 XOR Logical_Operator_out412_out1;

  Logical_Operator_out1436_out1 <= in822 XOR in824;

  Logical_Operator_out1437_out1 <= Logical_Operator_out413_out1 XOR Logical_Operator_out414_out1;

  Logical_Operator_out1438_out1 <= in826 XOR in828;

  Logical_Operator_out1439_out1 <= Logical_Operator_out415_out1 XOR Logical_Operator_out416_out1;

  Logical_Operator_out1440_out1 <= in830 XOR in832;

  Logical_Operator_out1441_out1 <= Logical_Operator_out417_out1 XOR Logical_Operator_out418_out1;

  Logical_Operator_out1442_out1 <= in834 XOR in836;

  Logical_Operator_out1443_out1 <= Logical_Operator_out419_out1 XOR Logical_Operator_out420_out1;

  Logical_Operator_out1444_out1 <= in838 XOR in840;

  Logical_Operator_out1445_out1 <= Logical_Operator_out421_out1 XOR Logical_Operator_out422_out1;

  Logical_Operator_out1446_out1 <= in842 XOR in844;

  Logical_Operator_out1447_out1 <= Logical_Operator_out423_out1 XOR Logical_Operator_out424_out1;

  Logical_Operator_out1448_out1 <= in846 XOR in848;

  Logical_Operator_out1449_out1 <= Logical_Operator_out425_out1 XOR Logical_Operator_out426_out1;

  Logical_Operator_out1450_out1 <= in850 XOR in852;

  Logical_Operator_out1451_out1 <= Logical_Operator_out427_out1 XOR Logical_Operator_out428_out1;

  Logical_Operator_out1452_out1 <= in854 XOR in856;

  Logical_Operator_out1453_out1 <= Logical_Operator_out429_out1 XOR Logical_Operator_out430_out1;

  Logical_Operator_out1454_out1 <= in858 XOR in860;

  Logical_Operator_out1455_out1 <= Logical_Operator_out431_out1 XOR Logical_Operator_out432_out1;

  Logical_Operator_out1456_out1 <= in862 XOR in864;

  Logical_Operator_out1457_out1 <= Logical_Operator_out433_out1 XOR Logical_Operator_out434_out1;

  Logical_Operator_out1458_out1 <= in866 XOR in868;

  Logical_Operator_out1459_out1 <= Logical_Operator_out435_out1 XOR Logical_Operator_out436_out1;

  Logical_Operator_out1460_out1 <= in870 XOR in872;

  Logical_Operator_out1461_out1 <= Logical_Operator_out437_out1 XOR Logical_Operator_out438_out1;

  Logical_Operator_out1462_out1 <= in874 XOR in876;

  Logical_Operator_out1463_out1 <= Logical_Operator_out439_out1 XOR Logical_Operator_out440_out1;

  Logical_Operator_out1464_out1 <= in878 XOR in880;

  Logical_Operator_out1465_out1 <= Logical_Operator_out441_out1 XOR Logical_Operator_out442_out1;

  Logical_Operator_out1466_out1 <= in882 XOR in884;

  Logical_Operator_out1467_out1 <= Logical_Operator_out443_out1 XOR Logical_Operator_out444_out1;

  Logical_Operator_out1468_out1 <= in886 XOR in888;

  Logical_Operator_out1469_out1 <= Logical_Operator_out445_out1 XOR Logical_Operator_out446_out1;

  Logical_Operator_out1470_out1 <= in890 XOR in892;

  Logical_Operator_out1471_out1 <= Logical_Operator_out447_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out1472_out1 <= in894 XOR in896;

  Logical_Operator_out1473_out1 <= Logical_Operator_out449_out1 XOR Logical_Operator_out450_out1;

  Logical_Operator_out1474_out1 <= in898 XOR in900;

  Logical_Operator_out1475_out1 <= Logical_Operator_out451_out1 XOR Logical_Operator_out452_out1;

  Logical_Operator_out1476_out1 <= in902 XOR in904;

  Logical_Operator_out1477_out1 <= Logical_Operator_out453_out1 XOR Logical_Operator_out454_out1;

  Logical_Operator_out1478_out1 <= in906 XOR in908;

  Logical_Operator_out1479_out1 <= Logical_Operator_out455_out1 XOR Logical_Operator_out456_out1;

  Logical_Operator_out1480_out1 <= in910 XOR in912;

  Logical_Operator_out1481_out1 <= Logical_Operator_out457_out1 XOR Logical_Operator_out458_out1;

  Logical_Operator_out1482_out1 <= in914 XOR in916;

  Logical_Operator_out1483_out1 <= Logical_Operator_out459_out1 XOR Logical_Operator_out460_out1;

  Logical_Operator_out1484_out1 <= in918 XOR in920;

  Logical_Operator_out1485_out1 <= Logical_Operator_out461_out1 XOR Logical_Operator_out462_out1;

  Logical_Operator_out1486_out1 <= in922 XOR in924;

  Logical_Operator_out1487_out1 <= Logical_Operator_out463_out1 XOR Logical_Operator_out464_out1;

  Logical_Operator_out1488_out1 <= in926 XOR in928;

  Logical_Operator_out1489_out1 <= Logical_Operator_out465_out1 XOR Logical_Operator_out466_out1;

  Logical_Operator_out1490_out1 <= in930 XOR in932;

  Logical_Operator_out1491_out1 <= Logical_Operator_out467_out1 XOR Logical_Operator_out468_out1;

  Logical_Operator_out1492_out1 <= in934 XOR in936;

  Logical_Operator_out1493_out1 <= Logical_Operator_out469_out1 XOR Logical_Operator_out470_out1;

  Logical_Operator_out1494_out1 <= in938 XOR in940;

  Logical_Operator_out1495_out1 <= Logical_Operator_out471_out1 XOR Logical_Operator_out472_out1;

  Logical_Operator_out1496_out1 <= in942 XOR in944;

  Logical_Operator_out1497_out1 <= Logical_Operator_out473_out1 XOR Logical_Operator_out474_out1;

  Logical_Operator_out1498_out1 <= in946 XOR in948;

  Logical_Operator_out1499_out1 <= Logical_Operator_out475_out1 XOR Logical_Operator_out476_out1;

  Logical_Operator_out1500_out1 <= in950 XOR in952;

  Logical_Operator_out1501_out1 <= Logical_Operator_out477_out1 XOR Logical_Operator_out478_out1;

  Logical_Operator_out1502_out1 <= in954 XOR in956;

  Logical_Operator_out1503_out1 <= Logical_Operator_out479_out1 XOR Logical_Operator_out480_out1;

  Logical_Operator_out1504_out1 <= in958 XOR in960;

  Logical_Operator_out1505_out1 <= Logical_Operator_out481_out1 XOR Logical_Operator_out482_out1;

  Logical_Operator_out1506_out1 <= in962 XOR in964;

  Logical_Operator_out1507_out1 <= Logical_Operator_out483_out1 XOR Logical_Operator_out484_out1;

  Logical_Operator_out1508_out1 <= in966 XOR in968;

  Logical_Operator_out1509_out1 <= Logical_Operator_out485_out1 XOR Logical_Operator_out486_out1;

  Logical_Operator_out1510_out1 <= in970 XOR in972;

  Logical_Operator_out1511_out1 <= Logical_Operator_out487_out1 XOR Logical_Operator_out488_out1;

  Logical_Operator_out1512_out1 <= in974 XOR in976;

  Logical_Operator_out1513_out1 <= Logical_Operator_out489_out1 XOR Logical_Operator_out490_out1;

  Logical_Operator_out1514_out1 <= in978 XOR in980;

  Logical_Operator_out1515_out1 <= Logical_Operator_out491_out1 XOR Logical_Operator_out492_out1;

  Logical_Operator_out1516_out1 <= in982 XOR in984;

  Logical_Operator_out1517_out1 <= Logical_Operator_out493_out1 XOR Logical_Operator_out494_out1;

  Logical_Operator_out1518_out1 <= in986 XOR in988;

  Logical_Operator_out1519_out1 <= Logical_Operator_out495_out1 XOR Logical_Operator_out496_out1;

  Logical_Operator_out1520_out1 <= in990 XOR in992;

  Logical_Operator_out1521_out1 <= Logical_Operator_out497_out1 XOR Logical_Operator_out498_out1;

  Logical_Operator_out1522_out1 <= in994 XOR in996;

  Logical_Operator_out1523_out1 <= Logical_Operator_out499_out1 XOR Logical_Operator_out500_out1;

  Logical_Operator_out1524_out1 <= in998 XOR in1000;

  Logical_Operator_out1525_out1 <= Logical_Operator_out501_out1 XOR Logical_Operator_out502_out1;

  Logical_Operator_out1526_out1 <= in1002 XOR in1004;

  Logical_Operator_out1527_out1 <= Logical_Operator_out503_out1 XOR Logical_Operator_out504_out1;

  Logical_Operator_out1528_out1 <= in1006 XOR in1008;

  Logical_Operator_out1529_out1 <= Logical_Operator_out505_out1 XOR Logical_Operator_out506_out1;

  Logical_Operator_out1530_out1 <= in1010 XOR in1012;

  Logical_Operator_out1531_out1 <= Logical_Operator_out507_out1 XOR Logical_Operator_out508_out1;

  Logical_Operator_out1532_out1 <= in1014 XOR in1016;

  Logical_Operator_out1533_out1 <= Logical_Operator_out509_out1 XOR Logical_Operator_out510_out1;

  Logical_Operator_out1534_out1 <= in1018 XOR in1020;

  Logical_Operator_out1535_out1 <= Logical_Operator_out511_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out1536_out1 <= in1022 XOR in1024;

  Logical_Operator_out1537_out1 <= Logical_Operator_out513_out1 XOR Logical_Operator_out514_out1;

  Logical_Operator_out1538_out1 <= in1026 XOR in1028;

  Logical_Operator_out1539_out1 <= Logical_Operator_out515_out1 XOR Logical_Operator_out516_out1;

  Logical_Operator_out1540_out1 <= in1030 XOR in1032;

  Logical_Operator_out1541_out1 <= Logical_Operator_out517_out1 XOR Logical_Operator_out518_out1;

  Logical_Operator_out1542_out1 <= in1034 XOR in1036;

  Logical_Operator_out1543_out1 <= Logical_Operator_out519_out1 XOR Logical_Operator_out520_out1;

  Logical_Operator_out1544_out1 <= in1038 XOR in1040;

  Logical_Operator_out1545_out1 <= Logical_Operator_out521_out1 XOR Logical_Operator_out522_out1;

  Logical_Operator_out1546_out1 <= in1042 XOR in1044;

  Logical_Operator_out1547_out1 <= Logical_Operator_out523_out1 XOR Logical_Operator_out524_out1;

  Logical_Operator_out1548_out1 <= in1046 XOR in1048;

  Logical_Operator_out1549_out1 <= Logical_Operator_out525_out1 XOR Logical_Operator_out526_out1;

  Logical_Operator_out1550_out1 <= in1050 XOR in1052;

  Logical_Operator_out1551_out1 <= Logical_Operator_out527_out1 XOR Logical_Operator_out528_out1;

  Logical_Operator_out1552_out1 <= in1054 XOR in1056;

  Logical_Operator_out1553_out1 <= Logical_Operator_out529_out1 XOR Logical_Operator_out530_out1;

  Logical_Operator_out1554_out1 <= in1058 XOR in1060;

  Logical_Operator_out1555_out1 <= Logical_Operator_out531_out1 XOR Logical_Operator_out532_out1;

  Logical_Operator_out1556_out1 <= in1062 XOR in1064;

  Logical_Operator_out1557_out1 <= Logical_Operator_out533_out1 XOR Logical_Operator_out534_out1;

  Logical_Operator_out1558_out1 <= in1066 XOR in1068;

  Logical_Operator_out1559_out1 <= Logical_Operator_out535_out1 XOR Logical_Operator_out536_out1;

  Logical_Operator_out1560_out1 <= in1070 XOR in1072;

  Logical_Operator_out1561_out1 <= Logical_Operator_out537_out1 XOR Logical_Operator_out538_out1;

  Logical_Operator_out1562_out1 <= in1074 XOR in1076;

  Logical_Operator_out1563_out1 <= Logical_Operator_out539_out1 XOR Logical_Operator_out540_out1;

  Logical_Operator_out1564_out1 <= in1078 XOR in1080;

  Logical_Operator_out1565_out1 <= Logical_Operator_out541_out1 XOR Logical_Operator_out542_out1;

  Logical_Operator_out1566_out1 <= in1082 XOR in1084;

  Logical_Operator_out1567_out1 <= Logical_Operator_out543_out1 XOR Logical_Operator_out544_out1;

  Logical_Operator_out1568_out1 <= in1086 XOR in1088;

  Logical_Operator_out1569_out1 <= Logical_Operator_out545_out1 XOR Logical_Operator_out546_out1;

  Logical_Operator_out1570_out1 <= in1090 XOR in1092;

  Logical_Operator_out1571_out1 <= Logical_Operator_out547_out1 XOR Logical_Operator_out548_out1;

  Logical_Operator_out1572_out1 <= in1094 XOR in1096;

  Logical_Operator_out1573_out1 <= Logical_Operator_out549_out1 XOR Logical_Operator_out550_out1;

  Logical_Operator_out1574_out1 <= in1098 XOR in1100;

  Logical_Operator_out1575_out1 <= Logical_Operator_out551_out1 XOR Logical_Operator_out552_out1;

  Logical_Operator_out1576_out1 <= in1102 XOR in1104;

  Logical_Operator_out1577_out1 <= Logical_Operator_out553_out1 XOR Logical_Operator_out554_out1;

  Logical_Operator_out1578_out1 <= in1106 XOR in1108;

  Logical_Operator_out1579_out1 <= Logical_Operator_out555_out1 XOR Logical_Operator_out556_out1;

  Logical_Operator_out1580_out1 <= in1110 XOR in1112;

  Logical_Operator_out1581_out1 <= Logical_Operator_out557_out1 XOR Logical_Operator_out558_out1;

  Logical_Operator_out1582_out1 <= in1114 XOR in1116;

  Logical_Operator_out1583_out1 <= Logical_Operator_out559_out1 XOR Logical_Operator_out560_out1;

  Logical_Operator_out1584_out1 <= in1118 XOR in1120;

  Logical_Operator_out1585_out1 <= Logical_Operator_out561_out1 XOR Logical_Operator_out562_out1;

  Logical_Operator_out1586_out1 <= in1122 XOR in1124;

  Logical_Operator_out1587_out1 <= Logical_Operator_out563_out1 XOR Logical_Operator_out564_out1;

  Logical_Operator_out1588_out1 <= in1126 XOR in1128;

  Logical_Operator_out1589_out1 <= Logical_Operator_out565_out1 XOR Logical_Operator_out566_out1;

  Logical_Operator_out1590_out1 <= in1130 XOR in1132;

  Logical_Operator_out1591_out1 <= Logical_Operator_out567_out1 XOR Logical_Operator_out568_out1;

  Logical_Operator_out1592_out1 <= in1134 XOR in1136;

  Logical_Operator_out1593_out1 <= Logical_Operator_out569_out1 XOR Logical_Operator_out570_out1;

  Logical_Operator_out1594_out1 <= in1138 XOR in1140;

  Logical_Operator_out1595_out1 <= Logical_Operator_out571_out1 XOR Logical_Operator_out572_out1;

  Logical_Operator_out1596_out1 <= in1142 XOR in1144;

  Logical_Operator_out1597_out1 <= Logical_Operator_out573_out1 XOR Logical_Operator_out574_out1;

  Logical_Operator_out1598_out1 <= in1146 XOR in1148;

  Logical_Operator_out1599_out1 <= Logical_Operator_out575_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out1600_out1 <= in1150 XOR in1152;

  Logical_Operator_out1601_out1 <= Logical_Operator_out577_out1 XOR Logical_Operator_out578_out1;

  Logical_Operator_out1602_out1 <= in1154 XOR in1156;

  Logical_Operator_out1603_out1 <= Logical_Operator_out579_out1 XOR Logical_Operator_out580_out1;

  Logical_Operator_out1604_out1 <= in1158 XOR in1160;

  Logical_Operator_out1605_out1 <= Logical_Operator_out581_out1 XOR Logical_Operator_out582_out1;

  Logical_Operator_out1606_out1 <= in1162 XOR in1164;

  Logical_Operator_out1607_out1 <= Logical_Operator_out583_out1 XOR Logical_Operator_out584_out1;

  Logical_Operator_out1608_out1 <= in1166 XOR in1168;

  Logical_Operator_out1609_out1 <= Logical_Operator_out585_out1 XOR Logical_Operator_out586_out1;

  Logical_Operator_out1610_out1 <= in1170 XOR in1172;

  Logical_Operator_out1611_out1 <= Logical_Operator_out587_out1 XOR Logical_Operator_out588_out1;

  Logical_Operator_out1612_out1 <= in1174 XOR in1176;

  Logical_Operator_out1613_out1 <= Logical_Operator_out589_out1 XOR Logical_Operator_out590_out1;

  Logical_Operator_out1614_out1 <= in1178 XOR in1180;

  Logical_Operator_out1615_out1 <= Logical_Operator_out591_out1 XOR Logical_Operator_out592_out1;

  Logical_Operator_out1616_out1 <= in1182 XOR in1184;

  Logical_Operator_out1617_out1 <= Logical_Operator_out593_out1 XOR Logical_Operator_out594_out1;

  Logical_Operator_out1618_out1 <= in1186 XOR in1188;

  Logical_Operator_out1619_out1 <= Logical_Operator_out595_out1 XOR Logical_Operator_out596_out1;

  Logical_Operator_out1620_out1 <= in1190 XOR in1192;

  Logical_Operator_out1621_out1 <= Logical_Operator_out597_out1 XOR Logical_Operator_out598_out1;

  Logical_Operator_out1622_out1 <= in1194 XOR in1196;

  Logical_Operator_out1623_out1 <= Logical_Operator_out599_out1 XOR Logical_Operator_out600_out1;

  Logical_Operator_out1624_out1 <= in1198 XOR in1200;

  Logical_Operator_out1625_out1 <= Logical_Operator_out601_out1 XOR Logical_Operator_out602_out1;

  Logical_Operator_out1626_out1 <= in1202 XOR in1204;

  Logical_Operator_out1627_out1 <= Logical_Operator_out603_out1 XOR Logical_Operator_out604_out1;

  Logical_Operator_out1628_out1 <= in1206 XOR in1208;

  Logical_Operator_out1629_out1 <= Logical_Operator_out605_out1 XOR Logical_Operator_out606_out1;

  Logical_Operator_out1630_out1 <= in1210 XOR in1212;

  Logical_Operator_out1631_out1 <= Logical_Operator_out607_out1 XOR Logical_Operator_out608_out1;

  Logical_Operator_out1632_out1 <= in1214 XOR in1216;

  Logical_Operator_out1633_out1 <= Logical_Operator_out609_out1 XOR Logical_Operator_out610_out1;

  Logical_Operator_out1634_out1 <= in1218 XOR in1220;

  Logical_Operator_out1635_out1 <= Logical_Operator_out611_out1 XOR Logical_Operator_out612_out1;

  Logical_Operator_out1636_out1 <= in1222 XOR in1224;

  Logical_Operator_out1637_out1 <= Logical_Operator_out613_out1 XOR Logical_Operator_out614_out1;

  Logical_Operator_out1638_out1 <= in1226 XOR in1228;

  Logical_Operator_out1639_out1 <= Logical_Operator_out615_out1 XOR Logical_Operator_out616_out1;

  Logical_Operator_out1640_out1 <= in1230 XOR in1232;

  Logical_Operator_out1641_out1 <= Logical_Operator_out617_out1 XOR Logical_Operator_out618_out1;

  Logical_Operator_out1642_out1 <= in1234 XOR in1236;

  Logical_Operator_out1643_out1 <= Logical_Operator_out619_out1 XOR Logical_Operator_out620_out1;

  Logical_Operator_out1644_out1 <= in1238 XOR in1240;

  Logical_Operator_out1645_out1 <= Logical_Operator_out621_out1 XOR Logical_Operator_out622_out1;

  Logical_Operator_out1646_out1 <= in1242 XOR in1244;

  Logical_Operator_out1647_out1 <= Logical_Operator_out623_out1 XOR Logical_Operator_out624_out1;

  Logical_Operator_out1648_out1 <= in1246 XOR in1248;

  Logical_Operator_out1649_out1 <= Logical_Operator_out625_out1 XOR Logical_Operator_out626_out1;

  Logical_Operator_out1650_out1 <= in1250 XOR in1252;

  Logical_Operator_out1651_out1 <= Logical_Operator_out627_out1 XOR Logical_Operator_out628_out1;

  Logical_Operator_out1652_out1 <= in1254 XOR in1256;

  Logical_Operator_out1653_out1 <= Logical_Operator_out629_out1 XOR Logical_Operator_out630_out1;

  Logical_Operator_out1654_out1 <= in1258 XOR in1260;

  Logical_Operator_out1655_out1 <= Logical_Operator_out631_out1 XOR Logical_Operator_out632_out1;

  Logical_Operator_out1656_out1 <= in1262 XOR in1264;

  Logical_Operator_out1657_out1 <= Logical_Operator_out633_out1 XOR Logical_Operator_out634_out1;

  Logical_Operator_out1658_out1 <= in1266 XOR in1268;

  Logical_Operator_out1659_out1 <= Logical_Operator_out635_out1 XOR Logical_Operator_out636_out1;

  Logical_Operator_out1660_out1 <= in1270 XOR in1272;

  Logical_Operator_out1661_out1 <= Logical_Operator_out637_out1 XOR Logical_Operator_out638_out1;

  Logical_Operator_out1662_out1 <= in1274 XOR in1276;

  Logical_Operator_out1663_out1 <= Logical_Operator_out639_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out1664_out1 <= in1278 XOR in1280;

  Logical_Operator_out1665_out1 <= Logical_Operator_out641_out1 XOR Logical_Operator_out642_out1;

  Logical_Operator_out1666_out1 <= in1282 XOR in1284;

  Logical_Operator_out1667_out1 <= Logical_Operator_out643_out1 XOR Logical_Operator_out644_out1;

  Logical_Operator_out1668_out1 <= in1286 XOR in1288;

  Logical_Operator_out1669_out1 <= Logical_Operator_out645_out1 XOR Logical_Operator_out646_out1;

  Logical_Operator_out1670_out1 <= in1290 XOR in1292;

  Logical_Operator_out1671_out1 <= Logical_Operator_out647_out1 XOR Logical_Operator_out648_out1;

  Logical_Operator_out1672_out1 <= in1294 XOR in1296;

  Logical_Operator_out1673_out1 <= Logical_Operator_out649_out1 XOR Logical_Operator_out650_out1;

  Logical_Operator_out1674_out1 <= in1298 XOR in1300;

  Logical_Operator_out1675_out1 <= Logical_Operator_out651_out1 XOR Logical_Operator_out652_out1;

  Logical_Operator_out1676_out1 <= in1302 XOR in1304;

  Logical_Operator_out1677_out1 <= Logical_Operator_out653_out1 XOR Logical_Operator_out654_out1;

  Logical_Operator_out1678_out1 <= in1306 XOR in1308;

  Logical_Operator_out1679_out1 <= Logical_Operator_out655_out1 XOR Logical_Operator_out656_out1;

  Logical_Operator_out1680_out1 <= in1310 XOR in1312;

  Logical_Operator_out1681_out1 <= Logical_Operator_out657_out1 XOR Logical_Operator_out658_out1;

  Logical_Operator_out1682_out1 <= in1314 XOR in1316;

  Logical_Operator_out1683_out1 <= Logical_Operator_out659_out1 XOR Logical_Operator_out660_out1;

  Logical_Operator_out1684_out1 <= in1318 XOR in1320;

  Logical_Operator_out1685_out1 <= Logical_Operator_out661_out1 XOR Logical_Operator_out662_out1;

  Logical_Operator_out1686_out1 <= in1322 XOR in1324;

  Logical_Operator_out1687_out1 <= Logical_Operator_out663_out1 XOR Logical_Operator_out664_out1;

  Logical_Operator_out1688_out1 <= in1326 XOR in1328;

  Logical_Operator_out1689_out1 <= Logical_Operator_out665_out1 XOR Logical_Operator_out666_out1;

  Logical_Operator_out1690_out1 <= in1330 XOR in1332;

  Logical_Operator_out1691_out1 <= Logical_Operator_out667_out1 XOR Logical_Operator_out668_out1;

  Logical_Operator_out1692_out1 <= in1334 XOR in1336;

  Logical_Operator_out1693_out1 <= Logical_Operator_out669_out1 XOR Logical_Operator_out670_out1;

  Logical_Operator_out1694_out1 <= in1338 XOR in1340;

  Logical_Operator_out1695_out1 <= Logical_Operator_out671_out1 XOR Logical_Operator_out672_out1;

  Logical_Operator_out1696_out1 <= in1342 XOR in1344;

  Logical_Operator_out1697_out1 <= Logical_Operator_out673_out1 XOR Logical_Operator_out674_out1;

  Logical_Operator_out1698_out1 <= in1346 XOR in1348;

  Logical_Operator_out1699_out1 <= Logical_Operator_out675_out1 XOR Logical_Operator_out676_out1;

  Logical_Operator_out1700_out1 <= in1350 XOR in1352;

  Logical_Operator_out1701_out1 <= Logical_Operator_out677_out1 XOR Logical_Operator_out678_out1;

  Logical_Operator_out1702_out1 <= in1354 XOR in1356;

  Logical_Operator_out1703_out1 <= Logical_Operator_out679_out1 XOR Logical_Operator_out680_out1;

  Logical_Operator_out1704_out1 <= in1358 XOR in1360;

  Logical_Operator_out1705_out1 <= Logical_Operator_out681_out1 XOR Logical_Operator_out682_out1;

  Logical_Operator_out1706_out1 <= in1362 XOR in1364;

  Logical_Operator_out1707_out1 <= Logical_Operator_out683_out1 XOR Logical_Operator_out684_out1;

  Logical_Operator_out1708_out1 <= in1366 XOR in1368;

  Logical_Operator_out1709_out1 <= Logical_Operator_out685_out1 XOR Logical_Operator_out686_out1;

  Logical_Operator_out1710_out1 <= in1370 XOR in1372;

  Logical_Operator_out1711_out1 <= Logical_Operator_out687_out1 XOR Logical_Operator_out688_out1;

  Logical_Operator_out1712_out1 <= in1374 XOR in1376;

  Logical_Operator_out1713_out1 <= Logical_Operator_out689_out1 XOR Logical_Operator_out690_out1;

  Logical_Operator_out1714_out1 <= in1378 XOR in1380;

  Logical_Operator_out1715_out1 <= Logical_Operator_out691_out1 XOR Logical_Operator_out692_out1;

  Logical_Operator_out1716_out1 <= in1382 XOR in1384;

  Logical_Operator_out1717_out1 <= Logical_Operator_out693_out1 XOR Logical_Operator_out694_out1;

  Logical_Operator_out1718_out1 <= in1386 XOR in1388;

  Logical_Operator_out1719_out1 <= Logical_Operator_out695_out1 XOR Logical_Operator_out696_out1;

  Logical_Operator_out1720_out1 <= in1390 XOR in1392;

  Logical_Operator_out1721_out1 <= Logical_Operator_out697_out1 XOR Logical_Operator_out698_out1;

  Logical_Operator_out1722_out1 <= in1394 XOR in1396;

  Logical_Operator_out1723_out1 <= Logical_Operator_out699_out1 XOR Logical_Operator_out700_out1;

  Logical_Operator_out1724_out1 <= in1398 XOR in1400;

  Logical_Operator_out1725_out1 <= Logical_Operator_out701_out1 XOR Logical_Operator_out702_out1;

  Logical_Operator_out1726_out1 <= in1402 XOR in1404;

  Logical_Operator_out1727_out1 <= Logical_Operator_out703_out1 XOR Logical_Operator_out704_out1;

  Logical_Operator_out1728_out1 <= in1406 XOR in1408;

  Logical_Operator_out1729_out1 <= Logical_Operator_out705_out1 XOR Logical_Operator_out706_out1;

  Logical_Operator_out1730_out1 <= in1410 XOR in1412;

  Logical_Operator_out1731_out1 <= Logical_Operator_out707_out1 XOR Logical_Operator_out708_out1;

  Logical_Operator_out1732_out1 <= in1414 XOR in1416;

  Logical_Operator_out1733_out1 <= Logical_Operator_out709_out1 XOR Logical_Operator_out710_out1;

  Logical_Operator_out1734_out1 <= in1418 XOR in1420;

  Logical_Operator_out1735_out1 <= Logical_Operator_out711_out1 XOR Logical_Operator_out712_out1;

  Logical_Operator_out1736_out1 <= in1422 XOR in1424;

  Logical_Operator_out1737_out1 <= Logical_Operator_out713_out1 XOR Logical_Operator_out714_out1;

  Logical_Operator_out1738_out1 <= in1426 XOR in1428;

  Logical_Operator_out1739_out1 <= Logical_Operator_out715_out1 XOR Logical_Operator_out716_out1;

  Logical_Operator_out1740_out1 <= in1430 XOR in1432;

  Logical_Operator_out1741_out1 <= Logical_Operator_out717_out1 XOR Logical_Operator_out718_out1;

  Logical_Operator_out1742_out1 <= in1434 XOR in1436;

  Logical_Operator_out1743_out1 <= Logical_Operator_out719_out1 XOR Logical_Operator_out720_out1;

  Logical_Operator_out1744_out1 <= in1438 XOR in1440;

  Logical_Operator_out1745_out1 <= Logical_Operator_out721_out1 XOR Logical_Operator_out722_out1;

  Logical_Operator_out1746_out1 <= in1442 XOR in1444;

  Logical_Operator_out1747_out1 <= Logical_Operator_out723_out1 XOR Logical_Operator_out724_out1;

  Logical_Operator_out1748_out1 <= in1446 XOR in1448;

  Logical_Operator_out1749_out1 <= Logical_Operator_out725_out1 XOR Logical_Operator_out726_out1;

  Logical_Operator_out1750_out1 <= in1450 XOR in1452;

  Logical_Operator_out1751_out1 <= Logical_Operator_out727_out1 XOR Logical_Operator_out728_out1;

  Logical_Operator_out1752_out1 <= in1454 XOR in1456;

  Logical_Operator_out1753_out1 <= Logical_Operator_out729_out1 XOR Logical_Operator_out730_out1;

  Logical_Operator_out1754_out1 <= in1458 XOR in1460;

  Logical_Operator_out1755_out1 <= Logical_Operator_out731_out1 XOR Logical_Operator_out732_out1;

  Logical_Operator_out1756_out1 <= in1462 XOR in1464;

  Logical_Operator_out1757_out1 <= Logical_Operator_out733_out1 XOR Logical_Operator_out734_out1;

  Logical_Operator_out1758_out1 <= in1466 XOR in1468;

  Logical_Operator_out1759_out1 <= Logical_Operator_out735_out1 XOR Logical_Operator_out736_out1;

  Logical_Operator_out1760_out1 <= in1470 XOR in1472;

  Logical_Operator_out1761_out1 <= Logical_Operator_out737_out1 XOR Logical_Operator_out738_out1;

  Logical_Operator_out1762_out1 <= in1474 XOR in1476;

  Logical_Operator_out1763_out1 <= Logical_Operator_out739_out1 XOR Logical_Operator_out740_out1;

  Logical_Operator_out1764_out1 <= in1478 XOR in1480;

  Logical_Operator_out1765_out1 <= Logical_Operator_out741_out1 XOR Logical_Operator_out742_out1;

  Logical_Operator_out1766_out1 <= in1482 XOR in1484;

  Logical_Operator_out1767_out1 <= Logical_Operator_out743_out1 XOR Logical_Operator_out744_out1;

  Logical_Operator_out1768_out1 <= in1486 XOR in1488;

  Logical_Operator_out1769_out1 <= Logical_Operator_out745_out1 XOR Logical_Operator_out746_out1;

  Logical_Operator_out1770_out1 <= in1490 XOR in1492;

  Logical_Operator_out1771_out1 <= Logical_Operator_out747_out1 XOR Logical_Operator_out748_out1;

  Logical_Operator_out1772_out1 <= in1494 XOR in1496;

  Logical_Operator_out1773_out1 <= Logical_Operator_out749_out1 XOR Logical_Operator_out750_out1;

  Logical_Operator_out1774_out1 <= in1498 XOR in1500;

  Logical_Operator_out1775_out1 <= Logical_Operator_out751_out1 XOR Logical_Operator_out752_out1;

  Logical_Operator_out1776_out1 <= in1502 XOR in1504;

  Logical_Operator_out1777_out1 <= Logical_Operator_out753_out1 XOR Logical_Operator_out754_out1;

  Logical_Operator_out1778_out1 <= in1506 XOR in1508;

  Logical_Operator_out1779_out1 <= Logical_Operator_out755_out1 XOR Logical_Operator_out756_out1;

  Logical_Operator_out1780_out1 <= in1510 XOR in1512;

  Logical_Operator_out1781_out1 <= Logical_Operator_out757_out1 XOR Logical_Operator_out758_out1;

  Logical_Operator_out1782_out1 <= in1514 XOR in1516;

  Logical_Operator_out1783_out1 <= Logical_Operator_out759_out1 XOR Logical_Operator_out760_out1;

  Logical_Operator_out1784_out1 <= in1518 XOR in1520;

  Logical_Operator_out1785_out1 <= Logical_Operator_out761_out1 XOR Logical_Operator_out762_out1;

  Logical_Operator_out1786_out1 <= in1522 XOR in1524;

  Logical_Operator_out1787_out1 <= Logical_Operator_out763_out1 XOR Logical_Operator_out764_out1;

  Logical_Operator_out1788_out1 <= in1526 XOR in1528;

  Logical_Operator_out1789_out1 <= Logical_Operator_out765_out1 XOR Logical_Operator_out766_out1;

  Logical_Operator_out1790_out1 <= in1530 XOR in1532;

  Logical_Operator_out1791_out1 <= Logical_Operator_out767_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out1792_out1 <= in1534 XOR in1536;

  Logical_Operator_out1793_out1 <= Logical_Operator_out769_out1 XOR Logical_Operator_out770_out1;

  Logical_Operator_out1794_out1 <= in1538 XOR in1540;

  Logical_Operator_out1795_out1 <= Logical_Operator_out771_out1 XOR Logical_Operator_out772_out1;

  Logical_Operator_out1796_out1 <= in1542 XOR in1544;

  Logical_Operator_out1797_out1 <= Logical_Operator_out773_out1 XOR Logical_Operator_out774_out1;

  Logical_Operator_out1798_out1 <= in1546 XOR in1548;

  Logical_Operator_out1799_out1 <= Logical_Operator_out775_out1 XOR Logical_Operator_out776_out1;

  Logical_Operator_out1800_out1 <= in1550 XOR in1552;

  Logical_Operator_out1801_out1 <= Logical_Operator_out777_out1 XOR Logical_Operator_out778_out1;

  Logical_Operator_out1802_out1 <= in1554 XOR in1556;

  Logical_Operator_out1803_out1 <= Logical_Operator_out779_out1 XOR Logical_Operator_out780_out1;

  Logical_Operator_out1804_out1 <= in1558 XOR in1560;

  Logical_Operator_out1805_out1 <= Logical_Operator_out781_out1 XOR Logical_Operator_out782_out1;

  Logical_Operator_out1806_out1 <= in1562 XOR in1564;

  Logical_Operator_out1807_out1 <= Logical_Operator_out783_out1 XOR Logical_Operator_out784_out1;

  Logical_Operator_out1808_out1 <= in1566 XOR in1568;

  Logical_Operator_out1809_out1 <= Logical_Operator_out785_out1 XOR Logical_Operator_out786_out1;

  Logical_Operator_out1810_out1 <= in1570 XOR in1572;

  Logical_Operator_out1811_out1 <= Logical_Operator_out787_out1 XOR Logical_Operator_out788_out1;

  Logical_Operator_out1812_out1 <= in1574 XOR in1576;

  Logical_Operator_out1813_out1 <= Logical_Operator_out789_out1 XOR Logical_Operator_out790_out1;

  Logical_Operator_out1814_out1 <= in1578 XOR in1580;

  Logical_Operator_out1815_out1 <= Logical_Operator_out791_out1 XOR Logical_Operator_out792_out1;

  Logical_Operator_out1816_out1 <= in1582 XOR in1584;

  Logical_Operator_out1817_out1 <= Logical_Operator_out793_out1 XOR Logical_Operator_out794_out1;

  Logical_Operator_out1818_out1 <= in1586 XOR in1588;

  Logical_Operator_out1819_out1 <= Logical_Operator_out795_out1 XOR Logical_Operator_out796_out1;

  Logical_Operator_out1820_out1 <= in1590 XOR in1592;

  Logical_Operator_out1821_out1 <= Logical_Operator_out797_out1 XOR Logical_Operator_out798_out1;

  Logical_Operator_out1822_out1 <= in1594 XOR in1596;

  Logical_Operator_out1823_out1 <= Logical_Operator_out799_out1 XOR Logical_Operator_out800_out1;

  Logical_Operator_out1824_out1 <= in1598 XOR in1600;

  Logical_Operator_out1825_out1 <= Logical_Operator_out801_out1 XOR Logical_Operator_out802_out1;

  Logical_Operator_out1826_out1 <= in1602 XOR in1604;

  Logical_Operator_out1827_out1 <= Logical_Operator_out803_out1 XOR Logical_Operator_out804_out1;

  Logical_Operator_out1828_out1 <= in1606 XOR in1608;

  Logical_Operator_out1829_out1 <= Logical_Operator_out805_out1 XOR Logical_Operator_out806_out1;

  Logical_Operator_out1830_out1 <= in1610 XOR in1612;

  Logical_Operator_out1831_out1 <= Logical_Operator_out807_out1 XOR Logical_Operator_out808_out1;

  Logical_Operator_out1832_out1 <= in1614 XOR in1616;

  Logical_Operator_out1833_out1 <= Logical_Operator_out809_out1 XOR Logical_Operator_out810_out1;

  Logical_Operator_out1834_out1 <= in1618 XOR in1620;

  Logical_Operator_out1835_out1 <= Logical_Operator_out811_out1 XOR Logical_Operator_out812_out1;

  Logical_Operator_out1836_out1 <= in1622 XOR in1624;

  Logical_Operator_out1837_out1 <= Logical_Operator_out813_out1 XOR Logical_Operator_out814_out1;

  Logical_Operator_out1838_out1 <= in1626 XOR in1628;

  Logical_Operator_out1839_out1 <= Logical_Operator_out815_out1 XOR Logical_Operator_out816_out1;

  Logical_Operator_out1840_out1 <= in1630 XOR in1632;

  Logical_Operator_out1841_out1 <= Logical_Operator_out817_out1 XOR Logical_Operator_out818_out1;

  Logical_Operator_out1842_out1 <= in1634 XOR in1636;

  Logical_Operator_out1843_out1 <= Logical_Operator_out819_out1 XOR Logical_Operator_out820_out1;

  Logical_Operator_out1844_out1 <= in1638 XOR in1640;

  Logical_Operator_out1845_out1 <= Logical_Operator_out821_out1 XOR Logical_Operator_out822_out1;

  Logical_Operator_out1846_out1 <= in1642 XOR in1644;

  Logical_Operator_out1847_out1 <= Logical_Operator_out823_out1 XOR Logical_Operator_out824_out1;

  Logical_Operator_out1848_out1 <= in1646 XOR in1648;

  Logical_Operator_out1849_out1 <= Logical_Operator_out825_out1 XOR Logical_Operator_out826_out1;

  Logical_Operator_out1850_out1 <= in1650 XOR in1652;

  Logical_Operator_out1851_out1 <= Logical_Operator_out827_out1 XOR Logical_Operator_out828_out1;

  Logical_Operator_out1852_out1 <= in1654 XOR in1656;

  Logical_Operator_out1853_out1 <= Logical_Operator_out829_out1 XOR Logical_Operator_out830_out1;

  Logical_Operator_out1854_out1 <= in1658 XOR in1660;

  Logical_Operator_out1855_out1 <= Logical_Operator_out831_out1 XOR Logical_Operator_out832_out1;

  Logical_Operator_out1856_out1 <= in1662 XOR in1664;

  Logical_Operator_out1857_out1 <= Logical_Operator_out833_out1 XOR Logical_Operator_out834_out1;

  Logical_Operator_out1858_out1 <= in1666 XOR in1668;

  Logical_Operator_out1859_out1 <= Logical_Operator_out835_out1 XOR Logical_Operator_out836_out1;

  Logical_Operator_out1860_out1 <= in1670 XOR in1672;

  Logical_Operator_out1861_out1 <= Logical_Operator_out837_out1 XOR Logical_Operator_out838_out1;

  Logical_Operator_out1862_out1 <= in1674 XOR in1676;

  Logical_Operator_out1863_out1 <= Logical_Operator_out839_out1 XOR Logical_Operator_out840_out1;

  Logical_Operator_out1864_out1 <= in1678 XOR in1680;

  Logical_Operator_out1865_out1 <= Logical_Operator_out841_out1 XOR Logical_Operator_out842_out1;

  Logical_Operator_out1866_out1 <= in1682 XOR in1684;

  Logical_Operator_out1867_out1 <= Logical_Operator_out843_out1 XOR Logical_Operator_out844_out1;

  Logical_Operator_out1868_out1 <= in1686 XOR in1688;

  Logical_Operator_out1869_out1 <= Logical_Operator_out845_out1 XOR Logical_Operator_out846_out1;

  Logical_Operator_out1870_out1 <= in1690 XOR in1692;

  Logical_Operator_out1871_out1 <= Logical_Operator_out847_out1 XOR Logical_Operator_out848_out1;

  Logical_Operator_out1872_out1 <= in1694 XOR in1696;

  Logical_Operator_out1873_out1 <= Logical_Operator_out849_out1 XOR Logical_Operator_out850_out1;

  Logical_Operator_out1874_out1 <= in1698 XOR in1700;

  Logical_Operator_out1875_out1 <= Logical_Operator_out851_out1 XOR Logical_Operator_out852_out1;

  Logical_Operator_out1876_out1 <= in1702 XOR in1704;

  Logical_Operator_out1877_out1 <= Logical_Operator_out853_out1 XOR Logical_Operator_out854_out1;

  Logical_Operator_out1878_out1 <= in1706 XOR in1708;

  Logical_Operator_out1879_out1 <= Logical_Operator_out855_out1 XOR Logical_Operator_out856_out1;

  Logical_Operator_out1880_out1 <= in1710 XOR in1712;

  Logical_Operator_out1881_out1 <= Logical_Operator_out857_out1 XOR Logical_Operator_out858_out1;

  Logical_Operator_out1882_out1 <= in1714 XOR in1716;

  Logical_Operator_out1883_out1 <= Logical_Operator_out859_out1 XOR Logical_Operator_out860_out1;

  Logical_Operator_out1884_out1 <= in1718 XOR in1720;

  Logical_Operator_out1885_out1 <= Logical_Operator_out861_out1 XOR Logical_Operator_out862_out1;

  Logical_Operator_out1886_out1 <= in1722 XOR in1724;

  Logical_Operator_out1887_out1 <= Logical_Operator_out863_out1 XOR Logical_Operator_out864_out1;

  Logical_Operator_out1888_out1 <= in1726 XOR in1728;

  Logical_Operator_out1889_out1 <= Logical_Operator_out865_out1 XOR Logical_Operator_out866_out1;

  Logical_Operator_out1890_out1 <= in1730 XOR in1732;

  Logical_Operator_out1891_out1 <= Logical_Operator_out867_out1 XOR Logical_Operator_out868_out1;

  Logical_Operator_out1892_out1 <= in1734 XOR in1736;

  Logical_Operator_out1893_out1 <= Logical_Operator_out869_out1 XOR Logical_Operator_out870_out1;

  Logical_Operator_out1894_out1 <= in1738 XOR in1740;

  Logical_Operator_out1895_out1 <= Logical_Operator_out871_out1 XOR Logical_Operator_out872_out1;

  Logical_Operator_out1896_out1 <= in1742 XOR in1744;

  Logical_Operator_out1897_out1 <= Logical_Operator_out873_out1 XOR Logical_Operator_out874_out1;

  Logical_Operator_out1898_out1 <= in1746 XOR in1748;

  Logical_Operator_out1899_out1 <= Logical_Operator_out875_out1 XOR Logical_Operator_out876_out1;

  Logical_Operator_out1900_out1 <= in1750 XOR in1752;

  Logical_Operator_out1901_out1 <= Logical_Operator_out877_out1 XOR Logical_Operator_out878_out1;

  Logical_Operator_out1902_out1 <= in1754 XOR in1756;

  Logical_Operator_out1903_out1 <= Logical_Operator_out879_out1 XOR Logical_Operator_out880_out1;

  Logical_Operator_out1904_out1 <= in1758 XOR in1760;

  Logical_Operator_out1905_out1 <= Logical_Operator_out881_out1 XOR Logical_Operator_out882_out1;

  Logical_Operator_out1906_out1 <= in1762 XOR in1764;

  Logical_Operator_out1907_out1 <= Logical_Operator_out883_out1 XOR Logical_Operator_out884_out1;

  Logical_Operator_out1908_out1 <= in1766 XOR in1768;

  Logical_Operator_out1909_out1 <= Logical_Operator_out885_out1 XOR Logical_Operator_out886_out1;

  Logical_Operator_out1910_out1 <= in1770 XOR in1772;

  Logical_Operator_out1911_out1 <= Logical_Operator_out887_out1 XOR Logical_Operator_out888_out1;

  Logical_Operator_out1912_out1 <= in1774 XOR in1776;

  Logical_Operator_out1913_out1 <= Logical_Operator_out889_out1 XOR Logical_Operator_out890_out1;

  Logical_Operator_out1914_out1 <= in1778 XOR in1780;

  Logical_Operator_out1915_out1 <= Logical_Operator_out891_out1 XOR Logical_Operator_out892_out1;

  Logical_Operator_out1916_out1 <= in1782 XOR in1784;

  Logical_Operator_out1917_out1 <= Logical_Operator_out893_out1 XOR Logical_Operator_out894_out1;

  Logical_Operator_out1918_out1 <= in1786 XOR in1788;

  Logical_Operator_out1919_out1 <= Logical_Operator_out895_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out1920_out1 <= in1790 XOR in1792;

  Logical_Operator_out1921_out1 <= Logical_Operator_out897_out1 XOR Logical_Operator_out898_out1;

  Logical_Operator_out1922_out1 <= in1794 XOR in1796;

  Logical_Operator_out1923_out1 <= Logical_Operator_out899_out1 XOR Logical_Operator_out900_out1;

  Logical_Operator_out1924_out1 <= in1798 XOR in1800;

  Logical_Operator_out1925_out1 <= Logical_Operator_out901_out1 XOR Logical_Operator_out902_out1;

  Logical_Operator_out1926_out1 <= in1802 XOR in1804;

  Logical_Operator_out1927_out1 <= Logical_Operator_out903_out1 XOR Logical_Operator_out904_out1;

  Logical_Operator_out1928_out1 <= in1806 XOR in1808;

  Logical_Operator_out1929_out1 <= Logical_Operator_out905_out1 XOR Logical_Operator_out906_out1;

  Logical_Operator_out1930_out1 <= in1810 XOR in1812;

  Logical_Operator_out1931_out1 <= Logical_Operator_out907_out1 XOR Logical_Operator_out908_out1;

  Logical_Operator_out1932_out1 <= in1814 XOR in1816;

  Logical_Operator_out1933_out1 <= Logical_Operator_out909_out1 XOR Logical_Operator_out910_out1;

  Logical_Operator_out1934_out1 <= in1818 XOR in1820;

  Logical_Operator_out1935_out1 <= Logical_Operator_out911_out1 XOR Logical_Operator_out912_out1;

  Logical_Operator_out1936_out1 <= in1822 XOR in1824;

  Logical_Operator_out1937_out1 <= Logical_Operator_out913_out1 XOR Logical_Operator_out914_out1;

  Logical_Operator_out1938_out1 <= in1826 XOR in1828;

  Logical_Operator_out1939_out1 <= Logical_Operator_out915_out1 XOR Logical_Operator_out916_out1;

  Logical_Operator_out1940_out1 <= in1830 XOR in1832;

  Logical_Operator_out1941_out1 <= Logical_Operator_out917_out1 XOR Logical_Operator_out918_out1;

  Logical_Operator_out1942_out1 <= in1834 XOR in1836;

  Logical_Operator_out1943_out1 <= Logical_Operator_out919_out1 XOR Logical_Operator_out920_out1;

  Logical_Operator_out1944_out1 <= in1838 XOR in1840;

  Logical_Operator_out1945_out1 <= Logical_Operator_out921_out1 XOR Logical_Operator_out922_out1;

  Logical_Operator_out1946_out1 <= in1842 XOR in1844;

  Logical_Operator_out1947_out1 <= Logical_Operator_out923_out1 XOR Logical_Operator_out924_out1;

  Logical_Operator_out1948_out1 <= in1846 XOR in1848;

  Logical_Operator_out1949_out1 <= Logical_Operator_out925_out1 XOR Logical_Operator_out926_out1;

  Logical_Operator_out1950_out1 <= in1850 XOR in1852;

  Logical_Operator_out1951_out1 <= Logical_Operator_out927_out1 XOR Logical_Operator_out928_out1;

  Logical_Operator_out1952_out1 <= in1854 XOR in1856;

  Logical_Operator_out1953_out1 <= Logical_Operator_out929_out1 XOR Logical_Operator_out930_out1;

  Logical_Operator_out1954_out1 <= in1858 XOR in1860;

  Logical_Operator_out1955_out1 <= Logical_Operator_out931_out1 XOR Logical_Operator_out932_out1;

  Logical_Operator_out1956_out1 <= in1862 XOR in1864;

  Logical_Operator_out1957_out1 <= Logical_Operator_out933_out1 XOR Logical_Operator_out934_out1;

  Logical_Operator_out1958_out1 <= in1866 XOR in1868;

  Logical_Operator_out1959_out1 <= Logical_Operator_out935_out1 XOR Logical_Operator_out936_out1;

  Logical_Operator_out1960_out1 <= in1870 XOR in1872;

  Logical_Operator_out1961_out1 <= Logical_Operator_out937_out1 XOR Logical_Operator_out938_out1;

  Logical_Operator_out1962_out1 <= in1874 XOR in1876;

  Logical_Operator_out1963_out1 <= Logical_Operator_out939_out1 XOR Logical_Operator_out940_out1;

  Logical_Operator_out1964_out1 <= in1878 XOR in1880;

  Logical_Operator_out1965_out1 <= Logical_Operator_out941_out1 XOR Logical_Operator_out942_out1;

  Logical_Operator_out1966_out1 <= in1882 XOR in1884;

  Logical_Operator_out1967_out1 <= Logical_Operator_out943_out1 XOR Logical_Operator_out944_out1;

  Logical_Operator_out1968_out1 <= in1886 XOR in1888;

  Logical_Operator_out1969_out1 <= Logical_Operator_out945_out1 XOR Logical_Operator_out946_out1;

  Logical_Operator_out1970_out1 <= in1890 XOR in1892;

  Logical_Operator_out1971_out1 <= Logical_Operator_out947_out1 XOR Logical_Operator_out948_out1;

  Logical_Operator_out1972_out1 <= in1894 XOR in1896;

  Logical_Operator_out1973_out1 <= Logical_Operator_out949_out1 XOR Logical_Operator_out950_out1;

  Logical_Operator_out1974_out1 <= in1898 XOR in1900;

  Logical_Operator_out1975_out1 <= Logical_Operator_out951_out1 XOR Logical_Operator_out952_out1;

  Logical_Operator_out1976_out1 <= in1902 XOR in1904;

  Logical_Operator_out1977_out1 <= Logical_Operator_out953_out1 XOR Logical_Operator_out954_out1;

  Logical_Operator_out1978_out1 <= in1906 XOR in1908;

  Logical_Operator_out1979_out1 <= Logical_Operator_out955_out1 XOR Logical_Operator_out956_out1;

  Logical_Operator_out1980_out1 <= in1910 XOR in1912;

  Logical_Operator_out1981_out1 <= Logical_Operator_out957_out1 XOR Logical_Operator_out958_out1;

  Logical_Operator_out1982_out1 <= in1914 XOR in1916;

  Logical_Operator_out1983_out1 <= Logical_Operator_out959_out1 XOR Logical_Operator_out960_out1;

  Logical_Operator_out1984_out1 <= in1918 XOR in1920;

  Logical_Operator_out1985_out1 <= Logical_Operator_out961_out1 XOR Logical_Operator_out962_out1;

  Logical_Operator_out1986_out1 <= in1922 XOR in1924;

  Logical_Operator_out1987_out1 <= Logical_Operator_out963_out1 XOR Logical_Operator_out964_out1;

  Logical_Operator_out1988_out1 <= in1926 XOR in1928;

  Logical_Operator_out1989_out1 <= Logical_Operator_out965_out1 XOR Logical_Operator_out966_out1;

  Logical_Operator_out1990_out1 <= in1930 XOR in1932;

  Logical_Operator_out1991_out1 <= Logical_Operator_out967_out1 XOR Logical_Operator_out968_out1;

  Logical_Operator_out1992_out1 <= in1934 XOR in1936;

  Logical_Operator_out1993_out1 <= Logical_Operator_out969_out1 XOR Logical_Operator_out970_out1;

  Logical_Operator_out1994_out1 <= in1938 XOR in1940;

  Logical_Operator_out1995_out1 <= Logical_Operator_out971_out1 XOR Logical_Operator_out972_out1;

  Logical_Operator_out1996_out1 <= in1942 XOR in1944;

  Logical_Operator_out1997_out1 <= Logical_Operator_out973_out1 XOR Logical_Operator_out974_out1;

  Logical_Operator_out1998_out1 <= in1946 XOR in1948;

  Logical_Operator_out1999_out1 <= Logical_Operator_out975_out1 XOR Logical_Operator_out976_out1;

  Logical_Operator_out2000_out1 <= in1950 XOR in1952;

  Logical_Operator_out2001_out1 <= Logical_Operator_out977_out1 XOR Logical_Operator_out978_out1;

  Logical_Operator_out2002_out1 <= in1954 XOR in1956;

  Logical_Operator_out2003_out1 <= Logical_Operator_out979_out1 XOR Logical_Operator_out980_out1;

  Logical_Operator_out2004_out1 <= in1958 XOR in1960;

  Logical_Operator_out2005_out1 <= Logical_Operator_out981_out1 XOR Logical_Operator_out982_out1;

  Logical_Operator_out2006_out1 <= in1962 XOR in1964;

  Logical_Operator_out2007_out1 <= Logical_Operator_out983_out1 XOR Logical_Operator_out984_out1;

  Logical_Operator_out2008_out1 <= in1966 XOR in1968;

  Logical_Operator_out2009_out1 <= Logical_Operator_out985_out1 XOR Logical_Operator_out986_out1;

  Logical_Operator_out2010_out1 <= in1970 XOR in1972;

  Logical_Operator_out2011_out1 <= Logical_Operator_out987_out1 XOR Logical_Operator_out988_out1;

  Logical_Operator_out2012_out1 <= in1974 XOR in1976;

  Logical_Operator_out2013_out1 <= Logical_Operator_out989_out1 XOR Logical_Operator_out990_out1;

  Logical_Operator_out2014_out1 <= in1978 XOR in1980;

  Logical_Operator_out2015_out1 <= Logical_Operator_out991_out1 XOR Logical_Operator_out992_out1;

  Logical_Operator_out2016_out1 <= in1982 XOR in1984;

  Logical_Operator_out2017_out1 <= Logical_Operator_out993_out1 XOR Logical_Operator_out994_out1;

  Logical_Operator_out2018_out1 <= in1986 XOR in1988;

  Logical_Operator_out2019_out1 <= Logical_Operator_out995_out1 XOR Logical_Operator_out996_out1;

  Logical_Operator_out2020_out1 <= in1990 XOR in1992;

  Logical_Operator_out2021_out1 <= Logical_Operator_out997_out1 XOR Logical_Operator_out998_out1;

  Logical_Operator_out2022_out1 <= in1994 XOR in1996;

  Logical_Operator_out2023_out1 <= Logical_Operator_out999_out1 XOR Logical_Operator_out1000_out1;

  Logical_Operator_out2024_out1 <= in1998 XOR in2000;

  Logical_Operator_out2025_out1 <= Logical_Operator_out1001_out1 XOR Logical_Operator_out1002_out1;

  Logical_Operator_out2026_out1 <= in2002 XOR in2004;

  Logical_Operator_out2027_out1 <= Logical_Operator_out1003_out1 XOR Logical_Operator_out1004_out1;

  Logical_Operator_out2028_out1 <= in2006 XOR in2008;

  Logical_Operator_out2029_out1 <= Logical_Operator_out1005_out1 XOR Logical_Operator_out1006_out1;

  Logical_Operator_out2030_out1 <= in2010 XOR in2012;

  Logical_Operator_out2031_out1 <= Logical_Operator_out1007_out1 XOR Logical_Operator_out1008_out1;

  Logical_Operator_out2032_out1 <= in2014 XOR in2016;

  Logical_Operator_out2033_out1 <= Logical_Operator_out1009_out1 XOR Logical_Operator_out1010_out1;

  Logical_Operator_out2034_out1 <= in2018 XOR in2020;

  Logical_Operator_out2035_out1 <= Logical_Operator_out1011_out1 XOR Logical_Operator_out1012_out1;

  Logical_Operator_out2036_out1 <= in2022 XOR in2024;

  Logical_Operator_out2037_out1 <= Logical_Operator_out1013_out1 XOR Logical_Operator_out1014_out1;

  Logical_Operator_out2038_out1 <= in2026 XOR in2028;

  Logical_Operator_out2039_out1 <= Logical_Operator_out1015_out1 XOR Logical_Operator_out1016_out1;

  Logical_Operator_out2040_out1 <= in2030 XOR in2032;

  Logical_Operator_out2041_out1 <= Logical_Operator_out1017_out1 XOR Logical_Operator_out1018_out1;

  Logical_Operator_out2042_out1 <= in2034 XOR in2036;

  Logical_Operator_out2043_out1 <= Logical_Operator_out1019_out1 XOR Logical_Operator_out1020_out1;

  Logical_Operator_out2044_out1 <= in2038 XOR in2040;

  Logical_Operator_out2045_out1 <= Logical_Operator_out1021_out1 XOR Logical_Operator_out1022_out1;

  Logical_Operator_out2046_out1 <= in2042 XOR in2044;

  Logical_Operator_out2047_out1 <= Logical_Operator_out1023_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out2048_out1 <= in2046 XOR in2048;

  Logical_Operator_out2049_out1 <= Logical_Operator_out1025_out1 XOR Logical_Operator_out1027_out1;

  Logical_Operator_out2050_out1 <= Logical_Operator_out1026_out1 XOR Logical_Operator_out1028_out1;

  Logical_Operator_out2051_out1 <= Logical_Operator_out2_out1 XOR Logical_Operator_out4_out1;

  Logical_Operator_out2052_out1 <= in4 XOR in8;

  Logical_Operator_out2053_out1 <= Logical_Operator_out1029_out1 XOR Logical_Operator_out1031_out1;

  Logical_Operator_out2054_out1 <= Logical_Operator_out1030_out1 XOR Logical_Operator_out1032_out1;

  Logical_Operator_out2055_out1 <= Logical_Operator_out6_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out2056_out1 <= in12 XOR in16;

  Logical_Operator_out2057_out1 <= Logical_Operator_out1033_out1 XOR Logical_Operator_out1035_out1;

  Logical_Operator_out2058_out1 <= Logical_Operator_out1034_out1 XOR Logical_Operator_out1036_out1;

  Logical_Operator_out2059_out1 <= Logical_Operator_out10_out1 XOR Logical_Operator_out12_out1;

  Logical_Operator_out2060_out1 <= in20 XOR in24;

  Logical_Operator_out2061_out1 <= Logical_Operator_out1037_out1 XOR Logical_Operator_out1039_out1;

  Logical_Operator_out2062_out1 <= Logical_Operator_out1038_out1 XOR Logical_Operator_out1040_out1;

  Logical_Operator_out2063_out1 <= Logical_Operator_out14_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out2064_out1 <= in28 XOR in32;

  Logical_Operator_out2065_out1 <= Logical_Operator_out1041_out1 XOR Logical_Operator_out1043_out1;

  Logical_Operator_out2066_out1 <= Logical_Operator_out1042_out1 XOR Logical_Operator_out1044_out1;

  Logical_Operator_out2067_out1 <= Logical_Operator_out18_out1 XOR Logical_Operator_out20_out1;

  Logical_Operator_out2068_out1 <= in36 XOR in40;

  Logical_Operator_out2069_out1 <= Logical_Operator_out1045_out1 XOR Logical_Operator_out1047_out1;

  Logical_Operator_out2070_out1 <= Logical_Operator_out1046_out1 XOR Logical_Operator_out1048_out1;

  Logical_Operator_out2071_out1 <= Logical_Operator_out22_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out2072_out1 <= in44 XOR in48;

  Logical_Operator_out2073_out1 <= Logical_Operator_out1049_out1 XOR Logical_Operator_out1051_out1;

  Logical_Operator_out2074_out1 <= Logical_Operator_out1050_out1 XOR Logical_Operator_out1052_out1;

  Logical_Operator_out2075_out1 <= Logical_Operator_out26_out1 XOR Logical_Operator_out28_out1;

  Logical_Operator_out2076_out1 <= in52 XOR in56;

  Logical_Operator_out2077_out1 <= Logical_Operator_out1053_out1 XOR Logical_Operator_out1055_out1;

  Logical_Operator_out2078_out1 <= Logical_Operator_out1054_out1 XOR Logical_Operator_out1056_out1;

  Logical_Operator_out2079_out1 <= Logical_Operator_out30_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out2080_out1 <= in60 XOR in64;

  Logical_Operator_out2081_out1 <= Logical_Operator_out1057_out1 XOR Logical_Operator_out1059_out1;

  Logical_Operator_out2082_out1 <= Logical_Operator_out1058_out1 XOR Logical_Operator_out1060_out1;

  Logical_Operator_out2083_out1 <= Logical_Operator_out34_out1 XOR Logical_Operator_out36_out1;

  Logical_Operator_out2084_out1 <= in68 XOR in72;

  Logical_Operator_out2085_out1 <= Logical_Operator_out1061_out1 XOR Logical_Operator_out1063_out1;

  Logical_Operator_out2086_out1 <= Logical_Operator_out1062_out1 XOR Logical_Operator_out1064_out1;

  Logical_Operator_out2087_out1 <= Logical_Operator_out38_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out2088_out1 <= in76 XOR in80;

  Logical_Operator_out2089_out1 <= Logical_Operator_out1065_out1 XOR Logical_Operator_out1067_out1;

  Logical_Operator_out2090_out1 <= Logical_Operator_out1066_out1 XOR Logical_Operator_out1068_out1;

  Logical_Operator_out2091_out1 <= Logical_Operator_out42_out1 XOR Logical_Operator_out44_out1;

  Logical_Operator_out2092_out1 <= in84 XOR in88;

  Logical_Operator_out2093_out1 <= Logical_Operator_out1069_out1 XOR Logical_Operator_out1071_out1;

  Logical_Operator_out2094_out1 <= Logical_Operator_out1070_out1 XOR Logical_Operator_out1072_out1;

  Logical_Operator_out2095_out1 <= Logical_Operator_out46_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out2096_out1 <= in92 XOR in96;

  Logical_Operator_out2097_out1 <= Logical_Operator_out1073_out1 XOR Logical_Operator_out1075_out1;

  Logical_Operator_out2098_out1 <= Logical_Operator_out1074_out1 XOR Logical_Operator_out1076_out1;

  Logical_Operator_out2099_out1 <= Logical_Operator_out50_out1 XOR Logical_Operator_out52_out1;

  Logical_Operator_out2100_out1 <= in100 XOR in104;

  Logical_Operator_out2101_out1 <= Logical_Operator_out1077_out1 XOR Logical_Operator_out1079_out1;

  Logical_Operator_out2102_out1 <= Logical_Operator_out1078_out1 XOR Logical_Operator_out1080_out1;

  Logical_Operator_out2103_out1 <= Logical_Operator_out54_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out2104_out1 <= in108 XOR in112;

  Logical_Operator_out2105_out1 <= Logical_Operator_out1081_out1 XOR Logical_Operator_out1083_out1;

  Logical_Operator_out2106_out1 <= Logical_Operator_out1082_out1 XOR Logical_Operator_out1084_out1;

  Logical_Operator_out2107_out1 <= Logical_Operator_out58_out1 XOR Logical_Operator_out60_out1;

  Logical_Operator_out2108_out1 <= in116 XOR in120;

  Logical_Operator_out2109_out1 <= Logical_Operator_out1085_out1 XOR Logical_Operator_out1087_out1;

  Logical_Operator_out2110_out1 <= Logical_Operator_out1086_out1 XOR Logical_Operator_out1088_out1;

  Logical_Operator_out2111_out1 <= Logical_Operator_out62_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out2112_out1 <= in124 XOR in128;

  Logical_Operator_out2113_out1 <= Logical_Operator_out1089_out1 XOR Logical_Operator_out1091_out1;

  Logical_Operator_out2114_out1 <= Logical_Operator_out1090_out1 XOR Logical_Operator_out1092_out1;

  Logical_Operator_out2115_out1 <= Logical_Operator_out66_out1 XOR Logical_Operator_out68_out1;

  Logical_Operator_out2116_out1 <= in132 XOR in136;

  Logical_Operator_out2117_out1 <= Logical_Operator_out1093_out1 XOR Logical_Operator_out1095_out1;

  Logical_Operator_out2118_out1 <= Logical_Operator_out1094_out1 XOR Logical_Operator_out1096_out1;

  Logical_Operator_out2119_out1 <= Logical_Operator_out70_out1 XOR Logical_Operator_out72_out1;

  Logical_Operator_out2120_out1 <= in140 XOR in144;

  Logical_Operator_out2121_out1 <= Logical_Operator_out1097_out1 XOR Logical_Operator_out1099_out1;

  Logical_Operator_out2122_out1 <= Logical_Operator_out1098_out1 XOR Logical_Operator_out1100_out1;

  Logical_Operator_out2123_out1 <= Logical_Operator_out74_out1 XOR Logical_Operator_out76_out1;

  Logical_Operator_out2124_out1 <= in148 XOR in152;

  Logical_Operator_out2125_out1 <= Logical_Operator_out1101_out1 XOR Logical_Operator_out1103_out1;

  Logical_Operator_out2126_out1 <= Logical_Operator_out1102_out1 XOR Logical_Operator_out1104_out1;

  Logical_Operator_out2127_out1 <= Logical_Operator_out78_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out2128_out1 <= in156 XOR in160;

  Logical_Operator_out2129_out1 <= Logical_Operator_out1105_out1 XOR Logical_Operator_out1107_out1;

  Logical_Operator_out2130_out1 <= Logical_Operator_out1106_out1 XOR Logical_Operator_out1108_out1;

  Logical_Operator_out2131_out1 <= Logical_Operator_out82_out1 XOR Logical_Operator_out84_out1;

  Logical_Operator_out2132_out1 <= in164 XOR in168;

  Logical_Operator_out2133_out1 <= Logical_Operator_out1109_out1 XOR Logical_Operator_out1111_out1;

  Logical_Operator_out2134_out1 <= Logical_Operator_out1110_out1 XOR Logical_Operator_out1112_out1;

  Logical_Operator_out2135_out1 <= Logical_Operator_out86_out1 XOR Logical_Operator_out88_out1;

  Logical_Operator_out2136_out1 <= in172 XOR in176;

  Logical_Operator_out2137_out1 <= Logical_Operator_out1113_out1 XOR Logical_Operator_out1115_out1;

  Logical_Operator_out2138_out1 <= Logical_Operator_out1114_out1 XOR Logical_Operator_out1116_out1;

  Logical_Operator_out2139_out1 <= Logical_Operator_out90_out1 XOR Logical_Operator_out92_out1;

  Logical_Operator_out2140_out1 <= in180 XOR in184;

  Logical_Operator_out2141_out1 <= Logical_Operator_out1117_out1 XOR Logical_Operator_out1119_out1;

  Logical_Operator_out2142_out1 <= Logical_Operator_out1118_out1 XOR Logical_Operator_out1120_out1;

  Logical_Operator_out2143_out1 <= Logical_Operator_out94_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out2144_out1 <= in188 XOR in192;

  Logical_Operator_out2145_out1 <= Logical_Operator_out1121_out1 XOR Logical_Operator_out1123_out1;

  Logical_Operator_out2146_out1 <= Logical_Operator_out1122_out1 XOR Logical_Operator_out1124_out1;

  Logical_Operator_out2147_out1 <= Logical_Operator_out98_out1 XOR Logical_Operator_out100_out1;

  Logical_Operator_out2148_out1 <= in196 XOR in200;

  Logical_Operator_out2149_out1 <= Logical_Operator_out1125_out1 XOR Logical_Operator_out1127_out1;

  Logical_Operator_out2150_out1 <= Logical_Operator_out1126_out1 XOR Logical_Operator_out1128_out1;

  Logical_Operator_out2151_out1 <= Logical_Operator_out102_out1 XOR Logical_Operator_out104_out1;

  Logical_Operator_out2152_out1 <= in204 XOR in208;

  Logical_Operator_out2153_out1 <= Logical_Operator_out1129_out1 XOR Logical_Operator_out1131_out1;

  Logical_Operator_out2154_out1 <= Logical_Operator_out1130_out1 XOR Logical_Operator_out1132_out1;

  Logical_Operator_out2155_out1 <= Logical_Operator_out106_out1 XOR Logical_Operator_out108_out1;

  Logical_Operator_out2156_out1 <= in212 XOR in216;

  Logical_Operator_out2157_out1 <= Logical_Operator_out1133_out1 XOR Logical_Operator_out1135_out1;

  Logical_Operator_out2158_out1 <= Logical_Operator_out1134_out1 XOR Logical_Operator_out1136_out1;

  Logical_Operator_out2159_out1 <= Logical_Operator_out110_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out2160_out1 <= in220 XOR in224;

  Logical_Operator_out2161_out1 <= Logical_Operator_out1137_out1 XOR Logical_Operator_out1139_out1;

  Logical_Operator_out2162_out1 <= Logical_Operator_out1138_out1 XOR Logical_Operator_out1140_out1;

  Logical_Operator_out2163_out1 <= Logical_Operator_out114_out1 XOR Logical_Operator_out116_out1;

  Logical_Operator_out2164_out1 <= in228 XOR in232;

  Logical_Operator_out2165_out1 <= Logical_Operator_out1141_out1 XOR Logical_Operator_out1143_out1;

  Logical_Operator_out2166_out1 <= Logical_Operator_out1142_out1 XOR Logical_Operator_out1144_out1;

  Logical_Operator_out2167_out1 <= Logical_Operator_out118_out1 XOR Logical_Operator_out120_out1;

  Logical_Operator_out2168_out1 <= in236 XOR in240;

  Logical_Operator_out2169_out1 <= Logical_Operator_out1145_out1 XOR Logical_Operator_out1147_out1;

  Logical_Operator_out2170_out1 <= Logical_Operator_out1146_out1 XOR Logical_Operator_out1148_out1;

  Logical_Operator_out2171_out1 <= Logical_Operator_out122_out1 XOR Logical_Operator_out124_out1;

  Logical_Operator_out2172_out1 <= in244 XOR in248;

  Logical_Operator_out2173_out1 <= Logical_Operator_out1149_out1 XOR Logical_Operator_out1151_out1;

  Logical_Operator_out2174_out1 <= Logical_Operator_out1150_out1 XOR Logical_Operator_out1152_out1;

  Logical_Operator_out2175_out1 <= Logical_Operator_out126_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out2176_out1 <= in252 XOR in256;

  Logical_Operator_out2177_out1 <= Logical_Operator_out1153_out1 XOR Logical_Operator_out1155_out1;

  Logical_Operator_out2178_out1 <= Logical_Operator_out1154_out1 XOR Logical_Operator_out1156_out1;

  Logical_Operator_out2179_out1 <= Logical_Operator_out130_out1 XOR Logical_Operator_out132_out1;

  Logical_Operator_out2180_out1 <= in260 XOR in264;

  Logical_Operator_out2181_out1 <= Logical_Operator_out1157_out1 XOR Logical_Operator_out1159_out1;

  Logical_Operator_out2182_out1 <= Logical_Operator_out1158_out1 XOR Logical_Operator_out1160_out1;

  Logical_Operator_out2183_out1 <= Logical_Operator_out134_out1 XOR Logical_Operator_out136_out1;

  Logical_Operator_out2184_out1 <= in268 XOR in272;

  Logical_Operator_out2185_out1 <= Logical_Operator_out1161_out1 XOR Logical_Operator_out1163_out1;

  Logical_Operator_out2186_out1 <= Logical_Operator_out1162_out1 XOR Logical_Operator_out1164_out1;

  Logical_Operator_out2187_out1 <= Logical_Operator_out138_out1 XOR Logical_Operator_out140_out1;

  Logical_Operator_out2188_out1 <= in276 XOR in280;

  Logical_Operator_out2189_out1 <= Logical_Operator_out1165_out1 XOR Logical_Operator_out1167_out1;

  Logical_Operator_out2190_out1 <= Logical_Operator_out1166_out1 XOR Logical_Operator_out1168_out1;

  Logical_Operator_out2191_out1 <= Logical_Operator_out142_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out2192_out1 <= in284 XOR in288;

  Logical_Operator_out2193_out1 <= Logical_Operator_out1169_out1 XOR Logical_Operator_out1171_out1;

  Logical_Operator_out2194_out1 <= Logical_Operator_out1170_out1 XOR Logical_Operator_out1172_out1;

  Logical_Operator_out2195_out1 <= Logical_Operator_out146_out1 XOR Logical_Operator_out148_out1;

  Logical_Operator_out2196_out1 <= in292 XOR in296;

  Logical_Operator_out2197_out1 <= Logical_Operator_out1173_out1 XOR Logical_Operator_out1175_out1;

  Logical_Operator_out2198_out1 <= Logical_Operator_out1174_out1 XOR Logical_Operator_out1176_out1;

  Logical_Operator_out2199_out1 <= Logical_Operator_out150_out1 XOR Logical_Operator_out152_out1;

  Logical_Operator_out2200_out1 <= in300 XOR in304;

  Logical_Operator_out2201_out1 <= Logical_Operator_out1177_out1 XOR Logical_Operator_out1179_out1;

  Logical_Operator_out2202_out1 <= Logical_Operator_out1178_out1 XOR Logical_Operator_out1180_out1;

  Logical_Operator_out2203_out1 <= Logical_Operator_out154_out1 XOR Logical_Operator_out156_out1;

  Logical_Operator_out2204_out1 <= in308 XOR in312;

  Logical_Operator_out2205_out1 <= Logical_Operator_out1181_out1 XOR Logical_Operator_out1183_out1;

  Logical_Operator_out2206_out1 <= Logical_Operator_out1182_out1 XOR Logical_Operator_out1184_out1;

  Logical_Operator_out2207_out1 <= Logical_Operator_out158_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out2208_out1 <= in316 XOR in320;

  Logical_Operator_out2209_out1 <= Logical_Operator_out1185_out1 XOR Logical_Operator_out1187_out1;

  Logical_Operator_out2210_out1 <= Logical_Operator_out1186_out1 XOR Logical_Operator_out1188_out1;

  Logical_Operator_out2211_out1 <= Logical_Operator_out162_out1 XOR Logical_Operator_out164_out1;

  Logical_Operator_out2212_out1 <= in324 XOR in328;

  Logical_Operator_out2213_out1 <= Logical_Operator_out1189_out1 XOR Logical_Operator_out1191_out1;

  Logical_Operator_out2214_out1 <= Logical_Operator_out1190_out1 XOR Logical_Operator_out1192_out1;

  Logical_Operator_out2215_out1 <= Logical_Operator_out166_out1 XOR Logical_Operator_out168_out1;

  Logical_Operator_out2216_out1 <= in332 XOR in336;

  Logical_Operator_out2217_out1 <= Logical_Operator_out1193_out1 XOR Logical_Operator_out1195_out1;

  Logical_Operator_out2218_out1 <= Logical_Operator_out1194_out1 XOR Logical_Operator_out1196_out1;

  Logical_Operator_out2219_out1 <= Logical_Operator_out170_out1 XOR Logical_Operator_out172_out1;

  Logical_Operator_out2220_out1 <= in340 XOR in344;

  Logical_Operator_out2221_out1 <= Logical_Operator_out1197_out1 XOR Logical_Operator_out1199_out1;

  Logical_Operator_out2222_out1 <= Logical_Operator_out1198_out1 XOR Logical_Operator_out1200_out1;

  Logical_Operator_out2223_out1 <= Logical_Operator_out174_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out2224_out1 <= in348 XOR in352;

  Logical_Operator_out2225_out1 <= Logical_Operator_out1201_out1 XOR Logical_Operator_out1203_out1;

  Logical_Operator_out2226_out1 <= Logical_Operator_out1202_out1 XOR Logical_Operator_out1204_out1;

  Logical_Operator_out2227_out1 <= Logical_Operator_out178_out1 XOR Logical_Operator_out180_out1;

  Logical_Operator_out2228_out1 <= in356 XOR in360;

  Logical_Operator_out2229_out1 <= Logical_Operator_out1205_out1 XOR Logical_Operator_out1207_out1;

  Logical_Operator_out2230_out1 <= Logical_Operator_out1206_out1 XOR Logical_Operator_out1208_out1;

  Logical_Operator_out2231_out1 <= Logical_Operator_out182_out1 XOR Logical_Operator_out184_out1;

  Logical_Operator_out2232_out1 <= in364 XOR in368;

  Logical_Operator_out2233_out1 <= Logical_Operator_out1209_out1 XOR Logical_Operator_out1211_out1;

  Logical_Operator_out2234_out1 <= Logical_Operator_out1210_out1 XOR Logical_Operator_out1212_out1;

  Logical_Operator_out2235_out1 <= Logical_Operator_out186_out1 XOR Logical_Operator_out188_out1;

  Logical_Operator_out2236_out1 <= in372 XOR in376;

  Logical_Operator_out2237_out1 <= Logical_Operator_out1213_out1 XOR Logical_Operator_out1215_out1;

  Logical_Operator_out2238_out1 <= Logical_Operator_out1214_out1 XOR Logical_Operator_out1216_out1;

  Logical_Operator_out2239_out1 <= Logical_Operator_out190_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out2240_out1 <= in380 XOR in384;

  Logical_Operator_out2241_out1 <= Logical_Operator_out1217_out1 XOR Logical_Operator_out1219_out1;

  Logical_Operator_out2242_out1 <= Logical_Operator_out1218_out1 XOR Logical_Operator_out1220_out1;

  Logical_Operator_out2243_out1 <= Logical_Operator_out194_out1 XOR Logical_Operator_out196_out1;

  Logical_Operator_out2244_out1 <= in388 XOR in392;

  Logical_Operator_out2245_out1 <= Logical_Operator_out1221_out1 XOR Logical_Operator_out1223_out1;

  Logical_Operator_out2246_out1 <= Logical_Operator_out1222_out1 XOR Logical_Operator_out1224_out1;

  Logical_Operator_out2247_out1 <= Logical_Operator_out198_out1 XOR Logical_Operator_out200_out1;

  Logical_Operator_out2248_out1 <= in396 XOR in400;

  Logical_Operator_out2249_out1 <= Logical_Operator_out1225_out1 XOR Logical_Operator_out1227_out1;

  Logical_Operator_out2250_out1 <= Logical_Operator_out1226_out1 XOR Logical_Operator_out1228_out1;

  Logical_Operator_out2251_out1 <= Logical_Operator_out202_out1 XOR Logical_Operator_out204_out1;

  Logical_Operator_out2252_out1 <= in404 XOR in408;

  Logical_Operator_out2253_out1 <= Logical_Operator_out1229_out1 XOR Logical_Operator_out1231_out1;

  Logical_Operator_out2254_out1 <= Logical_Operator_out1230_out1 XOR Logical_Operator_out1232_out1;

  Logical_Operator_out2255_out1 <= Logical_Operator_out206_out1 XOR Logical_Operator_out208_out1;

  Logical_Operator_out2256_out1 <= in412 XOR in416;

  Logical_Operator_out2257_out1 <= Logical_Operator_out1233_out1 XOR Logical_Operator_out1235_out1;

  Logical_Operator_out2258_out1 <= Logical_Operator_out1234_out1 XOR Logical_Operator_out1236_out1;

  Logical_Operator_out2259_out1 <= Logical_Operator_out210_out1 XOR Logical_Operator_out212_out1;

  Logical_Operator_out2260_out1 <= in420 XOR in424;

  Logical_Operator_out2261_out1 <= Logical_Operator_out1237_out1 XOR Logical_Operator_out1239_out1;

  Logical_Operator_out2262_out1 <= Logical_Operator_out1238_out1 XOR Logical_Operator_out1240_out1;

  Logical_Operator_out2263_out1 <= Logical_Operator_out214_out1 XOR Logical_Operator_out216_out1;

  Logical_Operator_out2264_out1 <= in428 XOR in432;

  Logical_Operator_out2265_out1 <= Logical_Operator_out1241_out1 XOR Logical_Operator_out1243_out1;

  Logical_Operator_out2266_out1 <= Logical_Operator_out1242_out1 XOR Logical_Operator_out1244_out1;

  Logical_Operator_out2267_out1 <= Logical_Operator_out218_out1 XOR Logical_Operator_out220_out1;

  Logical_Operator_out2268_out1 <= in436 XOR in440;

  Logical_Operator_out2269_out1 <= Logical_Operator_out1245_out1 XOR Logical_Operator_out1247_out1;

  Logical_Operator_out2270_out1 <= Logical_Operator_out1246_out1 XOR Logical_Operator_out1248_out1;

  Logical_Operator_out2271_out1 <= Logical_Operator_out222_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out2272_out1 <= in444 XOR in448;

  Logical_Operator_out2273_out1 <= Logical_Operator_out1249_out1 XOR Logical_Operator_out1251_out1;

  Logical_Operator_out2274_out1 <= Logical_Operator_out1250_out1 XOR Logical_Operator_out1252_out1;

  Logical_Operator_out2275_out1 <= Logical_Operator_out226_out1 XOR Logical_Operator_out228_out1;

  Logical_Operator_out2276_out1 <= in452 XOR in456;

  Logical_Operator_out2277_out1 <= Logical_Operator_out1253_out1 XOR Logical_Operator_out1255_out1;

  Logical_Operator_out2278_out1 <= Logical_Operator_out1254_out1 XOR Logical_Operator_out1256_out1;

  Logical_Operator_out2279_out1 <= Logical_Operator_out230_out1 XOR Logical_Operator_out232_out1;

  Logical_Operator_out2280_out1 <= in460 XOR in464;

  Logical_Operator_out2281_out1 <= Logical_Operator_out1257_out1 XOR Logical_Operator_out1259_out1;

  Logical_Operator_out2282_out1 <= Logical_Operator_out1258_out1 XOR Logical_Operator_out1260_out1;

  Logical_Operator_out2283_out1 <= Logical_Operator_out234_out1 XOR Logical_Operator_out236_out1;

  Logical_Operator_out2284_out1 <= in468 XOR in472;

  Logical_Operator_out2285_out1 <= Logical_Operator_out1261_out1 XOR Logical_Operator_out1263_out1;

  Logical_Operator_out2286_out1 <= Logical_Operator_out1262_out1 XOR Logical_Operator_out1264_out1;

  Logical_Operator_out2287_out1 <= Logical_Operator_out238_out1 XOR Logical_Operator_out240_out1;

  Logical_Operator_out2288_out1 <= in476 XOR in480;

  Logical_Operator_out2289_out1 <= Logical_Operator_out1265_out1 XOR Logical_Operator_out1267_out1;

  Logical_Operator_out2290_out1 <= Logical_Operator_out1266_out1 XOR Logical_Operator_out1268_out1;

  Logical_Operator_out2291_out1 <= Logical_Operator_out242_out1 XOR Logical_Operator_out244_out1;

  Logical_Operator_out2292_out1 <= in484 XOR in488;

  Logical_Operator_out2293_out1 <= Logical_Operator_out1269_out1 XOR Logical_Operator_out1271_out1;

  Logical_Operator_out2294_out1 <= Logical_Operator_out1270_out1 XOR Logical_Operator_out1272_out1;

  Logical_Operator_out2295_out1 <= Logical_Operator_out246_out1 XOR Logical_Operator_out248_out1;

  Logical_Operator_out2296_out1 <= in492 XOR in496;

  Logical_Operator_out2297_out1 <= Logical_Operator_out1273_out1 XOR Logical_Operator_out1275_out1;

  Logical_Operator_out2298_out1 <= Logical_Operator_out1274_out1 XOR Logical_Operator_out1276_out1;

  Logical_Operator_out2299_out1 <= Logical_Operator_out250_out1 XOR Logical_Operator_out252_out1;

  Logical_Operator_out2300_out1 <= in500 XOR in504;

  Logical_Operator_out2301_out1 <= Logical_Operator_out1277_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out2302_out1 <= Logical_Operator_out1278_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out2303_out1 <= Logical_Operator_out254_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out2304_out1 <= in508 XOR in512;

  Logical_Operator_out2305_out1 <= Logical_Operator_out1281_out1 XOR Logical_Operator_out1283_out1;

  Logical_Operator_out2306_out1 <= Logical_Operator_out1282_out1 XOR Logical_Operator_out1284_out1;

  Logical_Operator_out2307_out1 <= Logical_Operator_out258_out1 XOR Logical_Operator_out260_out1;

  Logical_Operator_out2308_out1 <= in516 XOR in520;

  Logical_Operator_out2309_out1 <= Logical_Operator_out1285_out1 XOR Logical_Operator_out1287_out1;

  Logical_Operator_out2310_out1 <= Logical_Operator_out1286_out1 XOR Logical_Operator_out1288_out1;

  Logical_Operator_out2311_out1 <= Logical_Operator_out262_out1 XOR Logical_Operator_out264_out1;

  Logical_Operator_out2312_out1 <= in524 XOR in528;

  Logical_Operator_out2313_out1 <= Logical_Operator_out1289_out1 XOR Logical_Operator_out1291_out1;

  Logical_Operator_out2314_out1 <= Logical_Operator_out1290_out1 XOR Logical_Operator_out1292_out1;

  Logical_Operator_out2315_out1 <= Logical_Operator_out266_out1 XOR Logical_Operator_out268_out1;

  Logical_Operator_out2316_out1 <= in532 XOR in536;

  Logical_Operator_out2317_out1 <= Logical_Operator_out1293_out1 XOR Logical_Operator_out1295_out1;

  Logical_Operator_out2318_out1 <= Logical_Operator_out1294_out1 XOR Logical_Operator_out1296_out1;

  Logical_Operator_out2319_out1 <= Logical_Operator_out270_out1 XOR Logical_Operator_out272_out1;

  Logical_Operator_out2320_out1 <= in540 XOR in544;

  Logical_Operator_out2321_out1 <= Logical_Operator_out1297_out1 XOR Logical_Operator_out1299_out1;

  Logical_Operator_out2322_out1 <= Logical_Operator_out1298_out1 XOR Logical_Operator_out1300_out1;

  Logical_Operator_out2323_out1 <= Logical_Operator_out274_out1 XOR Logical_Operator_out276_out1;

  Logical_Operator_out2324_out1 <= in548 XOR in552;

  Logical_Operator_out2325_out1 <= Logical_Operator_out1301_out1 XOR Logical_Operator_out1303_out1;

  Logical_Operator_out2326_out1 <= Logical_Operator_out1302_out1 XOR Logical_Operator_out1304_out1;

  Logical_Operator_out2327_out1 <= Logical_Operator_out278_out1 XOR Logical_Operator_out280_out1;

  Logical_Operator_out2328_out1 <= in556 XOR in560;

  Logical_Operator_out2329_out1 <= Logical_Operator_out1305_out1 XOR Logical_Operator_out1307_out1;

  Logical_Operator_out2330_out1 <= Logical_Operator_out1306_out1 XOR Logical_Operator_out1308_out1;

  Logical_Operator_out2331_out1 <= Logical_Operator_out282_out1 XOR Logical_Operator_out284_out1;

  Logical_Operator_out2332_out1 <= in564 XOR in568;

  Logical_Operator_out2333_out1 <= Logical_Operator_out1309_out1 XOR Logical_Operator_out1311_out1;

  Logical_Operator_out2334_out1 <= Logical_Operator_out1310_out1 XOR Logical_Operator_out1312_out1;

  Logical_Operator_out2335_out1 <= Logical_Operator_out286_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out2336_out1 <= in572 XOR in576;

  Logical_Operator_out2337_out1 <= Logical_Operator_out1313_out1 XOR Logical_Operator_out1315_out1;

  Logical_Operator_out2338_out1 <= Logical_Operator_out1314_out1 XOR Logical_Operator_out1316_out1;

  Logical_Operator_out2339_out1 <= Logical_Operator_out290_out1 XOR Logical_Operator_out292_out1;

  Logical_Operator_out2340_out1 <= in580 XOR in584;

  Logical_Operator_out2341_out1 <= Logical_Operator_out1317_out1 XOR Logical_Operator_out1319_out1;

  Logical_Operator_out2342_out1 <= Logical_Operator_out1318_out1 XOR Logical_Operator_out1320_out1;

  Logical_Operator_out2343_out1 <= Logical_Operator_out294_out1 XOR Logical_Operator_out296_out1;

  Logical_Operator_out2344_out1 <= in588 XOR in592;

  Logical_Operator_out2345_out1 <= Logical_Operator_out1321_out1 XOR Logical_Operator_out1323_out1;

  Logical_Operator_out2346_out1 <= Logical_Operator_out1322_out1 XOR Logical_Operator_out1324_out1;

  Logical_Operator_out2347_out1 <= Logical_Operator_out298_out1 XOR Logical_Operator_out300_out1;

  Logical_Operator_out2348_out1 <= in596 XOR in600;

  Logical_Operator_out2349_out1 <= Logical_Operator_out1325_out1 XOR Logical_Operator_out1327_out1;

  Logical_Operator_out2350_out1 <= Logical_Operator_out1326_out1 XOR Logical_Operator_out1328_out1;

  Logical_Operator_out2351_out1 <= Logical_Operator_out302_out1 XOR Logical_Operator_out304_out1;

  Logical_Operator_out2352_out1 <= in604 XOR in608;

  Logical_Operator_out2353_out1 <= Logical_Operator_out1329_out1 XOR Logical_Operator_out1331_out1;

  Logical_Operator_out2354_out1 <= Logical_Operator_out1330_out1 XOR Logical_Operator_out1332_out1;

  Logical_Operator_out2355_out1 <= Logical_Operator_out306_out1 XOR Logical_Operator_out308_out1;

  Logical_Operator_out2356_out1 <= in612 XOR in616;

  Logical_Operator_out2357_out1 <= Logical_Operator_out1333_out1 XOR Logical_Operator_out1335_out1;

  Logical_Operator_out2358_out1 <= Logical_Operator_out1334_out1 XOR Logical_Operator_out1336_out1;

  Logical_Operator_out2359_out1 <= Logical_Operator_out310_out1 XOR Logical_Operator_out312_out1;

  Logical_Operator_out2360_out1 <= in620 XOR in624;

  Logical_Operator_out2361_out1 <= Logical_Operator_out1337_out1 XOR Logical_Operator_out1339_out1;

  Logical_Operator_out2362_out1 <= Logical_Operator_out1338_out1 XOR Logical_Operator_out1340_out1;

  Logical_Operator_out2363_out1 <= Logical_Operator_out314_out1 XOR Logical_Operator_out316_out1;

  Logical_Operator_out2364_out1 <= in628 XOR in632;

  Logical_Operator_out2365_out1 <= Logical_Operator_out1341_out1 XOR Logical_Operator_out1343_out1;

  Logical_Operator_out2366_out1 <= Logical_Operator_out1342_out1 XOR Logical_Operator_out1344_out1;

  Logical_Operator_out2367_out1 <= Logical_Operator_out318_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out2368_out1 <= in636 XOR in640;

  Logical_Operator_out2369_out1 <= Logical_Operator_out1345_out1 XOR Logical_Operator_out1347_out1;

  Logical_Operator_out2370_out1 <= Logical_Operator_out1346_out1 XOR Logical_Operator_out1348_out1;

  Logical_Operator_out2371_out1 <= Logical_Operator_out322_out1 XOR Logical_Operator_out324_out1;

  Logical_Operator_out2372_out1 <= in644 XOR in648;

  Logical_Operator_out2373_out1 <= Logical_Operator_out1349_out1 XOR Logical_Operator_out1351_out1;

  Logical_Operator_out2374_out1 <= Logical_Operator_out1350_out1 XOR Logical_Operator_out1352_out1;

  Logical_Operator_out2375_out1 <= Logical_Operator_out326_out1 XOR Logical_Operator_out328_out1;

  Logical_Operator_out2376_out1 <= in652 XOR in656;

  Logical_Operator_out2377_out1 <= Logical_Operator_out1353_out1 XOR Logical_Operator_out1355_out1;

  Logical_Operator_out2378_out1 <= Logical_Operator_out1354_out1 XOR Logical_Operator_out1356_out1;

  Logical_Operator_out2379_out1 <= Logical_Operator_out330_out1 XOR Logical_Operator_out332_out1;

  Logical_Operator_out2380_out1 <= in660 XOR in664;

  Logical_Operator_out2381_out1 <= Logical_Operator_out1357_out1 XOR Logical_Operator_out1359_out1;

  Logical_Operator_out2382_out1 <= Logical_Operator_out1358_out1 XOR Logical_Operator_out1360_out1;

  Logical_Operator_out2383_out1 <= Logical_Operator_out334_out1 XOR Logical_Operator_out336_out1;

  Logical_Operator_out2384_out1 <= in668 XOR in672;

  Logical_Operator_out2385_out1 <= Logical_Operator_out1361_out1 XOR Logical_Operator_out1363_out1;

  Logical_Operator_out2386_out1 <= Logical_Operator_out1362_out1 XOR Logical_Operator_out1364_out1;

  Logical_Operator_out2387_out1 <= Logical_Operator_out338_out1 XOR Logical_Operator_out340_out1;

  Logical_Operator_out2388_out1 <= in676 XOR in680;

  Logical_Operator_out2389_out1 <= Logical_Operator_out1365_out1 XOR Logical_Operator_out1367_out1;

  Logical_Operator_out2390_out1 <= Logical_Operator_out1366_out1 XOR Logical_Operator_out1368_out1;

  Logical_Operator_out2391_out1 <= Logical_Operator_out342_out1 XOR Logical_Operator_out344_out1;

  Logical_Operator_out2392_out1 <= in684 XOR in688;

  Logical_Operator_out2393_out1 <= Logical_Operator_out1369_out1 XOR Logical_Operator_out1371_out1;

  Logical_Operator_out2394_out1 <= Logical_Operator_out1370_out1 XOR Logical_Operator_out1372_out1;

  Logical_Operator_out2395_out1 <= Logical_Operator_out346_out1 XOR Logical_Operator_out348_out1;

  Logical_Operator_out2396_out1 <= in692 XOR in696;

  Logical_Operator_out2397_out1 <= Logical_Operator_out1373_out1 XOR Logical_Operator_out1375_out1;

  Logical_Operator_out2398_out1 <= Logical_Operator_out1374_out1 XOR Logical_Operator_out1376_out1;

  Logical_Operator_out2399_out1 <= Logical_Operator_out350_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out2400_out1 <= in700 XOR in704;

  Logical_Operator_out2401_out1 <= Logical_Operator_out1377_out1 XOR Logical_Operator_out1379_out1;

  Logical_Operator_out2402_out1 <= Logical_Operator_out1378_out1 XOR Logical_Operator_out1380_out1;

  Logical_Operator_out2403_out1 <= Logical_Operator_out354_out1 XOR Logical_Operator_out356_out1;

  Logical_Operator_out2404_out1 <= in708 XOR in712;

  Logical_Operator_out2405_out1 <= Logical_Operator_out1381_out1 XOR Logical_Operator_out1383_out1;

  Logical_Operator_out2406_out1 <= Logical_Operator_out1382_out1 XOR Logical_Operator_out1384_out1;

  Logical_Operator_out2407_out1 <= Logical_Operator_out358_out1 XOR Logical_Operator_out360_out1;

  Logical_Operator_out2408_out1 <= in716 XOR in720;

  Logical_Operator_out2409_out1 <= Logical_Operator_out1385_out1 XOR Logical_Operator_out1387_out1;

  Logical_Operator_out2410_out1 <= Logical_Operator_out1386_out1 XOR Logical_Operator_out1388_out1;

  Logical_Operator_out2411_out1 <= Logical_Operator_out362_out1 XOR Logical_Operator_out364_out1;

  Logical_Operator_out2412_out1 <= in724 XOR in728;

  Logical_Operator_out2413_out1 <= Logical_Operator_out1389_out1 XOR Logical_Operator_out1391_out1;

  Logical_Operator_out2414_out1 <= Logical_Operator_out1390_out1 XOR Logical_Operator_out1392_out1;

  Logical_Operator_out2415_out1 <= Logical_Operator_out366_out1 XOR Logical_Operator_out368_out1;

  Logical_Operator_out2416_out1 <= in732 XOR in736;

  Logical_Operator_out2417_out1 <= Logical_Operator_out1393_out1 XOR Logical_Operator_out1395_out1;

  Logical_Operator_out2418_out1 <= Logical_Operator_out1394_out1 XOR Logical_Operator_out1396_out1;

  Logical_Operator_out2419_out1 <= Logical_Operator_out370_out1 XOR Logical_Operator_out372_out1;

  Logical_Operator_out2420_out1 <= in740 XOR in744;

  Logical_Operator_out2421_out1 <= Logical_Operator_out1397_out1 XOR Logical_Operator_out1399_out1;

  Logical_Operator_out2422_out1 <= Logical_Operator_out1398_out1 XOR Logical_Operator_out1400_out1;

  Logical_Operator_out2423_out1 <= Logical_Operator_out374_out1 XOR Logical_Operator_out376_out1;

  Logical_Operator_out2424_out1 <= in748 XOR in752;

  Logical_Operator_out2425_out1 <= Logical_Operator_out1401_out1 XOR Logical_Operator_out1403_out1;

  Logical_Operator_out2426_out1 <= Logical_Operator_out1402_out1 XOR Logical_Operator_out1404_out1;

  Logical_Operator_out2427_out1 <= Logical_Operator_out378_out1 XOR Logical_Operator_out380_out1;

  Logical_Operator_out2428_out1 <= in756 XOR in760;

  Logical_Operator_out2429_out1 <= Logical_Operator_out1405_out1 XOR Logical_Operator_out1407_out1;

  Logical_Operator_out2430_out1 <= Logical_Operator_out1406_out1 XOR Logical_Operator_out1408_out1;

  Logical_Operator_out2431_out1 <= Logical_Operator_out382_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out2432_out1 <= in764 XOR in768;

  Logical_Operator_out2433_out1 <= Logical_Operator_out1409_out1 XOR Logical_Operator_out1411_out1;

  Logical_Operator_out2434_out1 <= Logical_Operator_out1410_out1 XOR Logical_Operator_out1412_out1;

  Logical_Operator_out2435_out1 <= Logical_Operator_out386_out1 XOR Logical_Operator_out388_out1;

  Logical_Operator_out2436_out1 <= in772 XOR in776;

  Logical_Operator_out2437_out1 <= Logical_Operator_out1413_out1 XOR Logical_Operator_out1415_out1;

  Logical_Operator_out2438_out1 <= Logical_Operator_out1414_out1 XOR Logical_Operator_out1416_out1;

  Logical_Operator_out2439_out1 <= Logical_Operator_out390_out1 XOR Logical_Operator_out392_out1;

  Logical_Operator_out2440_out1 <= in780 XOR in784;

  Logical_Operator_out2441_out1 <= Logical_Operator_out1417_out1 XOR Logical_Operator_out1419_out1;

  Logical_Operator_out2442_out1 <= Logical_Operator_out1418_out1 XOR Logical_Operator_out1420_out1;

  Logical_Operator_out2443_out1 <= Logical_Operator_out394_out1 XOR Logical_Operator_out396_out1;

  Logical_Operator_out2444_out1 <= in788 XOR in792;

  Logical_Operator_out2445_out1 <= Logical_Operator_out1421_out1 XOR Logical_Operator_out1423_out1;

  Logical_Operator_out2446_out1 <= Logical_Operator_out1422_out1 XOR Logical_Operator_out1424_out1;

  Logical_Operator_out2447_out1 <= Logical_Operator_out398_out1 XOR Logical_Operator_out400_out1;

  Logical_Operator_out2448_out1 <= in796 XOR in800;

  Logical_Operator_out2449_out1 <= Logical_Operator_out1425_out1 XOR Logical_Operator_out1427_out1;

  Logical_Operator_out2450_out1 <= Logical_Operator_out1426_out1 XOR Logical_Operator_out1428_out1;

  Logical_Operator_out2451_out1 <= Logical_Operator_out402_out1 XOR Logical_Operator_out404_out1;

  Logical_Operator_out2452_out1 <= in804 XOR in808;

  Logical_Operator_out2453_out1 <= Logical_Operator_out1429_out1 XOR Logical_Operator_out1431_out1;

  Logical_Operator_out2454_out1 <= Logical_Operator_out1430_out1 XOR Logical_Operator_out1432_out1;

  Logical_Operator_out2455_out1 <= Logical_Operator_out406_out1 XOR Logical_Operator_out408_out1;

  Logical_Operator_out2456_out1 <= in812 XOR in816;

  Logical_Operator_out2457_out1 <= Logical_Operator_out1433_out1 XOR Logical_Operator_out1435_out1;

  Logical_Operator_out2458_out1 <= Logical_Operator_out1434_out1 XOR Logical_Operator_out1436_out1;

  Logical_Operator_out2459_out1 <= Logical_Operator_out410_out1 XOR Logical_Operator_out412_out1;

  Logical_Operator_out2460_out1 <= in820 XOR in824;

  Logical_Operator_out2461_out1 <= Logical_Operator_out1437_out1 XOR Logical_Operator_out1439_out1;

  Logical_Operator_out2462_out1 <= Logical_Operator_out1438_out1 XOR Logical_Operator_out1440_out1;

  Logical_Operator_out2463_out1 <= Logical_Operator_out414_out1 XOR Logical_Operator_out416_out1;

  Logical_Operator_out2464_out1 <= in828 XOR in832;

  Logical_Operator_out2465_out1 <= Logical_Operator_out1441_out1 XOR Logical_Operator_out1443_out1;

  Logical_Operator_out2466_out1 <= Logical_Operator_out1442_out1 XOR Logical_Operator_out1444_out1;

  Logical_Operator_out2467_out1 <= Logical_Operator_out418_out1 XOR Logical_Operator_out420_out1;

  Logical_Operator_out2468_out1 <= in836 XOR in840;

  Logical_Operator_out2469_out1 <= Logical_Operator_out1445_out1 XOR Logical_Operator_out1447_out1;

  Logical_Operator_out2470_out1 <= Logical_Operator_out1446_out1 XOR Logical_Operator_out1448_out1;

  Logical_Operator_out2471_out1 <= Logical_Operator_out422_out1 XOR Logical_Operator_out424_out1;

  Logical_Operator_out2472_out1 <= in844 XOR in848;

  Logical_Operator_out2473_out1 <= Logical_Operator_out1449_out1 XOR Logical_Operator_out1451_out1;

  Logical_Operator_out2474_out1 <= Logical_Operator_out1450_out1 XOR Logical_Operator_out1452_out1;

  Logical_Operator_out2475_out1 <= Logical_Operator_out426_out1 XOR Logical_Operator_out428_out1;

  Logical_Operator_out2476_out1 <= in852 XOR in856;

  Logical_Operator_out2477_out1 <= Logical_Operator_out1453_out1 XOR Logical_Operator_out1455_out1;

  Logical_Operator_out2478_out1 <= Logical_Operator_out1454_out1 XOR Logical_Operator_out1456_out1;

  Logical_Operator_out2479_out1 <= Logical_Operator_out430_out1 XOR Logical_Operator_out432_out1;

  Logical_Operator_out2480_out1 <= in860 XOR in864;

  Logical_Operator_out2481_out1 <= Logical_Operator_out1457_out1 XOR Logical_Operator_out1459_out1;

  Logical_Operator_out2482_out1 <= Logical_Operator_out1458_out1 XOR Logical_Operator_out1460_out1;

  Logical_Operator_out2483_out1 <= Logical_Operator_out434_out1 XOR Logical_Operator_out436_out1;

  Logical_Operator_out2484_out1 <= in868 XOR in872;

  Logical_Operator_out2485_out1 <= Logical_Operator_out1461_out1 XOR Logical_Operator_out1463_out1;

  Logical_Operator_out2486_out1 <= Logical_Operator_out1462_out1 XOR Logical_Operator_out1464_out1;

  Logical_Operator_out2487_out1 <= Logical_Operator_out438_out1 XOR Logical_Operator_out440_out1;

  Logical_Operator_out2488_out1 <= in876 XOR in880;

  Logical_Operator_out2489_out1 <= Logical_Operator_out1465_out1 XOR Logical_Operator_out1467_out1;

  Logical_Operator_out2490_out1 <= Logical_Operator_out1466_out1 XOR Logical_Operator_out1468_out1;

  Logical_Operator_out2491_out1 <= Logical_Operator_out442_out1 XOR Logical_Operator_out444_out1;

  Logical_Operator_out2492_out1 <= in884 XOR in888;

  Logical_Operator_out2493_out1 <= Logical_Operator_out1469_out1 XOR Logical_Operator_out1471_out1;

  Logical_Operator_out2494_out1 <= Logical_Operator_out1470_out1 XOR Logical_Operator_out1472_out1;

  Logical_Operator_out2495_out1 <= Logical_Operator_out446_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out2496_out1 <= in892 XOR in896;

  Logical_Operator_out2497_out1 <= Logical_Operator_out1473_out1 XOR Logical_Operator_out1475_out1;

  Logical_Operator_out2498_out1 <= Logical_Operator_out1474_out1 XOR Logical_Operator_out1476_out1;

  Logical_Operator_out2499_out1 <= Logical_Operator_out450_out1 XOR Logical_Operator_out452_out1;

  Logical_Operator_out2500_out1 <= in900 XOR in904;

  Logical_Operator_out2501_out1 <= Logical_Operator_out1477_out1 XOR Logical_Operator_out1479_out1;

  Logical_Operator_out2502_out1 <= Logical_Operator_out1478_out1 XOR Logical_Operator_out1480_out1;

  Logical_Operator_out2503_out1 <= Logical_Operator_out454_out1 XOR Logical_Operator_out456_out1;

  Logical_Operator_out2504_out1 <= in908 XOR in912;

  Logical_Operator_out2505_out1 <= Logical_Operator_out1481_out1 XOR Logical_Operator_out1483_out1;

  Logical_Operator_out2506_out1 <= Logical_Operator_out1482_out1 XOR Logical_Operator_out1484_out1;

  Logical_Operator_out2507_out1 <= Logical_Operator_out458_out1 XOR Logical_Operator_out460_out1;

  Logical_Operator_out2508_out1 <= in916 XOR in920;

  Logical_Operator_out2509_out1 <= Logical_Operator_out1485_out1 XOR Logical_Operator_out1487_out1;

  Logical_Operator_out2510_out1 <= Logical_Operator_out1486_out1 XOR Logical_Operator_out1488_out1;

  Logical_Operator_out2511_out1 <= Logical_Operator_out462_out1 XOR Logical_Operator_out464_out1;

  Logical_Operator_out2512_out1 <= in924 XOR in928;

  Logical_Operator_out2513_out1 <= Logical_Operator_out1489_out1 XOR Logical_Operator_out1491_out1;

  Logical_Operator_out2514_out1 <= Logical_Operator_out1490_out1 XOR Logical_Operator_out1492_out1;

  Logical_Operator_out2515_out1 <= Logical_Operator_out466_out1 XOR Logical_Operator_out468_out1;

  Logical_Operator_out2516_out1 <= in932 XOR in936;

  Logical_Operator_out2517_out1 <= Logical_Operator_out1493_out1 XOR Logical_Operator_out1495_out1;

  Logical_Operator_out2518_out1 <= Logical_Operator_out1494_out1 XOR Logical_Operator_out1496_out1;

  Logical_Operator_out2519_out1 <= Logical_Operator_out470_out1 XOR Logical_Operator_out472_out1;

  Logical_Operator_out2520_out1 <= in940 XOR in944;

  Logical_Operator_out2521_out1 <= Logical_Operator_out1497_out1 XOR Logical_Operator_out1499_out1;

  Logical_Operator_out2522_out1 <= Logical_Operator_out1498_out1 XOR Logical_Operator_out1500_out1;

  Logical_Operator_out2523_out1 <= Logical_Operator_out474_out1 XOR Logical_Operator_out476_out1;

  Logical_Operator_out2524_out1 <= in948 XOR in952;

  Logical_Operator_out2525_out1 <= Logical_Operator_out1501_out1 XOR Logical_Operator_out1503_out1;

  Logical_Operator_out2526_out1 <= Logical_Operator_out1502_out1 XOR Logical_Operator_out1504_out1;

  Logical_Operator_out2527_out1 <= Logical_Operator_out478_out1 XOR Logical_Operator_out480_out1;

  Logical_Operator_out2528_out1 <= in956 XOR in960;

  Logical_Operator_out2529_out1 <= Logical_Operator_out1505_out1 XOR Logical_Operator_out1507_out1;

  Logical_Operator_out2530_out1 <= Logical_Operator_out1506_out1 XOR Logical_Operator_out1508_out1;

  Logical_Operator_out2531_out1 <= Logical_Operator_out482_out1 XOR Logical_Operator_out484_out1;

  Logical_Operator_out2532_out1 <= in964 XOR in968;

  Logical_Operator_out2533_out1 <= Logical_Operator_out1509_out1 XOR Logical_Operator_out1511_out1;

  Logical_Operator_out2534_out1 <= Logical_Operator_out1510_out1 XOR Logical_Operator_out1512_out1;

  Logical_Operator_out2535_out1 <= Logical_Operator_out486_out1 XOR Logical_Operator_out488_out1;

  Logical_Operator_out2536_out1 <= in972 XOR in976;

  Logical_Operator_out2537_out1 <= Logical_Operator_out1513_out1 XOR Logical_Operator_out1515_out1;

  Logical_Operator_out2538_out1 <= Logical_Operator_out1514_out1 XOR Logical_Operator_out1516_out1;

  Logical_Operator_out2539_out1 <= Logical_Operator_out490_out1 XOR Logical_Operator_out492_out1;

  Logical_Operator_out2540_out1 <= in980 XOR in984;

  Logical_Operator_out2541_out1 <= Logical_Operator_out1517_out1 XOR Logical_Operator_out1519_out1;

  Logical_Operator_out2542_out1 <= Logical_Operator_out1518_out1 XOR Logical_Operator_out1520_out1;

  Logical_Operator_out2543_out1 <= Logical_Operator_out494_out1 XOR Logical_Operator_out496_out1;

  Logical_Operator_out2544_out1 <= in988 XOR in992;

  Logical_Operator_out2545_out1 <= Logical_Operator_out1521_out1 XOR Logical_Operator_out1523_out1;

  Logical_Operator_out2546_out1 <= Logical_Operator_out1522_out1 XOR Logical_Operator_out1524_out1;

  Logical_Operator_out2547_out1 <= Logical_Operator_out498_out1 XOR Logical_Operator_out500_out1;

  Logical_Operator_out2548_out1 <= in996 XOR in1000;

  Logical_Operator_out2549_out1 <= Logical_Operator_out1525_out1 XOR Logical_Operator_out1527_out1;

  Logical_Operator_out2550_out1 <= Logical_Operator_out1526_out1 XOR Logical_Operator_out1528_out1;

  Logical_Operator_out2551_out1 <= Logical_Operator_out502_out1 XOR Logical_Operator_out504_out1;

  Logical_Operator_out2552_out1 <= in1004 XOR in1008;

  Logical_Operator_out2553_out1 <= Logical_Operator_out1529_out1 XOR Logical_Operator_out1531_out1;

  Logical_Operator_out2554_out1 <= Logical_Operator_out1530_out1 XOR Logical_Operator_out1532_out1;

  Logical_Operator_out2555_out1 <= Logical_Operator_out506_out1 XOR Logical_Operator_out508_out1;

  Logical_Operator_out2556_out1 <= in1012 XOR in1016;

  Logical_Operator_out2557_out1 <= Logical_Operator_out1533_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out2558_out1 <= Logical_Operator_out1534_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out2559_out1 <= Logical_Operator_out510_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out2560_out1 <= in1020 XOR in1024;

  Logical_Operator_out2561_out1 <= Logical_Operator_out1537_out1 XOR Logical_Operator_out1539_out1;

  Logical_Operator_out2562_out1 <= Logical_Operator_out1538_out1 XOR Logical_Operator_out1540_out1;

  Logical_Operator_out2563_out1 <= Logical_Operator_out514_out1 XOR Logical_Operator_out516_out1;

  Logical_Operator_out2564_out1 <= in1028 XOR in1032;

  Logical_Operator_out2565_out1 <= Logical_Operator_out1541_out1 XOR Logical_Operator_out1543_out1;

  Logical_Operator_out2566_out1 <= Logical_Operator_out1542_out1 XOR Logical_Operator_out1544_out1;

  Logical_Operator_out2567_out1 <= Logical_Operator_out518_out1 XOR Logical_Operator_out520_out1;

  Logical_Operator_out2568_out1 <= in1036 XOR in1040;

  Logical_Operator_out2569_out1 <= Logical_Operator_out1545_out1 XOR Logical_Operator_out1547_out1;

  Logical_Operator_out2570_out1 <= Logical_Operator_out1546_out1 XOR Logical_Operator_out1548_out1;

  Logical_Operator_out2571_out1 <= Logical_Operator_out522_out1 XOR Logical_Operator_out524_out1;

  Logical_Operator_out2572_out1 <= in1044 XOR in1048;

  Logical_Operator_out2573_out1 <= Logical_Operator_out1549_out1 XOR Logical_Operator_out1551_out1;

  Logical_Operator_out2574_out1 <= Logical_Operator_out1550_out1 XOR Logical_Operator_out1552_out1;

  Logical_Operator_out2575_out1 <= Logical_Operator_out526_out1 XOR Logical_Operator_out528_out1;

  Logical_Operator_out2576_out1 <= in1052 XOR in1056;

  Logical_Operator_out2577_out1 <= Logical_Operator_out1553_out1 XOR Logical_Operator_out1555_out1;

  Logical_Operator_out2578_out1 <= Logical_Operator_out1554_out1 XOR Logical_Operator_out1556_out1;

  Logical_Operator_out2579_out1 <= Logical_Operator_out530_out1 XOR Logical_Operator_out532_out1;

  Logical_Operator_out2580_out1 <= in1060 XOR in1064;

  Logical_Operator_out2581_out1 <= Logical_Operator_out1557_out1 XOR Logical_Operator_out1559_out1;

  Logical_Operator_out2582_out1 <= Logical_Operator_out1558_out1 XOR Logical_Operator_out1560_out1;

  Logical_Operator_out2583_out1 <= Logical_Operator_out534_out1 XOR Logical_Operator_out536_out1;

  Logical_Operator_out2584_out1 <= in1068 XOR in1072;

  Logical_Operator_out2585_out1 <= Logical_Operator_out1561_out1 XOR Logical_Operator_out1563_out1;

  Logical_Operator_out2586_out1 <= Logical_Operator_out1562_out1 XOR Logical_Operator_out1564_out1;

  Logical_Operator_out2587_out1 <= Logical_Operator_out538_out1 XOR Logical_Operator_out540_out1;

  Logical_Operator_out2588_out1 <= in1076 XOR in1080;

  Logical_Operator_out2589_out1 <= Logical_Operator_out1565_out1 XOR Logical_Operator_out1567_out1;

  Logical_Operator_out2590_out1 <= Logical_Operator_out1566_out1 XOR Logical_Operator_out1568_out1;

  Logical_Operator_out2591_out1 <= Logical_Operator_out542_out1 XOR Logical_Operator_out544_out1;

  Logical_Operator_out2592_out1 <= in1084 XOR in1088;

  Logical_Operator_out2593_out1 <= Logical_Operator_out1569_out1 XOR Logical_Operator_out1571_out1;

  Logical_Operator_out2594_out1 <= Logical_Operator_out1570_out1 XOR Logical_Operator_out1572_out1;

  Logical_Operator_out2595_out1 <= Logical_Operator_out546_out1 XOR Logical_Operator_out548_out1;

  Logical_Operator_out2596_out1 <= in1092 XOR in1096;

  Logical_Operator_out2597_out1 <= Logical_Operator_out1573_out1 XOR Logical_Operator_out1575_out1;

  Logical_Operator_out2598_out1 <= Logical_Operator_out1574_out1 XOR Logical_Operator_out1576_out1;

  Logical_Operator_out2599_out1 <= Logical_Operator_out550_out1 XOR Logical_Operator_out552_out1;

  Logical_Operator_out2600_out1 <= in1100 XOR in1104;

  Logical_Operator_out2601_out1 <= Logical_Operator_out1577_out1 XOR Logical_Operator_out1579_out1;

  Logical_Operator_out2602_out1 <= Logical_Operator_out1578_out1 XOR Logical_Operator_out1580_out1;

  Logical_Operator_out2603_out1 <= Logical_Operator_out554_out1 XOR Logical_Operator_out556_out1;

  Logical_Operator_out2604_out1 <= in1108 XOR in1112;

  Logical_Operator_out2605_out1 <= Logical_Operator_out1581_out1 XOR Logical_Operator_out1583_out1;

  Logical_Operator_out2606_out1 <= Logical_Operator_out1582_out1 XOR Logical_Operator_out1584_out1;

  Logical_Operator_out2607_out1 <= Logical_Operator_out558_out1 XOR Logical_Operator_out560_out1;

  Logical_Operator_out2608_out1 <= in1116 XOR in1120;

  Logical_Operator_out2609_out1 <= Logical_Operator_out1585_out1 XOR Logical_Operator_out1587_out1;

  Logical_Operator_out2610_out1 <= Logical_Operator_out1586_out1 XOR Logical_Operator_out1588_out1;

  Logical_Operator_out2611_out1 <= Logical_Operator_out562_out1 XOR Logical_Operator_out564_out1;

  Logical_Operator_out2612_out1 <= in1124 XOR in1128;

  Logical_Operator_out2613_out1 <= Logical_Operator_out1589_out1 XOR Logical_Operator_out1591_out1;

  Logical_Operator_out2614_out1 <= Logical_Operator_out1590_out1 XOR Logical_Operator_out1592_out1;

  Logical_Operator_out2615_out1 <= Logical_Operator_out566_out1 XOR Logical_Operator_out568_out1;

  Logical_Operator_out2616_out1 <= in1132 XOR in1136;

  Logical_Operator_out2617_out1 <= Logical_Operator_out1593_out1 XOR Logical_Operator_out1595_out1;

  Logical_Operator_out2618_out1 <= Logical_Operator_out1594_out1 XOR Logical_Operator_out1596_out1;

  Logical_Operator_out2619_out1 <= Logical_Operator_out570_out1 XOR Logical_Operator_out572_out1;

  Logical_Operator_out2620_out1 <= in1140 XOR in1144;

  Logical_Operator_out2621_out1 <= Logical_Operator_out1597_out1 XOR Logical_Operator_out1599_out1;

  Logical_Operator_out2622_out1 <= Logical_Operator_out1598_out1 XOR Logical_Operator_out1600_out1;

  Logical_Operator_out2623_out1 <= Logical_Operator_out574_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out2624_out1 <= in1148 XOR in1152;

  Logical_Operator_out2625_out1 <= Logical_Operator_out1601_out1 XOR Logical_Operator_out1603_out1;

  Logical_Operator_out2626_out1 <= Logical_Operator_out1602_out1 XOR Logical_Operator_out1604_out1;

  Logical_Operator_out2627_out1 <= Logical_Operator_out578_out1 XOR Logical_Operator_out580_out1;

  Logical_Operator_out2628_out1 <= in1156 XOR in1160;

  Logical_Operator_out2629_out1 <= Logical_Operator_out1605_out1 XOR Logical_Operator_out1607_out1;

  Logical_Operator_out2630_out1 <= Logical_Operator_out1606_out1 XOR Logical_Operator_out1608_out1;

  Logical_Operator_out2631_out1 <= Logical_Operator_out582_out1 XOR Logical_Operator_out584_out1;

  Logical_Operator_out2632_out1 <= in1164 XOR in1168;

  Logical_Operator_out2633_out1 <= Logical_Operator_out1609_out1 XOR Logical_Operator_out1611_out1;

  Logical_Operator_out2634_out1 <= Logical_Operator_out1610_out1 XOR Logical_Operator_out1612_out1;

  Logical_Operator_out2635_out1 <= Logical_Operator_out586_out1 XOR Logical_Operator_out588_out1;

  Logical_Operator_out2636_out1 <= in1172 XOR in1176;

  Logical_Operator_out2637_out1 <= Logical_Operator_out1613_out1 XOR Logical_Operator_out1615_out1;

  Logical_Operator_out2638_out1 <= Logical_Operator_out1614_out1 XOR Logical_Operator_out1616_out1;

  Logical_Operator_out2639_out1 <= Logical_Operator_out590_out1 XOR Logical_Operator_out592_out1;

  Logical_Operator_out2640_out1 <= in1180 XOR in1184;

  Logical_Operator_out2641_out1 <= Logical_Operator_out1617_out1 XOR Logical_Operator_out1619_out1;

  Logical_Operator_out2642_out1 <= Logical_Operator_out1618_out1 XOR Logical_Operator_out1620_out1;

  Logical_Operator_out2643_out1 <= Logical_Operator_out594_out1 XOR Logical_Operator_out596_out1;

  Logical_Operator_out2644_out1 <= in1188 XOR in1192;

  Logical_Operator_out2645_out1 <= Logical_Operator_out1621_out1 XOR Logical_Operator_out1623_out1;

  Logical_Operator_out2646_out1 <= Logical_Operator_out1622_out1 XOR Logical_Operator_out1624_out1;

  Logical_Operator_out2647_out1 <= Logical_Operator_out598_out1 XOR Logical_Operator_out600_out1;

  Logical_Operator_out2648_out1 <= in1196 XOR in1200;

  Logical_Operator_out2649_out1 <= Logical_Operator_out1625_out1 XOR Logical_Operator_out1627_out1;

  Logical_Operator_out2650_out1 <= Logical_Operator_out1626_out1 XOR Logical_Operator_out1628_out1;

  Logical_Operator_out2651_out1 <= Logical_Operator_out602_out1 XOR Logical_Operator_out604_out1;

  Logical_Operator_out2652_out1 <= in1204 XOR in1208;

  Logical_Operator_out2653_out1 <= Logical_Operator_out1629_out1 XOR Logical_Operator_out1631_out1;

  Logical_Operator_out2654_out1 <= Logical_Operator_out1630_out1 XOR Logical_Operator_out1632_out1;

  Logical_Operator_out2655_out1 <= Logical_Operator_out606_out1 XOR Logical_Operator_out608_out1;

  Logical_Operator_out2656_out1 <= in1212 XOR in1216;

  Logical_Operator_out2657_out1 <= Logical_Operator_out1633_out1 XOR Logical_Operator_out1635_out1;

  Logical_Operator_out2658_out1 <= Logical_Operator_out1634_out1 XOR Logical_Operator_out1636_out1;

  Logical_Operator_out2659_out1 <= Logical_Operator_out610_out1 XOR Logical_Operator_out612_out1;

  Logical_Operator_out2660_out1 <= in1220 XOR in1224;

  Logical_Operator_out2661_out1 <= Logical_Operator_out1637_out1 XOR Logical_Operator_out1639_out1;

  Logical_Operator_out2662_out1 <= Logical_Operator_out1638_out1 XOR Logical_Operator_out1640_out1;

  Logical_Operator_out2663_out1 <= Logical_Operator_out614_out1 XOR Logical_Operator_out616_out1;

  Logical_Operator_out2664_out1 <= in1228 XOR in1232;

  Logical_Operator_out2665_out1 <= Logical_Operator_out1641_out1 XOR Logical_Operator_out1643_out1;

  Logical_Operator_out2666_out1 <= Logical_Operator_out1642_out1 XOR Logical_Operator_out1644_out1;

  Logical_Operator_out2667_out1 <= Logical_Operator_out618_out1 XOR Logical_Operator_out620_out1;

  Logical_Operator_out2668_out1 <= in1236 XOR in1240;

  Logical_Operator_out2669_out1 <= Logical_Operator_out1645_out1 XOR Logical_Operator_out1647_out1;

  Logical_Operator_out2670_out1 <= Logical_Operator_out1646_out1 XOR Logical_Operator_out1648_out1;

  Logical_Operator_out2671_out1 <= Logical_Operator_out622_out1 XOR Logical_Operator_out624_out1;

  Logical_Operator_out2672_out1 <= in1244 XOR in1248;

  Logical_Operator_out2673_out1 <= Logical_Operator_out1649_out1 XOR Logical_Operator_out1651_out1;

  Logical_Operator_out2674_out1 <= Logical_Operator_out1650_out1 XOR Logical_Operator_out1652_out1;

  Logical_Operator_out2675_out1 <= Logical_Operator_out626_out1 XOR Logical_Operator_out628_out1;

  Logical_Operator_out2676_out1 <= in1252 XOR in1256;

  Logical_Operator_out2677_out1 <= Logical_Operator_out1653_out1 XOR Logical_Operator_out1655_out1;

  Logical_Operator_out2678_out1 <= Logical_Operator_out1654_out1 XOR Logical_Operator_out1656_out1;

  Logical_Operator_out2679_out1 <= Logical_Operator_out630_out1 XOR Logical_Operator_out632_out1;

  Logical_Operator_out2680_out1 <= in1260 XOR in1264;

  Logical_Operator_out2681_out1 <= Logical_Operator_out1657_out1 XOR Logical_Operator_out1659_out1;

  Logical_Operator_out2682_out1 <= Logical_Operator_out1658_out1 XOR Logical_Operator_out1660_out1;

  Logical_Operator_out2683_out1 <= Logical_Operator_out634_out1 XOR Logical_Operator_out636_out1;

  Logical_Operator_out2684_out1 <= in1268 XOR in1272;

  Logical_Operator_out2685_out1 <= Logical_Operator_out1661_out1 XOR Logical_Operator_out1663_out1;

  Logical_Operator_out2686_out1 <= Logical_Operator_out1662_out1 XOR Logical_Operator_out1664_out1;

  Logical_Operator_out2687_out1 <= Logical_Operator_out638_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out2688_out1 <= in1276 XOR in1280;

  Logical_Operator_out2689_out1 <= Logical_Operator_out1665_out1 XOR Logical_Operator_out1667_out1;

  Logical_Operator_out2690_out1 <= Logical_Operator_out1666_out1 XOR Logical_Operator_out1668_out1;

  Logical_Operator_out2691_out1 <= Logical_Operator_out642_out1 XOR Logical_Operator_out644_out1;

  Logical_Operator_out2692_out1 <= in1284 XOR in1288;

  Logical_Operator_out2693_out1 <= Logical_Operator_out1669_out1 XOR Logical_Operator_out1671_out1;

  Logical_Operator_out2694_out1 <= Logical_Operator_out1670_out1 XOR Logical_Operator_out1672_out1;

  Logical_Operator_out2695_out1 <= Logical_Operator_out646_out1 XOR Logical_Operator_out648_out1;

  Logical_Operator_out2696_out1 <= in1292 XOR in1296;

  Logical_Operator_out2697_out1 <= Logical_Operator_out1673_out1 XOR Logical_Operator_out1675_out1;

  Logical_Operator_out2698_out1 <= Logical_Operator_out1674_out1 XOR Logical_Operator_out1676_out1;

  Logical_Operator_out2699_out1 <= Logical_Operator_out650_out1 XOR Logical_Operator_out652_out1;

  Logical_Operator_out2700_out1 <= in1300 XOR in1304;

  Logical_Operator_out2701_out1 <= Logical_Operator_out1677_out1 XOR Logical_Operator_out1679_out1;

  Logical_Operator_out2702_out1 <= Logical_Operator_out1678_out1 XOR Logical_Operator_out1680_out1;

  Logical_Operator_out2703_out1 <= Logical_Operator_out654_out1 XOR Logical_Operator_out656_out1;

  Logical_Operator_out2704_out1 <= in1308 XOR in1312;

  Logical_Operator_out2705_out1 <= Logical_Operator_out1681_out1 XOR Logical_Operator_out1683_out1;

  Logical_Operator_out2706_out1 <= Logical_Operator_out1682_out1 XOR Logical_Operator_out1684_out1;

  Logical_Operator_out2707_out1 <= Logical_Operator_out658_out1 XOR Logical_Operator_out660_out1;

  Logical_Operator_out2708_out1 <= in1316 XOR in1320;

  Logical_Operator_out2709_out1 <= Logical_Operator_out1685_out1 XOR Logical_Operator_out1687_out1;

  Logical_Operator_out2710_out1 <= Logical_Operator_out1686_out1 XOR Logical_Operator_out1688_out1;

  Logical_Operator_out2711_out1 <= Logical_Operator_out662_out1 XOR Logical_Operator_out664_out1;

  Logical_Operator_out2712_out1 <= in1324 XOR in1328;

  Logical_Operator_out2713_out1 <= Logical_Operator_out1689_out1 XOR Logical_Operator_out1691_out1;

  Logical_Operator_out2714_out1 <= Logical_Operator_out1690_out1 XOR Logical_Operator_out1692_out1;

  Logical_Operator_out2715_out1 <= Logical_Operator_out666_out1 XOR Logical_Operator_out668_out1;

  Logical_Operator_out2716_out1 <= in1332 XOR in1336;

  Logical_Operator_out2717_out1 <= Logical_Operator_out1693_out1 XOR Logical_Operator_out1695_out1;

  Logical_Operator_out2718_out1 <= Logical_Operator_out1694_out1 XOR Logical_Operator_out1696_out1;

  Logical_Operator_out2719_out1 <= Logical_Operator_out670_out1 XOR Logical_Operator_out672_out1;

  Logical_Operator_out2720_out1 <= in1340 XOR in1344;

  Logical_Operator_out2721_out1 <= Logical_Operator_out1697_out1 XOR Logical_Operator_out1699_out1;

  Logical_Operator_out2722_out1 <= Logical_Operator_out1698_out1 XOR Logical_Operator_out1700_out1;

  Logical_Operator_out2723_out1 <= Logical_Operator_out674_out1 XOR Logical_Operator_out676_out1;

  Logical_Operator_out2724_out1 <= in1348 XOR in1352;

  Logical_Operator_out2725_out1 <= Logical_Operator_out1701_out1 XOR Logical_Operator_out1703_out1;

  Logical_Operator_out2726_out1 <= Logical_Operator_out1702_out1 XOR Logical_Operator_out1704_out1;

  Logical_Operator_out2727_out1 <= Logical_Operator_out678_out1 XOR Logical_Operator_out680_out1;

  Logical_Operator_out2728_out1 <= in1356 XOR in1360;

  Logical_Operator_out2729_out1 <= Logical_Operator_out1705_out1 XOR Logical_Operator_out1707_out1;

  Logical_Operator_out2730_out1 <= Logical_Operator_out1706_out1 XOR Logical_Operator_out1708_out1;

  Logical_Operator_out2731_out1 <= Logical_Operator_out682_out1 XOR Logical_Operator_out684_out1;

  Logical_Operator_out2732_out1 <= in1364 XOR in1368;

  Logical_Operator_out2733_out1 <= Logical_Operator_out1709_out1 XOR Logical_Operator_out1711_out1;

  Logical_Operator_out2734_out1 <= Logical_Operator_out1710_out1 XOR Logical_Operator_out1712_out1;

  Logical_Operator_out2735_out1 <= Logical_Operator_out686_out1 XOR Logical_Operator_out688_out1;

  Logical_Operator_out2736_out1 <= in1372 XOR in1376;

  Logical_Operator_out2737_out1 <= Logical_Operator_out1713_out1 XOR Logical_Operator_out1715_out1;

  Logical_Operator_out2738_out1 <= Logical_Operator_out1714_out1 XOR Logical_Operator_out1716_out1;

  Logical_Operator_out2739_out1 <= Logical_Operator_out690_out1 XOR Logical_Operator_out692_out1;

  Logical_Operator_out2740_out1 <= in1380 XOR in1384;

  Logical_Operator_out2741_out1 <= Logical_Operator_out1717_out1 XOR Logical_Operator_out1719_out1;

  Logical_Operator_out2742_out1 <= Logical_Operator_out1718_out1 XOR Logical_Operator_out1720_out1;

  Logical_Operator_out2743_out1 <= Logical_Operator_out694_out1 XOR Logical_Operator_out696_out1;

  Logical_Operator_out2744_out1 <= in1388 XOR in1392;

  Logical_Operator_out2745_out1 <= Logical_Operator_out1721_out1 XOR Logical_Operator_out1723_out1;

  Logical_Operator_out2746_out1 <= Logical_Operator_out1722_out1 XOR Logical_Operator_out1724_out1;

  Logical_Operator_out2747_out1 <= Logical_Operator_out698_out1 XOR Logical_Operator_out700_out1;

  Logical_Operator_out2748_out1 <= in1396 XOR in1400;

  Logical_Operator_out2749_out1 <= Logical_Operator_out1725_out1 XOR Logical_Operator_out1727_out1;

  Logical_Operator_out2750_out1 <= Logical_Operator_out1726_out1 XOR Logical_Operator_out1728_out1;

  Logical_Operator_out2751_out1 <= Logical_Operator_out702_out1 XOR Logical_Operator_out704_out1;

  Logical_Operator_out2752_out1 <= in1404 XOR in1408;

  Logical_Operator_out2753_out1 <= Logical_Operator_out1729_out1 XOR Logical_Operator_out1731_out1;

  Logical_Operator_out2754_out1 <= Logical_Operator_out1730_out1 XOR Logical_Operator_out1732_out1;

  Logical_Operator_out2755_out1 <= Logical_Operator_out706_out1 XOR Logical_Operator_out708_out1;

  Logical_Operator_out2756_out1 <= in1412 XOR in1416;

  Logical_Operator_out2757_out1 <= Logical_Operator_out1733_out1 XOR Logical_Operator_out1735_out1;

  Logical_Operator_out2758_out1 <= Logical_Operator_out1734_out1 XOR Logical_Operator_out1736_out1;

  Logical_Operator_out2759_out1 <= Logical_Operator_out710_out1 XOR Logical_Operator_out712_out1;

  Logical_Operator_out2760_out1 <= in1420 XOR in1424;

  Logical_Operator_out2761_out1 <= Logical_Operator_out1737_out1 XOR Logical_Operator_out1739_out1;

  Logical_Operator_out2762_out1 <= Logical_Operator_out1738_out1 XOR Logical_Operator_out1740_out1;

  Logical_Operator_out2763_out1 <= Logical_Operator_out714_out1 XOR Logical_Operator_out716_out1;

  Logical_Operator_out2764_out1 <= in1428 XOR in1432;

  Logical_Operator_out2765_out1 <= Logical_Operator_out1741_out1 XOR Logical_Operator_out1743_out1;

  Logical_Operator_out2766_out1 <= Logical_Operator_out1742_out1 XOR Logical_Operator_out1744_out1;

  Logical_Operator_out2767_out1 <= Logical_Operator_out718_out1 XOR Logical_Operator_out720_out1;

  Logical_Operator_out2768_out1 <= in1436 XOR in1440;

  Logical_Operator_out2769_out1 <= Logical_Operator_out1745_out1 XOR Logical_Operator_out1747_out1;

  Logical_Operator_out2770_out1 <= Logical_Operator_out1746_out1 XOR Logical_Operator_out1748_out1;

  Logical_Operator_out2771_out1 <= Logical_Operator_out722_out1 XOR Logical_Operator_out724_out1;

  Logical_Operator_out2772_out1 <= in1444 XOR in1448;

  Logical_Operator_out2773_out1 <= Logical_Operator_out1749_out1 XOR Logical_Operator_out1751_out1;

  Logical_Operator_out2774_out1 <= Logical_Operator_out1750_out1 XOR Logical_Operator_out1752_out1;

  Logical_Operator_out2775_out1 <= Logical_Operator_out726_out1 XOR Logical_Operator_out728_out1;

  Logical_Operator_out2776_out1 <= in1452 XOR in1456;

  Logical_Operator_out2777_out1 <= Logical_Operator_out1753_out1 XOR Logical_Operator_out1755_out1;

  Logical_Operator_out2778_out1 <= Logical_Operator_out1754_out1 XOR Logical_Operator_out1756_out1;

  Logical_Operator_out2779_out1 <= Logical_Operator_out730_out1 XOR Logical_Operator_out732_out1;

  Logical_Operator_out2780_out1 <= in1460 XOR in1464;

  Logical_Operator_out2781_out1 <= Logical_Operator_out1757_out1 XOR Logical_Operator_out1759_out1;

  Logical_Operator_out2782_out1 <= Logical_Operator_out1758_out1 XOR Logical_Operator_out1760_out1;

  Logical_Operator_out2783_out1 <= Logical_Operator_out734_out1 XOR Logical_Operator_out736_out1;

  Logical_Operator_out2784_out1 <= in1468 XOR in1472;

  Logical_Operator_out2785_out1 <= Logical_Operator_out1761_out1 XOR Logical_Operator_out1763_out1;

  Logical_Operator_out2786_out1 <= Logical_Operator_out1762_out1 XOR Logical_Operator_out1764_out1;

  Logical_Operator_out2787_out1 <= Logical_Operator_out738_out1 XOR Logical_Operator_out740_out1;

  Logical_Operator_out2788_out1 <= in1476 XOR in1480;

  Logical_Operator_out2789_out1 <= Logical_Operator_out1765_out1 XOR Logical_Operator_out1767_out1;

  Logical_Operator_out2790_out1 <= Logical_Operator_out1766_out1 XOR Logical_Operator_out1768_out1;

  Logical_Operator_out2791_out1 <= Logical_Operator_out742_out1 XOR Logical_Operator_out744_out1;

  Logical_Operator_out2792_out1 <= in1484 XOR in1488;

  Logical_Operator_out2793_out1 <= Logical_Operator_out1769_out1 XOR Logical_Operator_out1771_out1;

  Logical_Operator_out2794_out1 <= Logical_Operator_out1770_out1 XOR Logical_Operator_out1772_out1;

  Logical_Operator_out2795_out1 <= Logical_Operator_out746_out1 XOR Logical_Operator_out748_out1;

  Logical_Operator_out2796_out1 <= in1492 XOR in1496;

  Logical_Operator_out2797_out1 <= Logical_Operator_out1773_out1 XOR Logical_Operator_out1775_out1;

  Logical_Operator_out2798_out1 <= Logical_Operator_out1774_out1 XOR Logical_Operator_out1776_out1;

  Logical_Operator_out2799_out1 <= Logical_Operator_out750_out1 XOR Logical_Operator_out752_out1;

  Logical_Operator_out2800_out1 <= in1500 XOR in1504;

  Logical_Operator_out2801_out1 <= Logical_Operator_out1777_out1 XOR Logical_Operator_out1779_out1;

  Logical_Operator_out2802_out1 <= Logical_Operator_out1778_out1 XOR Logical_Operator_out1780_out1;

  Logical_Operator_out2803_out1 <= Logical_Operator_out754_out1 XOR Logical_Operator_out756_out1;

  Logical_Operator_out2804_out1 <= in1508 XOR in1512;

  Logical_Operator_out2805_out1 <= Logical_Operator_out1781_out1 XOR Logical_Operator_out1783_out1;

  Logical_Operator_out2806_out1 <= Logical_Operator_out1782_out1 XOR Logical_Operator_out1784_out1;

  Logical_Operator_out2807_out1 <= Logical_Operator_out758_out1 XOR Logical_Operator_out760_out1;

  Logical_Operator_out2808_out1 <= in1516 XOR in1520;

  Logical_Operator_out2809_out1 <= Logical_Operator_out1785_out1 XOR Logical_Operator_out1787_out1;

  Logical_Operator_out2810_out1 <= Logical_Operator_out1786_out1 XOR Logical_Operator_out1788_out1;

  Logical_Operator_out2811_out1 <= Logical_Operator_out762_out1 XOR Logical_Operator_out764_out1;

  Logical_Operator_out2812_out1 <= in1524 XOR in1528;

  Logical_Operator_out2813_out1 <= Logical_Operator_out1789_out1 XOR Logical_Operator_out1791_out1;

  Logical_Operator_out2814_out1 <= Logical_Operator_out1790_out1 XOR Logical_Operator_out1792_out1;

  Logical_Operator_out2815_out1 <= Logical_Operator_out766_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out2816_out1 <= in1532 XOR in1536;

  Logical_Operator_out2817_out1 <= Logical_Operator_out1793_out1 XOR Logical_Operator_out1795_out1;

  Logical_Operator_out2818_out1 <= Logical_Operator_out1794_out1 XOR Logical_Operator_out1796_out1;

  Logical_Operator_out2819_out1 <= Logical_Operator_out770_out1 XOR Logical_Operator_out772_out1;

  Logical_Operator_out2820_out1 <= in1540 XOR in1544;

  Logical_Operator_out2821_out1 <= Logical_Operator_out1797_out1 XOR Logical_Operator_out1799_out1;

  Logical_Operator_out2822_out1 <= Logical_Operator_out1798_out1 XOR Logical_Operator_out1800_out1;

  Logical_Operator_out2823_out1 <= Logical_Operator_out774_out1 XOR Logical_Operator_out776_out1;

  Logical_Operator_out2824_out1 <= in1548 XOR in1552;

  Logical_Operator_out2825_out1 <= Logical_Operator_out1801_out1 XOR Logical_Operator_out1803_out1;

  Logical_Operator_out2826_out1 <= Logical_Operator_out1802_out1 XOR Logical_Operator_out1804_out1;

  Logical_Operator_out2827_out1 <= Logical_Operator_out778_out1 XOR Logical_Operator_out780_out1;

  Logical_Operator_out2828_out1 <= in1556 XOR in1560;

  Logical_Operator_out2829_out1 <= Logical_Operator_out1805_out1 XOR Logical_Operator_out1807_out1;

  Logical_Operator_out2830_out1 <= Logical_Operator_out1806_out1 XOR Logical_Operator_out1808_out1;

  Logical_Operator_out2831_out1 <= Logical_Operator_out782_out1 XOR Logical_Operator_out784_out1;

  Logical_Operator_out2832_out1 <= in1564 XOR in1568;

  Logical_Operator_out2833_out1 <= Logical_Operator_out1809_out1 XOR Logical_Operator_out1811_out1;

  Logical_Operator_out2834_out1 <= Logical_Operator_out1810_out1 XOR Logical_Operator_out1812_out1;

  Logical_Operator_out2835_out1 <= Logical_Operator_out786_out1 XOR Logical_Operator_out788_out1;

  Logical_Operator_out2836_out1 <= in1572 XOR in1576;

  Logical_Operator_out2837_out1 <= Logical_Operator_out1813_out1 XOR Logical_Operator_out1815_out1;

  Logical_Operator_out2838_out1 <= Logical_Operator_out1814_out1 XOR Logical_Operator_out1816_out1;

  Logical_Operator_out2839_out1 <= Logical_Operator_out790_out1 XOR Logical_Operator_out792_out1;

  Logical_Operator_out2840_out1 <= in1580 XOR in1584;

  Logical_Operator_out2841_out1 <= Logical_Operator_out1817_out1 XOR Logical_Operator_out1819_out1;

  Logical_Operator_out2842_out1 <= Logical_Operator_out1818_out1 XOR Logical_Operator_out1820_out1;

  Logical_Operator_out2843_out1 <= Logical_Operator_out794_out1 XOR Logical_Operator_out796_out1;

  Logical_Operator_out2844_out1 <= in1588 XOR in1592;

  Logical_Operator_out2845_out1 <= Logical_Operator_out1821_out1 XOR Logical_Operator_out1823_out1;

  Logical_Operator_out2846_out1 <= Logical_Operator_out1822_out1 XOR Logical_Operator_out1824_out1;

  Logical_Operator_out2847_out1 <= Logical_Operator_out798_out1 XOR Logical_Operator_out800_out1;

  Logical_Operator_out2848_out1 <= in1596 XOR in1600;

  Logical_Operator_out2849_out1 <= Logical_Operator_out1825_out1 XOR Logical_Operator_out1827_out1;

  Logical_Operator_out2850_out1 <= Logical_Operator_out1826_out1 XOR Logical_Operator_out1828_out1;

  Logical_Operator_out2851_out1 <= Logical_Operator_out802_out1 XOR Logical_Operator_out804_out1;

  Logical_Operator_out2852_out1 <= in1604 XOR in1608;

  Logical_Operator_out2853_out1 <= Logical_Operator_out1829_out1 XOR Logical_Operator_out1831_out1;

  Logical_Operator_out2854_out1 <= Logical_Operator_out1830_out1 XOR Logical_Operator_out1832_out1;

  Logical_Operator_out2855_out1 <= Logical_Operator_out806_out1 XOR Logical_Operator_out808_out1;

  Logical_Operator_out2856_out1 <= in1612 XOR in1616;

  Logical_Operator_out2857_out1 <= Logical_Operator_out1833_out1 XOR Logical_Operator_out1835_out1;

  Logical_Operator_out2858_out1 <= Logical_Operator_out1834_out1 XOR Logical_Operator_out1836_out1;

  Logical_Operator_out2859_out1 <= Logical_Operator_out810_out1 XOR Logical_Operator_out812_out1;

  Logical_Operator_out2860_out1 <= in1620 XOR in1624;

  Logical_Operator_out2861_out1 <= Logical_Operator_out1837_out1 XOR Logical_Operator_out1839_out1;

  Logical_Operator_out2862_out1 <= Logical_Operator_out1838_out1 XOR Logical_Operator_out1840_out1;

  Logical_Operator_out2863_out1 <= Logical_Operator_out814_out1 XOR Logical_Operator_out816_out1;

  Logical_Operator_out2864_out1 <= in1628 XOR in1632;

  Logical_Operator_out2865_out1 <= Logical_Operator_out1841_out1 XOR Logical_Operator_out1843_out1;

  Logical_Operator_out2866_out1 <= Logical_Operator_out1842_out1 XOR Logical_Operator_out1844_out1;

  Logical_Operator_out2867_out1 <= Logical_Operator_out818_out1 XOR Logical_Operator_out820_out1;

  Logical_Operator_out2868_out1 <= in1636 XOR in1640;

  Logical_Operator_out2869_out1 <= Logical_Operator_out1845_out1 XOR Logical_Operator_out1847_out1;

  Logical_Operator_out2870_out1 <= Logical_Operator_out1846_out1 XOR Logical_Operator_out1848_out1;

  Logical_Operator_out2871_out1 <= Logical_Operator_out822_out1 XOR Logical_Operator_out824_out1;

  Logical_Operator_out2872_out1 <= in1644 XOR in1648;

  Logical_Operator_out2873_out1 <= Logical_Operator_out1849_out1 XOR Logical_Operator_out1851_out1;

  Logical_Operator_out2874_out1 <= Logical_Operator_out1850_out1 XOR Logical_Operator_out1852_out1;

  Logical_Operator_out2875_out1 <= Logical_Operator_out826_out1 XOR Logical_Operator_out828_out1;

  Logical_Operator_out2876_out1 <= in1652 XOR in1656;

  Logical_Operator_out2877_out1 <= Logical_Operator_out1853_out1 XOR Logical_Operator_out1855_out1;

  Logical_Operator_out2878_out1 <= Logical_Operator_out1854_out1 XOR Logical_Operator_out1856_out1;

  Logical_Operator_out2879_out1 <= Logical_Operator_out830_out1 XOR Logical_Operator_out832_out1;

  Logical_Operator_out2880_out1 <= in1660 XOR in1664;

  Logical_Operator_out2881_out1 <= Logical_Operator_out1857_out1 XOR Logical_Operator_out1859_out1;

  Logical_Operator_out2882_out1 <= Logical_Operator_out1858_out1 XOR Logical_Operator_out1860_out1;

  Logical_Operator_out2883_out1 <= Logical_Operator_out834_out1 XOR Logical_Operator_out836_out1;

  Logical_Operator_out2884_out1 <= in1668 XOR in1672;

  Logical_Operator_out2885_out1 <= Logical_Operator_out1861_out1 XOR Logical_Operator_out1863_out1;

  Logical_Operator_out2886_out1 <= Logical_Operator_out1862_out1 XOR Logical_Operator_out1864_out1;

  Logical_Operator_out2887_out1 <= Logical_Operator_out838_out1 XOR Logical_Operator_out840_out1;

  Logical_Operator_out2888_out1 <= in1676 XOR in1680;

  Logical_Operator_out2889_out1 <= Logical_Operator_out1865_out1 XOR Logical_Operator_out1867_out1;

  Logical_Operator_out2890_out1 <= Logical_Operator_out1866_out1 XOR Logical_Operator_out1868_out1;

  Logical_Operator_out2891_out1 <= Logical_Operator_out842_out1 XOR Logical_Operator_out844_out1;

  Logical_Operator_out2892_out1 <= in1684 XOR in1688;

  Logical_Operator_out2893_out1 <= Logical_Operator_out1869_out1 XOR Logical_Operator_out1871_out1;

  Logical_Operator_out2894_out1 <= Logical_Operator_out1870_out1 XOR Logical_Operator_out1872_out1;

  Logical_Operator_out2895_out1 <= Logical_Operator_out846_out1 XOR Logical_Operator_out848_out1;

  Logical_Operator_out2896_out1 <= in1692 XOR in1696;

  Logical_Operator_out2897_out1 <= Logical_Operator_out1873_out1 XOR Logical_Operator_out1875_out1;

  Logical_Operator_out2898_out1 <= Logical_Operator_out1874_out1 XOR Logical_Operator_out1876_out1;

  Logical_Operator_out2899_out1 <= Logical_Operator_out850_out1 XOR Logical_Operator_out852_out1;

  Logical_Operator_out2900_out1 <= in1700 XOR in1704;

  Logical_Operator_out2901_out1 <= Logical_Operator_out1877_out1 XOR Logical_Operator_out1879_out1;

  Logical_Operator_out2902_out1 <= Logical_Operator_out1878_out1 XOR Logical_Operator_out1880_out1;

  Logical_Operator_out2903_out1 <= Logical_Operator_out854_out1 XOR Logical_Operator_out856_out1;

  Logical_Operator_out2904_out1 <= in1708 XOR in1712;

  Logical_Operator_out2905_out1 <= Logical_Operator_out1881_out1 XOR Logical_Operator_out1883_out1;

  Logical_Operator_out2906_out1 <= Logical_Operator_out1882_out1 XOR Logical_Operator_out1884_out1;

  Logical_Operator_out2907_out1 <= Logical_Operator_out858_out1 XOR Logical_Operator_out860_out1;

  Logical_Operator_out2908_out1 <= in1716 XOR in1720;

  Logical_Operator_out2909_out1 <= Logical_Operator_out1885_out1 XOR Logical_Operator_out1887_out1;

  Logical_Operator_out2910_out1 <= Logical_Operator_out1886_out1 XOR Logical_Operator_out1888_out1;

  Logical_Operator_out2911_out1 <= Logical_Operator_out862_out1 XOR Logical_Operator_out864_out1;

  Logical_Operator_out2912_out1 <= in1724 XOR in1728;

  Logical_Operator_out2913_out1 <= Logical_Operator_out1889_out1 XOR Logical_Operator_out1891_out1;

  Logical_Operator_out2914_out1 <= Logical_Operator_out1890_out1 XOR Logical_Operator_out1892_out1;

  Logical_Operator_out2915_out1 <= Logical_Operator_out866_out1 XOR Logical_Operator_out868_out1;

  Logical_Operator_out2916_out1 <= in1732 XOR in1736;

  Logical_Operator_out2917_out1 <= Logical_Operator_out1893_out1 XOR Logical_Operator_out1895_out1;

  Logical_Operator_out2918_out1 <= Logical_Operator_out1894_out1 XOR Logical_Operator_out1896_out1;

  Logical_Operator_out2919_out1 <= Logical_Operator_out870_out1 XOR Logical_Operator_out872_out1;

  Logical_Operator_out2920_out1 <= in1740 XOR in1744;

  Logical_Operator_out2921_out1 <= Logical_Operator_out1897_out1 XOR Logical_Operator_out1899_out1;

  Logical_Operator_out2922_out1 <= Logical_Operator_out1898_out1 XOR Logical_Operator_out1900_out1;

  Logical_Operator_out2923_out1 <= Logical_Operator_out874_out1 XOR Logical_Operator_out876_out1;

  Logical_Operator_out2924_out1 <= in1748 XOR in1752;

  Logical_Operator_out2925_out1 <= Logical_Operator_out1901_out1 XOR Logical_Operator_out1903_out1;

  Logical_Operator_out2926_out1 <= Logical_Operator_out1902_out1 XOR Logical_Operator_out1904_out1;

  Logical_Operator_out2927_out1 <= Logical_Operator_out878_out1 XOR Logical_Operator_out880_out1;

  Logical_Operator_out2928_out1 <= in1756 XOR in1760;

  Logical_Operator_out2929_out1 <= Logical_Operator_out1905_out1 XOR Logical_Operator_out1907_out1;

  Logical_Operator_out2930_out1 <= Logical_Operator_out1906_out1 XOR Logical_Operator_out1908_out1;

  Logical_Operator_out2931_out1 <= Logical_Operator_out882_out1 XOR Logical_Operator_out884_out1;

  Logical_Operator_out2932_out1 <= in1764 XOR in1768;

  Logical_Operator_out2933_out1 <= Logical_Operator_out1909_out1 XOR Logical_Operator_out1911_out1;

  Logical_Operator_out2934_out1 <= Logical_Operator_out1910_out1 XOR Logical_Operator_out1912_out1;

  Logical_Operator_out2935_out1 <= Logical_Operator_out886_out1 XOR Logical_Operator_out888_out1;

  Logical_Operator_out2936_out1 <= in1772 XOR in1776;

  Logical_Operator_out2937_out1 <= Logical_Operator_out1913_out1 XOR Logical_Operator_out1915_out1;

  Logical_Operator_out2938_out1 <= Logical_Operator_out1914_out1 XOR Logical_Operator_out1916_out1;

  Logical_Operator_out2939_out1 <= Logical_Operator_out890_out1 XOR Logical_Operator_out892_out1;

  Logical_Operator_out2940_out1 <= in1780 XOR in1784;

  Logical_Operator_out2941_out1 <= Logical_Operator_out1917_out1 XOR Logical_Operator_out1919_out1;

  Logical_Operator_out2942_out1 <= Logical_Operator_out1918_out1 XOR Logical_Operator_out1920_out1;

  Logical_Operator_out2943_out1 <= Logical_Operator_out894_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out2944_out1 <= in1788 XOR in1792;

  Logical_Operator_out2945_out1 <= Logical_Operator_out1921_out1 XOR Logical_Operator_out1923_out1;

  Logical_Operator_out2946_out1 <= Logical_Operator_out1922_out1 XOR Logical_Operator_out1924_out1;

  Logical_Operator_out2947_out1 <= Logical_Operator_out898_out1 XOR Logical_Operator_out900_out1;

  Logical_Operator_out2948_out1 <= in1796 XOR in1800;

  Logical_Operator_out2949_out1 <= Logical_Operator_out1925_out1 XOR Logical_Operator_out1927_out1;

  Logical_Operator_out2950_out1 <= Logical_Operator_out1926_out1 XOR Logical_Operator_out1928_out1;

  Logical_Operator_out2951_out1 <= Logical_Operator_out902_out1 XOR Logical_Operator_out904_out1;

  Logical_Operator_out2952_out1 <= in1804 XOR in1808;

  Logical_Operator_out2953_out1 <= Logical_Operator_out1929_out1 XOR Logical_Operator_out1931_out1;

  Logical_Operator_out2954_out1 <= Logical_Operator_out1930_out1 XOR Logical_Operator_out1932_out1;

  Logical_Operator_out2955_out1 <= Logical_Operator_out906_out1 XOR Logical_Operator_out908_out1;

  Logical_Operator_out2956_out1 <= in1812 XOR in1816;

  Logical_Operator_out2957_out1 <= Logical_Operator_out1933_out1 XOR Logical_Operator_out1935_out1;

  Logical_Operator_out2958_out1 <= Logical_Operator_out1934_out1 XOR Logical_Operator_out1936_out1;

  Logical_Operator_out2959_out1 <= Logical_Operator_out910_out1 XOR Logical_Operator_out912_out1;

  Logical_Operator_out2960_out1 <= in1820 XOR in1824;

  Logical_Operator_out2961_out1 <= Logical_Operator_out1937_out1 XOR Logical_Operator_out1939_out1;

  Logical_Operator_out2962_out1 <= Logical_Operator_out1938_out1 XOR Logical_Operator_out1940_out1;

  Logical_Operator_out2963_out1 <= Logical_Operator_out914_out1 XOR Logical_Operator_out916_out1;

  Logical_Operator_out2964_out1 <= in1828 XOR in1832;

  Logical_Operator_out2965_out1 <= Logical_Operator_out1941_out1 XOR Logical_Operator_out1943_out1;

  Logical_Operator_out2966_out1 <= Logical_Operator_out1942_out1 XOR Logical_Operator_out1944_out1;

  Logical_Operator_out2967_out1 <= Logical_Operator_out918_out1 XOR Logical_Operator_out920_out1;

  Logical_Operator_out2968_out1 <= in1836 XOR in1840;

  Logical_Operator_out2969_out1 <= Logical_Operator_out1945_out1 XOR Logical_Operator_out1947_out1;

  Logical_Operator_out2970_out1 <= Logical_Operator_out1946_out1 XOR Logical_Operator_out1948_out1;

  Logical_Operator_out2971_out1 <= Logical_Operator_out922_out1 XOR Logical_Operator_out924_out1;

  Logical_Operator_out2972_out1 <= in1844 XOR in1848;

  Logical_Operator_out2973_out1 <= Logical_Operator_out1949_out1 XOR Logical_Operator_out1951_out1;

  Logical_Operator_out2974_out1 <= Logical_Operator_out1950_out1 XOR Logical_Operator_out1952_out1;

  Logical_Operator_out2975_out1 <= Logical_Operator_out926_out1 XOR Logical_Operator_out928_out1;

  Logical_Operator_out2976_out1 <= in1852 XOR in1856;

  Logical_Operator_out2977_out1 <= Logical_Operator_out1953_out1 XOR Logical_Operator_out1955_out1;

  Logical_Operator_out2978_out1 <= Logical_Operator_out1954_out1 XOR Logical_Operator_out1956_out1;

  Logical_Operator_out2979_out1 <= Logical_Operator_out930_out1 XOR Logical_Operator_out932_out1;

  Logical_Operator_out2980_out1 <= in1860 XOR in1864;

  Logical_Operator_out2981_out1 <= Logical_Operator_out1957_out1 XOR Logical_Operator_out1959_out1;

  Logical_Operator_out2982_out1 <= Logical_Operator_out1958_out1 XOR Logical_Operator_out1960_out1;

  Logical_Operator_out2983_out1 <= Logical_Operator_out934_out1 XOR Logical_Operator_out936_out1;

  Logical_Operator_out2984_out1 <= in1868 XOR in1872;

  Logical_Operator_out2985_out1 <= Logical_Operator_out1961_out1 XOR Logical_Operator_out1963_out1;

  Logical_Operator_out2986_out1 <= Logical_Operator_out1962_out1 XOR Logical_Operator_out1964_out1;

  Logical_Operator_out2987_out1 <= Logical_Operator_out938_out1 XOR Logical_Operator_out940_out1;

  Logical_Operator_out2988_out1 <= in1876 XOR in1880;

  Logical_Operator_out2989_out1 <= Logical_Operator_out1965_out1 XOR Logical_Operator_out1967_out1;

  Logical_Operator_out2990_out1 <= Logical_Operator_out1966_out1 XOR Logical_Operator_out1968_out1;

  Logical_Operator_out2991_out1 <= Logical_Operator_out942_out1 XOR Logical_Operator_out944_out1;

  Logical_Operator_out2992_out1 <= in1884 XOR in1888;

  Logical_Operator_out2993_out1 <= Logical_Operator_out1969_out1 XOR Logical_Operator_out1971_out1;

  Logical_Operator_out2994_out1 <= Logical_Operator_out1970_out1 XOR Logical_Operator_out1972_out1;

  Logical_Operator_out2995_out1 <= Logical_Operator_out946_out1 XOR Logical_Operator_out948_out1;

  Logical_Operator_out2996_out1 <= in1892 XOR in1896;

  Logical_Operator_out2997_out1 <= Logical_Operator_out1973_out1 XOR Logical_Operator_out1975_out1;

  Logical_Operator_out2998_out1 <= Logical_Operator_out1974_out1 XOR Logical_Operator_out1976_out1;

  Logical_Operator_out2999_out1 <= Logical_Operator_out950_out1 XOR Logical_Operator_out952_out1;

  Logical_Operator_out3000_out1 <= in1900 XOR in1904;

  Logical_Operator_out3001_out1 <= Logical_Operator_out1977_out1 XOR Logical_Operator_out1979_out1;

  Logical_Operator_out3002_out1 <= Logical_Operator_out1978_out1 XOR Logical_Operator_out1980_out1;

  Logical_Operator_out3003_out1 <= Logical_Operator_out954_out1 XOR Logical_Operator_out956_out1;

  Logical_Operator_out3004_out1 <= in1908 XOR in1912;

  Logical_Operator_out3005_out1 <= Logical_Operator_out1981_out1 XOR Logical_Operator_out1983_out1;

  Logical_Operator_out3006_out1 <= Logical_Operator_out1982_out1 XOR Logical_Operator_out1984_out1;

  Logical_Operator_out3007_out1 <= Logical_Operator_out958_out1 XOR Logical_Operator_out960_out1;

  Logical_Operator_out3008_out1 <= in1916 XOR in1920;

  Logical_Operator_out3009_out1 <= Logical_Operator_out1985_out1 XOR Logical_Operator_out1987_out1;

  Logical_Operator_out3010_out1 <= Logical_Operator_out1986_out1 XOR Logical_Operator_out1988_out1;

  Logical_Operator_out3011_out1 <= Logical_Operator_out962_out1 XOR Logical_Operator_out964_out1;

  Logical_Operator_out3012_out1 <= in1924 XOR in1928;

  Logical_Operator_out3013_out1 <= Logical_Operator_out1989_out1 XOR Logical_Operator_out1991_out1;

  Logical_Operator_out3014_out1 <= Logical_Operator_out1990_out1 XOR Logical_Operator_out1992_out1;

  Logical_Operator_out3015_out1 <= Logical_Operator_out966_out1 XOR Logical_Operator_out968_out1;

  Logical_Operator_out3016_out1 <= in1932 XOR in1936;

  Logical_Operator_out3017_out1 <= Logical_Operator_out1993_out1 XOR Logical_Operator_out1995_out1;

  Logical_Operator_out3018_out1 <= Logical_Operator_out1994_out1 XOR Logical_Operator_out1996_out1;

  Logical_Operator_out3019_out1 <= Logical_Operator_out970_out1 XOR Logical_Operator_out972_out1;

  Logical_Operator_out3020_out1 <= in1940 XOR in1944;

  Logical_Operator_out3021_out1 <= Logical_Operator_out1997_out1 XOR Logical_Operator_out1999_out1;

  Logical_Operator_out3022_out1 <= Logical_Operator_out1998_out1 XOR Logical_Operator_out2000_out1;

  Logical_Operator_out3023_out1 <= Logical_Operator_out974_out1 XOR Logical_Operator_out976_out1;

  Logical_Operator_out3024_out1 <= in1948 XOR in1952;

  Logical_Operator_out3025_out1 <= Logical_Operator_out2001_out1 XOR Logical_Operator_out2003_out1;

  Logical_Operator_out3026_out1 <= Logical_Operator_out2002_out1 XOR Logical_Operator_out2004_out1;

  Logical_Operator_out3027_out1 <= Logical_Operator_out978_out1 XOR Logical_Operator_out980_out1;

  Logical_Operator_out3028_out1 <= in1956 XOR in1960;

  Logical_Operator_out3029_out1 <= Logical_Operator_out2005_out1 XOR Logical_Operator_out2007_out1;

  Logical_Operator_out3030_out1 <= Logical_Operator_out2006_out1 XOR Logical_Operator_out2008_out1;

  Logical_Operator_out3031_out1 <= Logical_Operator_out982_out1 XOR Logical_Operator_out984_out1;

  Logical_Operator_out3032_out1 <= in1964 XOR in1968;

  Logical_Operator_out3033_out1 <= Logical_Operator_out2009_out1 XOR Logical_Operator_out2011_out1;

  Logical_Operator_out3034_out1 <= Logical_Operator_out2010_out1 XOR Logical_Operator_out2012_out1;

  Logical_Operator_out3035_out1 <= Logical_Operator_out986_out1 XOR Logical_Operator_out988_out1;

  Logical_Operator_out3036_out1 <= in1972 XOR in1976;

  Logical_Operator_out3037_out1 <= Logical_Operator_out2013_out1 XOR Logical_Operator_out2015_out1;

  Logical_Operator_out3038_out1 <= Logical_Operator_out2014_out1 XOR Logical_Operator_out2016_out1;

  Logical_Operator_out3039_out1 <= Logical_Operator_out990_out1 XOR Logical_Operator_out992_out1;

  Logical_Operator_out3040_out1 <= in1980 XOR in1984;

  Logical_Operator_out3041_out1 <= Logical_Operator_out2017_out1 XOR Logical_Operator_out2019_out1;

  Logical_Operator_out3042_out1 <= Logical_Operator_out2018_out1 XOR Logical_Operator_out2020_out1;

  Logical_Operator_out3043_out1 <= Logical_Operator_out994_out1 XOR Logical_Operator_out996_out1;

  Logical_Operator_out3044_out1 <= in1988 XOR in1992;

  Logical_Operator_out3045_out1 <= Logical_Operator_out2021_out1 XOR Logical_Operator_out2023_out1;

  Logical_Operator_out3046_out1 <= Logical_Operator_out2022_out1 XOR Logical_Operator_out2024_out1;

  Logical_Operator_out3047_out1 <= Logical_Operator_out998_out1 XOR Logical_Operator_out1000_out1;

  Logical_Operator_out3048_out1 <= in1996 XOR in2000;

  Logical_Operator_out3049_out1 <= Logical_Operator_out2025_out1 XOR Logical_Operator_out2027_out1;

  Logical_Operator_out3050_out1 <= Logical_Operator_out2026_out1 XOR Logical_Operator_out2028_out1;

  Logical_Operator_out3051_out1 <= Logical_Operator_out1002_out1 XOR Logical_Operator_out1004_out1;

  Logical_Operator_out3052_out1 <= in2004 XOR in2008;

  Logical_Operator_out3053_out1 <= Logical_Operator_out2029_out1 XOR Logical_Operator_out2031_out1;

  Logical_Operator_out3054_out1 <= Logical_Operator_out2030_out1 XOR Logical_Operator_out2032_out1;

  Logical_Operator_out3055_out1 <= Logical_Operator_out1006_out1 XOR Logical_Operator_out1008_out1;

  Logical_Operator_out3056_out1 <= in2012 XOR in2016;

  Logical_Operator_out3057_out1 <= Logical_Operator_out2033_out1 XOR Logical_Operator_out2035_out1;

  Logical_Operator_out3058_out1 <= Logical_Operator_out2034_out1 XOR Logical_Operator_out2036_out1;

  Logical_Operator_out3059_out1 <= Logical_Operator_out1010_out1 XOR Logical_Operator_out1012_out1;

  Logical_Operator_out3060_out1 <= in2020 XOR in2024;

  Logical_Operator_out3061_out1 <= Logical_Operator_out2037_out1 XOR Logical_Operator_out2039_out1;

  Logical_Operator_out3062_out1 <= Logical_Operator_out2038_out1 XOR Logical_Operator_out2040_out1;

  Logical_Operator_out3063_out1 <= Logical_Operator_out1014_out1 XOR Logical_Operator_out1016_out1;

  Logical_Operator_out3064_out1 <= in2028 XOR in2032;

  Logical_Operator_out3065_out1 <= Logical_Operator_out2041_out1 XOR Logical_Operator_out2043_out1;

  Logical_Operator_out3066_out1 <= Logical_Operator_out2042_out1 XOR Logical_Operator_out2044_out1;

  Logical_Operator_out3067_out1 <= Logical_Operator_out1018_out1 XOR Logical_Operator_out1020_out1;

  Logical_Operator_out3068_out1 <= in2036 XOR in2040;

  Logical_Operator_out3069_out1 <= Logical_Operator_out2045_out1 XOR Logical_Operator_out2047_out1;

  Logical_Operator_out3070_out1 <= Logical_Operator_out2046_out1 XOR Logical_Operator_out2048_out1;

  Logical_Operator_out3071_out1 <= Logical_Operator_out1022_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out3072_out1 <= in2044 XOR in2048;

  Logical_Operator_out3073_out1 <= Logical_Operator_out2049_out1 XOR Logical_Operator_out2053_out1;

  Logical_Operator_out3074_out1 <= Logical_Operator_out2050_out1 XOR Logical_Operator_out2054_out1;

  Logical_Operator_out3075_out1 <= Logical_Operator_out2051_out1 XOR Logical_Operator_out2055_out1;

  Logical_Operator_out3076_out1 <= Logical_Operator_out2052_out1 XOR Logical_Operator_out2056_out1;

  Logical_Operator_out3077_out1 <= Logical_Operator_out1027_out1 XOR Logical_Operator_out1031_out1;

  Logical_Operator_out3078_out1 <= Logical_Operator_out1028_out1 XOR Logical_Operator_out1032_out1;

  Logical_Operator_out3079_out1 <= Logical_Operator_out4_out1 XOR Logical_Operator_out8_out1;

  Logical_Operator_out3080_out1 <= in8 XOR in16;

  Logical_Operator_out3081_out1 <= Logical_Operator_out2057_out1 XOR Logical_Operator_out2061_out1;

  Logical_Operator_out3082_out1 <= Logical_Operator_out2058_out1 XOR Logical_Operator_out2062_out1;

  Logical_Operator_out3083_out1 <= Logical_Operator_out2059_out1 XOR Logical_Operator_out2063_out1;

  Logical_Operator_out3084_out1 <= Logical_Operator_out2060_out1 XOR Logical_Operator_out2064_out1;

  Logical_Operator_out3085_out1 <= Logical_Operator_out1035_out1 XOR Logical_Operator_out1039_out1;

  Logical_Operator_out3086_out1 <= Logical_Operator_out1036_out1 XOR Logical_Operator_out1040_out1;

  Logical_Operator_out3087_out1 <= Logical_Operator_out12_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out3088_out1 <= in24 XOR in32;

  Logical_Operator_out3089_out1 <= Logical_Operator_out2065_out1 XOR Logical_Operator_out2069_out1;

  Logical_Operator_out3090_out1 <= Logical_Operator_out2066_out1 XOR Logical_Operator_out2070_out1;

  Logical_Operator_out3091_out1 <= Logical_Operator_out2067_out1 XOR Logical_Operator_out2071_out1;

  Logical_Operator_out3092_out1 <= Logical_Operator_out2068_out1 XOR Logical_Operator_out2072_out1;

  Logical_Operator_out3093_out1 <= Logical_Operator_out1043_out1 XOR Logical_Operator_out1047_out1;

  Logical_Operator_out3094_out1 <= Logical_Operator_out1044_out1 XOR Logical_Operator_out1048_out1;

  Logical_Operator_out3095_out1 <= Logical_Operator_out20_out1 XOR Logical_Operator_out24_out1;

  Logical_Operator_out3096_out1 <= in40 XOR in48;

  Logical_Operator_out3097_out1 <= Logical_Operator_out2073_out1 XOR Logical_Operator_out2077_out1;

  Logical_Operator_out3098_out1 <= Logical_Operator_out2074_out1 XOR Logical_Operator_out2078_out1;

  Logical_Operator_out3099_out1 <= Logical_Operator_out2075_out1 XOR Logical_Operator_out2079_out1;

  Logical_Operator_out3100_out1 <= Logical_Operator_out2076_out1 XOR Logical_Operator_out2080_out1;

  Logical_Operator_out3101_out1 <= Logical_Operator_out1051_out1 XOR Logical_Operator_out1055_out1;

  Logical_Operator_out3102_out1 <= Logical_Operator_out1052_out1 XOR Logical_Operator_out1056_out1;

  Logical_Operator_out3103_out1 <= Logical_Operator_out28_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out3104_out1 <= in56 XOR in64;

  Logical_Operator_out3105_out1 <= Logical_Operator_out2081_out1 XOR Logical_Operator_out2085_out1;

  Logical_Operator_out3106_out1 <= Logical_Operator_out2082_out1 XOR Logical_Operator_out2086_out1;

  Logical_Operator_out3107_out1 <= Logical_Operator_out2083_out1 XOR Logical_Operator_out2087_out1;

  Logical_Operator_out3108_out1 <= Logical_Operator_out2084_out1 XOR Logical_Operator_out2088_out1;

  Logical_Operator_out3109_out1 <= Logical_Operator_out1059_out1 XOR Logical_Operator_out1063_out1;

  Logical_Operator_out3110_out1 <= Logical_Operator_out1060_out1 XOR Logical_Operator_out1064_out1;

  Logical_Operator_out3111_out1 <= Logical_Operator_out36_out1 XOR Logical_Operator_out40_out1;

  Logical_Operator_out3112_out1 <= in72 XOR in80;

  Logical_Operator_out3113_out1 <= Logical_Operator_out2089_out1 XOR Logical_Operator_out2093_out1;

  Logical_Operator_out3114_out1 <= Logical_Operator_out2090_out1 XOR Logical_Operator_out2094_out1;

  Logical_Operator_out3115_out1 <= Logical_Operator_out2091_out1 XOR Logical_Operator_out2095_out1;

  Logical_Operator_out3116_out1 <= Logical_Operator_out2092_out1 XOR Logical_Operator_out2096_out1;

  Logical_Operator_out3117_out1 <= Logical_Operator_out1067_out1 XOR Logical_Operator_out1071_out1;

  Logical_Operator_out3118_out1 <= Logical_Operator_out1068_out1 XOR Logical_Operator_out1072_out1;

  Logical_Operator_out3119_out1 <= Logical_Operator_out44_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out3120_out1 <= in88 XOR in96;

  Logical_Operator_out3121_out1 <= Logical_Operator_out2097_out1 XOR Logical_Operator_out2101_out1;

  Logical_Operator_out3122_out1 <= Logical_Operator_out2098_out1 XOR Logical_Operator_out2102_out1;

  Logical_Operator_out3123_out1 <= Logical_Operator_out2099_out1 XOR Logical_Operator_out2103_out1;

  Logical_Operator_out3124_out1 <= Logical_Operator_out2100_out1 XOR Logical_Operator_out2104_out1;

  Logical_Operator_out3125_out1 <= Logical_Operator_out1075_out1 XOR Logical_Operator_out1079_out1;

  Logical_Operator_out3126_out1 <= Logical_Operator_out1076_out1 XOR Logical_Operator_out1080_out1;

  Logical_Operator_out3127_out1 <= Logical_Operator_out52_out1 XOR Logical_Operator_out56_out1;

  Logical_Operator_out3128_out1 <= in104 XOR in112;

  Logical_Operator_out3129_out1 <= Logical_Operator_out2105_out1 XOR Logical_Operator_out2109_out1;

  Logical_Operator_out3130_out1 <= Logical_Operator_out2106_out1 XOR Logical_Operator_out2110_out1;

  Logical_Operator_out3131_out1 <= Logical_Operator_out2107_out1 XOR Logical_Operator_out2111_out1;

  Logical_Operator_out3132_out1 <= Logical_Operator_out2108_out1 XOR Logical_Operator_out2112_out1;

  Logical_Operator_out3133_out1 <= Logical_Operator_out1083_out1 XOR Logical_Operator_out1087_out1;

  Logical_Operator_out3134_out1 <= Logical_Operator_out1084_out1 XOR Logical_Operator_out1088_out1;

  Logical_Operator_out3135_out1 <= Logical_Operator_out60_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out3136_out1 <= in120 XOR in128;

  Logical_Operator_out3137_out1 <= Logical_Operator_out2113_out1 XOR Logical_Operator_out2117_out1;

  Logical_Operator_out3138_out1 <= Logical_Operator_out2114_out1 XOR Logical_Operator_out2118_out1;

  Logical_Operator_out3139_out1 <= Logical_Operator_out2115_out1 XOR Logical_Operator_out2119_out1;

  Logical_Operator_out3140_out1 <= Logical_Operator_out2116_out1 XOR Logical_Operator_out2120_out1;

  Logical_Operator_out3141_out1 <= Logical_Operator_out1091_out1 XOR Logical_Operator_out1095_out1;

  Logical_Operator_out3142_out1 <= Logical_Operator_out1092_out1 XOR Logical_Operator_out1096_out1;

  Logical_Operator_out3143_out1 <= Logical_Operator_out68_out1 XOR Logical_Operator_out72_out1;

  Logical_Operator_out3144_out1 <= in136 XOR in144;

  Logical_Operator_out3145_out1 <= Logical_Operator_out2121_out1 XOR Logical_Operator_out2125_out1;

  Logical_Operator_out3146_out1 <= Logical_Operator_out2122_out1 XOR Logical_Operator_out2126_out1;

  Logical_Operator_out3147_out1 <= Logical_Operator_out2123_out1 XOR Logical_Operator_out2127_out1;

  Logical_Operator_out3148_out1 <= Logical_Operator_out2124_out1 XOR Logical_Operator_out2128_out1;

  Logical_Operator_out3149_out1 <= Logical_Operator_out1099_out1 XOR Logical_Operator_out1103_out1;

  Logical_Operator_out3150_out1 <= Logical_Operator_out1100_out1 XOR Logical_Operator_out1104_out1;

  Logical_Operator_out3151_out1 <= Logical_Operator_out76_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out3152_out1 <= in152 XOR in160;

  Logical_Operator_out3153_out1 <= Logical_Operator_out2129_out1 XOR Logical_Operator_out2133_out1;

  Logical_Operator_out3154_out1 <= Logical_Operator_out2130_out1 XOR Logical_Operator_out2134_out1;

  Logical_Operator_out3155_out1 <= Logical_Operator_out2131_out1 XOR Logical_Operator_out2135_out1;

  Logical_Operator_out3156_out1 <= Logical_Operator_out2132_out1 XOR Logical_Operator_out2136_out1;

  Logical_Operator_out3157_out1 <= Logical_Operator_out1107_out1 XOR Logical_Operator_out1111_out1;

  Logical_Operator_out3158_out1 <= Logical_Operator_out1108_out1 XOR Logical_Operator_out1112_out1;

  Logical_Operator_out3159_out1 <= Logical_Operator_out84_out1 XOR Logical_Operator_out88_out1;

  Logical_Operator_out3160_out1 <= in168 XOR in176;

  Logical_Operator_out3161_out1 <= Logical_Operator_out2137_out1 XOR Logical_Operator_out2141_out1;

  Logical_Operator_out3162_out1 <= Logical_Operator_out2138_out1 XOR Logical_Operator_out2142_out1;

  Logical_Operator_out3163_out1 <= Logical_Operator_out2139_out1 XOR Logical_Operator_out2143_out1;

  Logical_Operator_out3164_out1 <= Logical_Operator_out2140_out1 XOR Logical_Operator_out2144_out1;

  Logical_Operator_out3165_out1 <= Logical_Operator_out1115_out1 XOR Logical_Operator_out1119_out1;

  Logical_Operator_out3166_out1 <= Logical_Operator_out1116_out1 XOR Logical_Operator_out1120_out1;

  Logical_Operator_out3167_out1 <= Logical_Operator_out92_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out3168_out1 <= in184 XOR in192;

  Logical_Operator_out3169_out1 <= Logical_Operator_out2145_out1 XOR Logical_Operator_out2149_out1;

  Logical_Operator_out3170_out1 <= Logical_Operator_out2146_out1 XOR Logical_Operator_out2150_out1;

  Logical_Operator_out3171_out1 <= Logical_Operator_out2147_out1 XOR Logical_Operator_out2151_out1;

  Logical_Operator_out3172_out1 <= Logical_Operator_out2148_out1 XOR Logical_Operator_out2152_out1;

  Logical_Operator_out3173_out1 <= Logical_Operator_out1123_out1 XOR Logical_Operator_out1127_out1;

  Logical_Operator_out3174_out1 <= Logical_Operator_out1124_out1 XOR Logical_Operator_out1128_out1;

  Logical_Operator_out3175_out1 <= Logical_Operator_out100_out1 XOR Logical_Operator_out104_out1;

  Logical_Operator_out3176_out1 <= in200 XOR in208;

  Logical_Operator_out3177_out1 <= Logical_Operator_out2153_out1 XOR Logical_Operator_out2157_out1;

  Logical_Operator_out3178_out1 <= Logical_Operator_out2154_out1 XOR Logical_Operator_out2158_out1;

  Logical_Operator_out3179_out1 <= Logical_Operator_out2155_out1 XOR Logical_Operator_out2159_out1;

  Logical_Operator_out3180_out1 <= Logical_Operator_out2156_out1 XOR Logical_Operator_out2160_out1;

  Logical_Operator_out3181_out1 <= Logical_Operator_out1131_out1 XOR Logical_Operator_out1135_out1;

  Logical_Operator_out3182_out1 <= Logical_Operator_out1132_out1 XOR Logical_Operator_out1136_out1;

  Logical_Operator_out3183_out1 <= Logical_Operator_out108_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out3184_out1 <= in216 XOR in224;

  Logical_Operator_out3185_out1 <= Logical_Operator_out2161_out1 XOR Logical_Operator_out2165_out1;

  Logical_Operator_out3186_out1 <= Logical_Operator_out2162_out1 XOR Logical_Operator_out2166_out1;

  Logical_Operator_out3187_out1 <= Logical_Operator_out2163_out1 XOR Logical_Operator_out2167_out1;

  Logical_Operator_out3188_out1 <= Logical_Operator_out2164_out1 XOR Logical_Operator_out2168_out1;

  Logical_Operator_out3189_out1 <= Logical_Operator_out1139_out1 XOR Logical_Operator_out1143_out1;

  Logical_Operator_out3190_out1 <= Logical_Operator_out1140_out1 XOR Logical_Operator_out1144_out1;

  Logical_Operator_out3191_out1 <= Logical_Operator_out116_out1 XOR Logical_Operator_out120_out1;

  Logical_Operator_out3192_out1 <= in232 XOR in240;

  Logical_Operator_out3193_out1 <= Logical_Operator_out2169_out1 XOR Logical_Operator_out2173_out1;

  Logical_Operator_out3194_out1 <= Logical_Operator_out2170_out1 XOR Logical_Operator_out2174_out1;

  Logical_Operator_out3195_out1 <= Logical_Operator_out2171_out1 XOR Logical_Operator_out2175_out1;

  Logical_Operator_out3196_out1 <= Logical_Operator_out2172_out1 XOR Logical_Operator_out2176_out1;

  Logical_Operator_out3197_out1 <= Logical_Operator_out1147_out1 XOR Logical_Operator_out1151_out1;

  Logical_Operator_out3198_out1 <= Logical_Operator_out1148_out1 XOR Logical_Operator_out1152_out1;

  Logical_Operator_out3199_out1 <= Logical_Operator_out124_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out3200_out1 <= in248 XOR in256;

  Logical_Operator_out3201_out1 <= Logical_Operator_out2177_out1 XOR Logical_Operator_out2181_out1;

  Logical_Operator_out3202_out1 <= Logical_Operator_out2178_out1 XOR Logical_Operator_out2182_out1;

  Logical_Operator_out3203_out1 <= Logical_Operator_out2179_out1 XOR Logical_Operator_out2183_out1;

  Logical_Operator_out3204_out1 <= Logical_Operator_out2180_out1 XOR Logical_Operator_out2184_out1;

  Logical_Operator_out3205_out1 <= Logical_Operator_out1155_out1 XOR Logical_Operator_out1159_out1;

  Logical_Operator_out3206_out1 <= Logical_Operator_out1156_out1 XOR Logical_Operator_out1160_out1;

  Logical_Operator_out3207_out1 <= Logical_Operator_out132_out1 XOR Logical_Operator_out136_out1;

  Logical_Operator_out3208_out1 <= in264 XOR in272;

  Logical_Operator_out3209_out1 <= Logical_Operator_out2185_out1 XOR Logical_Operator_out2189_out1;

  Logical_Operator_out3210_out1 <= Logical_Operator_out2186_out1 XOR Logical_Operator_out2190_out1;

  Logical_Operator_out3211_out1 <= Logical_Operator_out2187_out1 XOR Logical_Operator_out2191_out1;

  Logical_Operator_out3212_out1 <= Logical_Operator_out2188_out1 XOR Logical_Operator_out2192_out1;

  Logical_Operator_out3213_out1 <= Logical_Operator_out1163_out1 XOR Logical_Operator_out1167_out1;

  Logical_Operator_out3214_out1 <= Logical_Operator_out1164_out1 XOR Logical_Operator_out1168_out1;

  Logical_Operator_out3215_out1 <= Logical_Operator_out140_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out3216_out1 <= in280 XOR in288;

  Logical_Operator_out3217_out1 <= Logical_Operator_out2193_out1 XOR Logical_Operator_out2197_out1;

  Logical_Operator_out3218_out1 <= Logical_Operator_out2194_out1 XOR Logical_Operator_out2198_out1;

  Logical_Operator_out3219_out1 <= Logical_Operator_out2195_out1 XOR Logical_Operator_out2199_out1;

  Logical_Operator_out3220_out1 <= Logical_Operator_out2196_out1 XOR Logical_Operator_out2200_out1;

  Logical_Operator_out3221_out1 <= Logical_Operator_out1171_out1 XOR Logical_Operator_out1175_out1;

  Logical_Operator_out3222_out1 <= Logical_Operator_out1172_out1 XOR Logical_Operator_out1176_out1;

  Logical_Operator_out3223_out1 <= Logical_Operator_out148_out1 XOR Logical_Operator_out152_out1;

  Logical_Operator_out3224_out1 <= in296 XOR in304;

  Logical_Operator_out3225_out1 <= Logical_Operator_out2201_out1 XOR Logical_Operator_out2205_out1;

  Logical_Operator_out3226_out1 <= Logical_Operator_out2202_out1 XOR Logical_Operator_out2206_out1;

  Logical_Operator_out3227_out1 <= Logical_Operator_out2203_out1 XOR Logical_Operator_out2207_out1;

  Logical_Operator_out3228_out1 <= Logical_Operator_out2204_out1 XOR Logical_Operator_out2208_out1;

  Logical_Operator_out3229_out1 <= Logical_Operator_out1179_out1 XOR Logical_Operator_out1183_out1;

  Logical_Operator_out3230_out1 <= Logical_Operator_out1180_out1 XOR Logical_Operator_out1184_out1;

  Logical_Operator_out3231_out1 <= Logical_Operator_out156_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out3232_out1 <= in312 XOR in320;

  Logical_Operator_out3233_out1 <= Logical_Operator_out2209_out1 XOR Logical_Operator_out2213_out1;

  Logical_Operator_out3234_out1 <= Logical_Operator_out2210_out1 XOR Logical_Operator_out2214_out1;

  Logical_Operator_out3235_out1 <= Logical_Operator_out2211_out1 XOR Logical_Operator_out2215_out1;

  Logical_Operator_out3236_out1 <= Logical_Operator_out2212_out1 XOR Logical_Operator_out2216_out1;

  Logical_Operator_out3237_out1 <= Logical_Operator_out1187_out1 XOR Logical_Operator_out1191_out1;

  Logical_Operator_out3238_out1 <= Logical_Operator_out1188_out1 XOR Logical_Operator_out1192_out1;

  Logical_Operator_out3239_out1 <= Logical_Operator_out164_out1 XOR Logical_Operator_out168_out1;

  Logical_Operator_out3240_out1 <= in328 XOR in336;

  Logical_Operator_out3241_out1 <= Logical_Operator_out2217_out1 XOR Logical_Operator_out2221_out1;

  Logical_Operator_out3242_out1 <= Logical_Operator_out2218_out1 XOR Logical_Operator_out2222_out1;

  Logical_Operator_out3243_out1 <= Logical_Operator_out2219_out1 XOR Logical_Operator_out2223_out1;

  Logical_Operator_out3244_out1 <= Logical_Operator_out2220_out1 XOR Logical_Operator_out2224_out1;

  Logical_Operator_out3245_out1 <= Logical_Operator_out1195_out1 XOR Logical_Operator_out1199_out1;

  Logical_Operator_out3246_out1 <= Logical_Operator_out1196_out1 XOR Logical_Operator_out1200_out1;

  Logical_Operator_out3247_out1 <= Logical_Operator_out172_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out3248_out1 <= in344 XOR in352;

  Logical_Operator_out3249_out1 <= Logical_Operator_out2225_out1 XOR Logical_Operator_out2229_out1;

  Logical_Operator_out3250_out1 <= Logical_Operator_out2226_out1 XOR Logical_Operator_out2230_out1;

  Logical_Operator_out3251_out1 <= Logical_Operator_out2227_out1 XOR Logical_Operator_out2231_out1;

  Logical_Operator_out3252_out1 <= Logical_Operator_out2228_out1 XOR Logical_Operator_out2232_out1;

  Logical_Operator_out3253_out1 <= Logical_Operator_out1203_out1 XOR Logical_Operator_out1207_out1;

  Logical_Operator_out3254_out1 <= Logical_Operator_out1204_out1 XOR Logical_Operator_out1208_out1;

  Logical_Operator_out3255_out1 <= Logical_Operator_out180_out1 XOR Logical_Operator_out184_out1;

  Logical_Operator_out3256_out1 <= in360 XOR in368;

  Logical_Operator_out3257_out1 <= Logical_Operator_out2233_out1 XOR Logical_Operator_out2237_out1;

  Logical_Operator_out3258_out1 <= Logical_Operator_out2234_out1 XOR Logical_Operator_out2238_out1;

  Logical_Operator_out3259_out1 <= Logical_Operator_out2235_out1 XOR Logical_Operator_out2239_out1;

  Logical_Operator_out3260_out1 <= Logical_Operator_out2236_out1 XOR Logical_Operator_out2240_out1;

  Logical_Operator_out3261_out1 <= Logical_Operator_out1211_out1 XOR Logical_Operator_out1215_out1;

  Logical_Operator_out3262_out1 <= Logical_Operator_out1212_out1 XOR Logical_Operator_out1216_out1;

  Logical_Operator_out3263_out1 <= Logical_Operator_out188_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out3264_out1 <= in376 XOR in384;

  Logical_Operator_out3265_out1 <= Logical_Operator_out2241_out1 XOR Logical_Operator_out2245_out1;

  Logical_Operator_out3266_out1 <= Logical_Operator_out2242_out1 XOR Logical_Operator_out2246_out1;

  Logical_Operator_out3267_out1 <= Logical_Operator_out2243_out1 XOR Logical_Operator_out2247_out1;

  Logical_Operator_out3268_out1 <= Logical_Operator_out2244_out1 XOR Logical_Operator_out2248_out1;

  Logical_Operator_out3269_out1 <= Logical_Operator_out1219_out1 XOR Logical_Operator_out1223_out1;

  Logical_Operator_out3270_out1 <= Logical_Operator_out1220_out1 XOR Logical_Operator_out1224_out1;

  Logical_Operator_out3271_out1 <= Logical_Operator_out196_out1 XOR Logical_Operator_out200_out1;

  Logical_Operator_out3272_out1 <= in392 XOR in400;

  Logical_Operator_out3273_out1 <= Logical_Operator_out2249_out1 XOR Logical_Operator_out2253_out1;

  Logical_Operator_out3274_out1 <= Logical_Operator_out2250_out1 XOR Logical_Operator_out2254_out1;

  Logical_Operator_out3275_out1 <= Logical_Operator_out2251_out1 XOR Logical_Operator_out2255_out1;

  Logical_Operator_out3276_out1 <= Logical_Operator_out2252_out1 XOR Logical_Operator_out2256_out1;

  Logical_Operator_out3277_out1 <= Logical_Operator_out1227_out1 XOR Logical_Operator_out1231_out1;

  Logical_Operator_out3278_out1 <= Logical_Operator_out1228_out1 XOR Logical_Operator_out1232_out1;

  Logical_Operator_out3279_out1 <= Logical_Operator_out204_out1 XOR Logical_Operator_out208_out1;

  Logical_Operator_out3280_out1 <= in408 XOR in416;

  Logical_Operator_out3281_out1 <= Logical_Operator_out2257_out1 XOR Logical_Operator_out2261_out1;

  Logical_Operator_out3282_out1 <= Logical_Operator_out2258_out1 XOR Logical_Operator_out2262_out1;

  Logical_Operator_out3283_out1 <= Logical_Operator_out2259_out1 XOR Logical_Operator_out2263_out1;

  Logical_Operator_out3284_out1 <= Logical_Operator_out2260_out1 XOR Logical_Operator_out2264_out1;

  Logical_Operator_out3285_out1 <= Logical_Operator_out1235_out1 XOR Logical_Operator_out1239_out1;

  Logical_Operator_out3286_out1 <= Logical_Operator_out1236_out1 XOR Logical_Operator_out1240_out1;

  Logical_Operator_out3287_out1 <= Logical_Operator_out212_out1 XOR Logical_Operator_out216_out1;

  Logical_Operator_out3288_out1 <= in424 XOR in432;

  Logical_Operator_out3289_out1 <= Logical_Operator_out2265_out1 XOR Logical_Operator_out2269_out1;

  Logical_Operator_out3290_out1 <= Logical_Operator_out2266_out1 XOR Logical_Operator_out2270_out1;

  Logical_Operator_out3291_out1 <= Logical_Operator_out2267_out1 XOR Logical_Operator_out2271_out1;

  Logical_Operator_out3292_out1 <= Logical_Operator_out2268_out1 XOR Logical_Operator_out2272_out1;

  Logical_Operator_out3293_out1 <= Logical_Operator_out1243_out1 XOR Logical_Operator_out1247_out1;

  Logical_Operator_out3294_out1 <= Logical_Operator_out1244_out1 XOR Logical_Operator_out1248_out1;

  Logical_Operator_out3295_out1 <= Logical_Operator_out220_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out3296_out1 <= in440 XOR in448;

  Logical_Operator_out3297_out1 <= Logical_Operator_out2273_out1 XOR Logical_Operator_out2277_out1;

  Logical_Operator_out3298_out1 <= Logical_Operator_out2274_out1 XOR Logical_Operator_out2278_out1;

  Logical_Operator_out3299_out1 <= Logical_Operator_out2275_out1 XOR Logical_Operator_out2279_out1;

  Logical_Operator_out3300_out1 <= Logical_Operator_out2276_out1 XOR Logical_Operator_out2280_out1;

  Logical_Operator_out3301_out1 <= Logical_Operator_out1251_out1 XOR Logical_Operator_out1255_out1;

  Logical_Operator_out3302_out1 <= Logical_Operator_out1252_out1 XOR Logical_Operator_out1256_out1;

  Logical_Operator_out3303_out1 <= Logical_Operator_out228_out1 XOR Logical_Operator_out232_out1;

  Logical_Operator_out3304_out1 <= in456 XOR in464;

  Logical_Operator_out3305_out1 <= Logical_Operator_out2281_out1 XOR Logical_Operator_out2285_out1;

  Logical_Operator_out3306_out1 <= Logical_Operator_out2282_out1 XOR Logical_Operator_out2286_out1;

  Logical_Operator_out3307_out1 <= Logical_Operator_out2283_out1 XOR Logical_Operator_out2287_out1;

  Logical_Operator_out3308_out1 <= Logical_Operator_out2284_out1 XOR Logical_Operator_out2288_out1;

  Logical_Operator_out3309_out1 <= Logical_Operator_out1259_out1 XOR Logical_Operator_out1263_out1;

  Logical_Operator_out3310_out1 <= Logical_Operator_out1260_out1 XOR Logical_Operator_out1264_out1;

  Logical_Operator_out3311_out1 <= Logical_Operator_out236_out1 XOR Logical_Operator_out240_out1;

  Logical_Operator_out3312_out1 <= in472 XOR in480;

  Logical_Operator_out3313_out1 <= Logical_Operator_out2289_out1 XOR Logical_Operator_out2293_out1;

  Logical_Operator_out3314_out1 <= Logical_Operator_out2290_out1 XOR Logical_Operator_out2294_out1;

  Logical_Operator_out3315_out1 <= Logical_Operator_out2291_out1 XOR Logical_Operator_out2295_out1;

  Logical_Operator_out3316_out1 <= Logical_Operator_out2292_out1 XOR Logical_Operator_out2296_out1;

  Logical_Operator_out3317_out1 <= Logical_Operator_out1267_out1 XOR Logical_Operator_out1271_out1;

  Logical_Operator_out3318_out1 <= Logical_Operator_out1268_out1 XOR Logical_Operator_out1272_out1;

  Logical_Operator_out3319_out1 <= Logical_Operator_out244_out1 XOR Logical_Operator_out248_out1;

  Logical_Operator_out3320_out1 <= in488 XOR in496;

  Logical_Operator_out3321_out1 <= Logical_Operator_out2297_out1 XOR Logical_Operator_out2301_out1;

  Logical_Operator_out3322_out1 <= Logical_Operator_out2298_out1 XOR Logical_Operator_out2302_out1;

  Logical_Operator_out3323_out1 <= Logical_Operator_out2299_out1 XOR Logical_Operator_out2303_out1;

  Logical_Operator_out3324_out1 <= Logical_Operator_out2300_out1 XOR Logical_Operator_out2304_out1;

  Logical_Operator_out3325_out1 <= Logical_Operator_out1275_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out3326_out1 <= Logical_Operator_out1276_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out3327_out1 <= Logical_Operator_out252_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out3328_out1 <= in504 XOR in512;

  Logical_Operator_out3329_out1 <= Logical_Operator_out2305_out1 XOR Logical_Operator_out2309_out1;

  Logical_Operator_out3330_out1 <= Logical_Operator_out2306_out1 XOR Logical_Operator_out2310_out1;

  Logical_Operator_out3331_out1 <= Logical_Operator_out2307_out1 XOR Logical_Operator_out2311_out1;

  Logical_Operator_out3332_out1 <= Logical_Operator_out2308_out1 XOR Logical_Operator_out2312_out1;

  Logical_Operator_out3333_out1 <= Logical_Operator_out1283_out1 XOR Logical_Operator_out1287_out1;

  Logical_Operator_out3334_out1 <= Logical_Operator_out1284_out1 XOR Logical_Operator_out1288_out1;

  Logical_Operator_out3335_out1 <= Logical_Operator_out260_out1 XOR Logical_Operator_out264_out1;

  Logical_Operator_out3336_out1 <= in520 XOR in528;

  Logical_Operator_out3337_out1 <= Logical_Operator_out2313_out1 XOR Logical_Operator_out2317_out1;

  Logical_Operator_out3338_out1 <= Logical_Operator_out2314_out1 XOR Logical_Operator_out2318_out1;

  Logical_Operator_out3339_out1 <= Logical_Operator_out2315_out1 XOR Logical_Operator_out2319_out1;

  Logical_Operator_out3340_out1 <= Logical_Operator_out2316_out1 XOR Logical_Operator_out2320_out1;

  Logical_Operator_out3341_out1 <= Logical_Operator_out1291_out1 XOR Logical_Operator_out1295_out1;

  Logical_Operator_out3342_out1 <= Logical_Operator_out1292_out1 XOR Logical_Operator_out1296_out1;

  Logical_Operator_out3343_out1 <= Logical_Operator_out268_out1 XOR Logical_Operator_out272_out1;

  Logical_Operator_out3344_out1 <= in536 XOR in544;

  Logical_Operator_out3345_out1 <= Logical_Operator_out2321_out1 XOR Logical_Operator_out2325_out1;

  Logical_Operator_out3346_out1 <= Logical_Operator_out2322_out1 XOR Logical_Operator_out2326_out1;

  Logical_Operator_out3347_out1 <= Logical_Operator_out2323_out1 XOR Logical_Operator_out2327_out1;

  Logical_Operator_out3348_out1 <= Logical_Operator_out2324_out1 XOR Logical_Operator_out2328_out1;

  Logical_Operator_out3349_out1 <= Logical_Operator_out1299_out1 XOR Logical_Operator_out1303_out1;

  Logical_Operator_out3350_out1 <= Logical_Operator_out1300_out1 XOR Logical_Operator_out1304_out1;

  Logical_Operator_out3351_out1 <= Logical_Operator_out276_out1 XOR Logical_Operator_out280_out1;

  Logical_Operator_out3352_out1 <= in552 XOR in560;

  Logical_Operator_out3353_out1 <= Logical_Operator_out2329_out1 XOR Logical_Operator_out2333_out1;

  Logical_Operator_out3354_out1 <= Logical_Operator_out2330_out1 XOR Logical_Operator_out2334_out1;

  Logical_Operator_out3355_out1 <= Logical_Operator_out2331_out1 XOR Logical_Operator_out2335_out1;

  Logical_Operator_out3356_out1 <= Logical_Operator_out2332_out1 XOR Logical_Operator_out2336_out1;

  Logical_Operator_out3357_out1 <= Logical_Operator_out1307_out1 XOR Logical_Operator_out1311_out1;

  Logical_Operator_out3358_out1 <= Logical_Operator_out1308_out1 XOR Logical_Operator_out1312_out1;

  Logical_Operator_out3359_out1 <= Logical_Operator_out284_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out3360_out1 <= in568 XOR in576;

  Logical_Operator_out3361_out1 <= Logical_Operator_out2337_out1 XOR Logical_Operator_out2341_out1;

  Logical_Operator_out3362_out1 <= Logical_Operator_out2338_out1 XOR Logical_Operator_out2342_out1;

  Logical_Operator_out3363_out1 <= Logical_Operator_out2339_out1 XOR Logical_Operator_out2343_out1;

  Logical_Operator_out3364_out1 <= Logical_Operator_out2340_out1 XOR Logical_Operator_out2344_out1;

  Logical_Operator_out3365_out1 <= Logical_Operator_out1315_out1 XOR Logical_Operator_out1319_out1;

  Logical_Operator_out3366_out1 <= Logical_Operator_out1316_out1 XOR Logical_Operator_out1320_out1;

  Logical_Operator_out3367_out1 <= Logical_Operator_out292_out1 XOR Logical_Operator_out296_out1;

  Logical_Operator_out3368_out1 <= in584 XOR in592;

  Logical_Operator_out3369_out1 <= Logical_Operator_out2345_out1 XOR Logical_Operator_out2349_out1;

  Logical_Operator_out3370_out1 <= Logical_Operator_out2346_out1 XOR Logical_Operator_out2350_out1;

  Logical_Operator_out3371_out1 <= Logical_Operator_out2347_out1 XOR Logical_Operator_out2351_out1;

  Logical_Operator_out3372_out1 <= Logical_Operator_out2348_out1 XOR Logical_Operator_out2352_out1;

  Logical_Operator_out3373_out1 <= Logical_Operator_out1323_out1 XOR Logical_Operator_out1327_out1;

  Logical_Operator_out3374_out1 <= Logical_Operator_out1324_out1 XOR Logical_Operator_out1328_out1;

  Logical_Operator_out3375_out1 <= Logical_Operator_out300_out1 XOR Logical_Operator_out304_out1;

  Logical_Operator_out3376_out1 <= in600 XOR in608;

  Logical_Operator_out3377_out1 <= Logical_Operator_out2353_out1 XOR Logical_Operator_out2357_out1;

  Logical_Operator_out3378_out1 <= Logical_Operator_out2354_out1 XOR Logical_Operator_out2358_out1;

  Logical_Operator_out3379_out1 <= Logical_Operator_out2355_out1 XOR Logical_Operator_out2359_out1;

  Logical_Operator_out3380_out1 <= Logical_Operator_out2356_out1 XOR Logical_Operator_out2360_out1;

  Logical_Operator_out3381_out1 <= Logical_Operator_out1331_out1 XOR Logical_Operator_out1335_out1;

  Logical_Operator_out3382_out1 <= Logical_Operator_out1332_out1 XOR Logical_Operator_out1336_out1;

  Logical_Operator_out3383_out1 <= Logical_Operator_out308_out1 XOR Logical_Operator_out312_out1;

  Logical_Operator_out3384_out1 <= in616 XOR in624;

  Logical_Operator_out3385_out1 <= Logical_Operator_out2361_out1 XOR Logical_Operator_out2365_out1;

  Logical_Operator_out3386_out1 <= Logical_Operator_out2362_out1 XOR Logical_Operator_out2366_out1;

  Logical_Operator_out3387_out1 <= Logical_Operator_out2363_out1 XOR Logical_Operator_out2367_out1;

  Logical_Operator_out3388_out1 <= Logical_Operator_out2364_out1 XOR Logical_Operator_out2368_out1;

  Logical_Operator_out3389_out1 <= Logical_Operator_out1339_out1 XOR Logical_Operator_out1343_out1;

  Logical_Operator_out3390_out1 <= Logical_Operator_out1340_out1 XOR Logical_Operator_out1344_out1;

  Logical_Operator_out3391_out1 <= Logical_Operator_out316_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out3392_out1 <= in632 XOR in640;

  Logical_Operator_out3393_out1 <= Logical_Operator_out2369_out1 XOR Logical_Operator_out2373_out1;

  Logical_Operator_out3394_out1 <= Logical_Operator_out2370_out1 XOR Logical_Operator_out2374_out1;

  Logical_Operator_out3395_out1 <= Logical_Operator_out2371_out1 XOR Logical_Operator_out2375_out1;

  Logical_Operator_out3396_out1 <= Logical_Operator_out2372_out1 XOR Logical_Operator_out2376_out1;

  Logical_Operator_out3397_out1 <= Logical_Operator_out1347_out1 XOR Logical_Operator_out1351_out1;

  Logical_Operator_out3398_out1 <= Logical_Operator_out1348_out1 XOR Logical_Operator_out1352_out1;

  Logical_Operator_out3399_out1 <= Logical_Operator_out324_out1 XOR Logical_Operator_out328_out1;

  Logical_Operator_out3400_out1 <= in648 XOR in656;

  Logical_Operator_out3401_out1 <= Logical_Operator_out2377_out1 XOR Logical_Operator_out2381_out1;

  Logical_Operator_out3402_out1 <= Logical_Operator_out2378_out1 XOR Logical_Operator_out2382_out1;

  Logical_Operator_out3403_out1 <= Logical_Operator_out2379_out1 XOR Logical_Operator_out2383_out1;

  Logical_Operator_out3404_out1 <= Logical_Operator_out2380_out1 XOR Logical_Operator_out2384_out1;

  Logical_Operator_out3405_out1 <= Logical_Operator_out1355_out1 XOR Logical_Operator_out1359_out1;

  Logical_Operator_out3406_out1 <= Logical_Operator_out1356_out1 XOR Logical_Operator_out1360_out1;

  Logical_Operator_out3407_out1 <= Logical_Operator_out332_out1 XOR Logical_Operator_out336_out1;

  Logical_Operator_out3408_out1 <= in664 XOR in672;

  Logical_Operator_out3409_out1 <= Logical_Operator_out2385_out1 XOR Logical_Operator_out2389_out1;

  Logical_Operator_out3410_out1 <= Logical_Operator_out2386_out1 XOR Logical_Operator_out2390_out1;

  Logical_Operator_out3411_out1 <= Logical_Operator_out2387_out1 XOR Logical_Operator_out2391_out1;

  Logical_Operator_out3412_out1 <= Logical_Operator_out2388_out1 XOR Logical_Operator_out2392_out1;

  Logical_Operator_out3413_out1 <= Logical_Operator_out1363_out1 XOR Logical_Operator_out1367_out1;

  Logical_Operator_out3414_out1 <= Logical_Operator_out1364_out1 XOR Logical_Operator_out1368_out1;

  Logical_Operator_out3415_out1 <= Logical_Operator_out340_out1 XOR Logical_Operator_out344_out1;

  Logical_Operator_out3416_out1 <= in680 XOR in688;

  Logical_Operator_out3417_out1 <= Logical_Operator_out2393_out1 XOR Logical_Operator_out2397_out1;

  Logical_Operator_out3418_out1 <= Logical_Operator_out2394_out1 XOR Logical_Operator_out2398_out1;

  Logical_Operator_out3419_out1 <= Logical_Operator_out2395_out1 XOR Logical_Operator_out2399_out1;

  Logical_Operator_out3420_out1 <= Logical_Operator_out2396_out1 XOR Logical_Operator_out2400_out1;

  Logical_Operator_out3421_out1 <= Logical_Operator_out1371_out1 XOR Logical_Operator_out1375_out1;

  Logical_Operator_out3422_out1 <= Logical_Operator_out1372_out1 XOR Logical_Operator_out1376_out1;

  Logical_Operator_out3423_out1 <= Logical_Operator_out348_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out3424_out1 <= in696 XOR in704;

  Logical_Operator_out3425_out1 <= Logical_Operator_out2401_out1 XOR Logical_Operator_out2405_out1;

  Logical_Operator_out3426_out1 <= Logical_Operator_out2402_out1 XOR Logical_Operator_out2406_out1;

  Logical_Operator_out3427_out1 <= Logical_Operator_out2403_out1 XOR Logical_Operator_out2407_out1;

  Logical_Operator_out3428_out1 <= Logical_Operator_out2404_out1 XOR Logical_Operator_out2408_out1;

  Logical_Operator_out3429_out1 <= Logical_Operator_out1379_out1 XOR Logical_Operator_out1383_out1;

  Logical_Operator_out3430_out1 <= Logical_Operator_out1380_out1 XOR Logical_Operator_out1384_out1;

  Logical_Operator_out3431_out1 <= Logical_Operator_out356_out1 XOR Logical_Operator_out360_out1;

  Logical_Operator_out3432_out1 <= in712 XOR in720;

  Logical_Operator_out3433_out1 <= Logical_Operator_out2409_out1 XOR Logical_Operator_out2413_out1;

  Logical_Operator_out3434_out1 <= Logical_Operator_out2410_out1 XOR Logical_Operator_out2414_out1;

  Logical_Operator_out3435_out1 <= Logical_Operator_out2411_out1 XOR Logical_Operator_out2415_out1;

  Logical_Operator_out3436_out1 <= Logical_Operator_out2412_out1 XOR Logical_Operator_out2416_out1;

  Logical_Operator_out3437_out1 <= Logical_Operator_out1387_out1 XOR Logical_Operator_out1391_out1;

  Logical_Operator_out3438_out1 <= Logical_Operator_out1388_out1 XOR Logical_Operator_out1392_out1;

  Logical_Operator_out3439_out1 <= Logical_Operator_out364_out1 XOR Logical_Operator_out368_out1;

  Logical_Operator_out3440_out1 <= in728 XOR in736;

  Logical_Operator_out3441_out1 <= Logical_Operator_out2417_out1 XOR Logical_Operator_out2421_out1;

  Logical_Operator_out3442_out1 <= Logical_Operator_out2418_out1 XOR Logical_Operator_out2422_out1;

  Logical_Operator_out3443_out1 <= Logical_Operator_out2419_out1 XOR Logical_Operator_out2423_out1;

  Logical_Operator_out3444_out1 <= Logical_Operator_out2420_out1 XOR Logical_Operator_out2424_out1;

  Logical_Operator_out3445_out1 <= Logical_Operator_out1395_out1 XOR Logical_Operator_out1399_out1;

  Logical_Operator_out3446_out1 <= Logical_Operator_out1396_out1 XOR Logical_Operator_out1400_out1;

  Logical_Operator_out3447_out1 <= Logical_Operator_out372_out1 XOR Logical_Operator_out376_out1;

  Logical_Operator_out3448_out1 <= in744 XOR in752;

  Logical_Operator_out3449_out1 <= Logical_Operator_out2425_out1 XOR Logical_Operator_out2429_out1;

  Logical_Operator_out3450_out1 <= Logical_Operator_out2426_out1 XOR Logical_Operator_out2430_out1;

  Logical_Operator_out3451_out1 <= Logical_Operator_out2427_out1 XOR Logical_Operator_out2431_out1;

  Logical_Operator_out3452_out1 <= Logical_Operator_out2428_out1 XOR Logical_Operator_out2432_out1;

  Logical_Operator_out3453_out1 <= Logical_Operator_out1403_out1 XOR Logical_Operator_out1407_out1;

  Logical_Operator_out3454_out1 <= Logical_Operator_out1404_out1 XOR Logical_Operator_out1408_out1;

  Logical_Operator_out3455_out1 <= Logical_Operator_out380_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out3456_out1 <= in760 XOR in768;

  Logical_Operator_out3457_out1 <= Logical_Operator_out2433_out1 XOR Logical_Operator_out2437_out1;

  Logical_Operator_out3458_out1 <= Logical_Operator_out2434_out1 XOR Logical_Operator_out2438_out1;

  Logical_Operator_out3459_out1 <= Logical_Operator_out2435_out1 XOR Logical_Operator_out2439_out1;

  Logical_Operator_out3460_out1 <= Logical_Operator_out2436_out1 XOR Logical_Operator_out2440_out1;

  Logical_Operator_out3461_out1 <= Logical_Operator_out1411_out1 XOR Logical_Operator_out1415_out1;

  Logical_Operator_out3462_out1 <= Logical_Operator_out1412_out1 XOR Logical_Operator_out1416_out1;

  Logical_Operator_out3463_out1 <= Logical_Operator_out388_out1 XOR Logical_Operator_out392_out1;

  Logical_Operator_out3464_out1 <= in776 XOR in784;

  Logical_Operator_out3465_out1 <= Logical_Operator_out2441_out1 XOR Logical_Operator_out2445_out1;

  Logical_Operator_out3466_out1 <= Logical_Operator_out2442_out1 XOR Logical_Operator_out2446_out1;

  Logical_Operator_out3467_out1 <= Logical_Operator_out2443_out1 XOR Logical_Operator_out2447_out1;

  Logical_Operator_out3468_out1 <= Logical_Operator_out2444_out1 XOR Logical_Operator_out2448_out1;

  Logical_Operator_out3469_out1 <= Logical_Operator_out1419_out1 XOR Logical_Operator_out1423_out1;

  Logical_Operator_out3470_out1 <= Logical_Operator_out1420_out1 XOR Logical_Operator_out1424_out1;

  Logical_Operator_out3471_out1 <= Logical_Operator_out396_out1 XOR Logical_Operator_out400_out1;

  Logical_Operator_out3472_out1 <= in792 XOR in800;

  Logical_Operator_out3473_out1 <= Logical_Operator_out2449_out1 XOR Logical_Operator_out2453_out1;

  Logical_Operator_out3474_out1 <= Logical_Operator_out2450_out1 XOR Logical_Operator_out2454_out1;

  Logical_Operator_out3475_out1 <= Logical_Operator_out2451_out1 XOR Logical_Operator_out2455_out1;

  Logical_Operator_out3476_out1 <= Logical_Operator_out2452_out1 XOR Logical_Operator_out2456_out1;

  Logical_Operator_out3477_out1 <= Logical_Operator_out1427_out1 XOR Logical_Operator_out1431_out1;

  Logical_Operator_out3478_out1 <= Logical_Operator_out1428_out1 XOR Logical_Operator_out1432_out1;

  Logical_Operator_out3479_out1 <= Logical_Operator_out404_out1 XOR Logical_Operator_out408_out1;

  Logical_Operator_out3480_out1 <= in808 XOR in816;

  Logical_Operator_out3481_out1 <= Logical_Operator_out2457_out1 XOR Logical_Operator_out2461_out1;

  Logical_Operator_out3482_out1 <= Logical_Operator_out2458_out1 XOR Logical_Operator_out2462_out1;

  Logical_Operator_out3483_out1 <= Logical_Operator_out2459_out1 XOR Logical_Operator_out2463_out1;

  Logical_Operator_out3484_out1 <= Logical_Operator_out2460_out1 XOR Logical_Operator_out2464_out1;

  Logical_Operator_out3485_out1 <= Logical_Operator_out1435_out1 XOR Logical_Operator_out1439_out1;

  Logical_Operator_out3486_out1 <= Logical_Operator_out1436_out1 XOR Logical_Operator_out1440_out1;

  Logical_Operator_out3487_out1 <= Logical_Operator_out412_out1 XOR Logical_Operator_out416_out1;

  Logical_Operator_out3488_out1 <= in824 XOR in832;

  Logical_Operator_out3489_out1 <= Logical_Operator_out2465_out1 XOR Logical_Operator_out2469_out1;

  Logical_Operator_out3490_out1 <= Logical_Operator_out2466_out1 XOR Logical_Operator_out2470_out1;

  Logical_Operator_out3491_out1 <= Logical_Operator_out2467_out1 XOR Logical_Operator_out2471_out1;

  Logical_Operator_out3492_out1 <= Logical_Operator_out2468_out1 XOR Logical_Operator_out2472_out1;

  Logical_Operator_out3493_out1 <= Logical_Operator_out1443_out1 XOR Logical_Operator_out1447_out1;

  Logical_Operator_out3494_out1 <= Logical_Operator_out1444_out1 XOR Logical_Operator_out1448_out1;

  Logical_Operator_out3495_out1 <= Logical_Operator_out420_out1 XOR Logical_Operator_out424_out1;

  Logical_Operator_out3496_out1 <= in840 XOR in848;

  Logical_Operator_out3497_out1 <= Logical_Operator_out2473_out1 XOR Logical_Operator_out2477_out1;

  Logical_Operator_out3498_out1 <= Logical_Operator_out2474_out1 XOR Logical_Operator_out2478_out1;

  Logical_Operator_out3499_out1 <= Logical_Operator_out2475_out1 XOR Logical_Operator_out2479_out1;

  Logical_Operator_out3500_out1 <= Logical_Operator_out2476_out1 XOR Logical_Operator_out2480_out1;

  Logical_Operator_out3501_out1 <= Logical_Operator_out1451_out1 XOR Logical_Operator_out1455_out1;

  Logical_Operator_out3502_out1 <= Logical_Operator_out1452_out1 XOR Logical_Operator_out1456_out1;

  Logical_Operator_out3503_out1 <= Logical_Operator_out428_out1 XOR Logical_Operator_out432_out1;

  Logical_Operator_out3504_out1 <= in856 XOR in864;

  Logical_Operator_out3505_out1 <= Logical_Operator_out2481_out1 XOR Logical_Operator_out2485_out1;

  Logical_Operator_out3506_out1 <= Logical_Operator_out2482_out1 XOR Logical_Operator_out2486_out1;

  Logical_Operator_out3507_out1 <= Logical_Operator_out2483_out1 XOR Logical_Operator_out2487_out1;

  Logical_Operator_out3508_out1 <= Logical_Operator_out2484_out1 XOR Logical_Operator_out2488_out1;

  Logical_Operator_out3509_out1 <= Logical_Operator_out1459_out1 XOR Logical_Operator_out1463_out1;

  Logical_Operator_out3510_out1 <= Logical_Operator_out1460_out1 XOR Logical_Operator_out1464_out1;

  Logical_Operator_out3511_out1 <= Logical_Operator_out436_out1 XOR Logical_Operator_out440_out1;

  Logical_Operator_out3512_out1 <= in872 XOR in880;

  Logical_Operator_out3513_out1 <= Logical_Operator_out2489_out1 XOR Logical_Operator_out2493_out1;

  Logical_Operator_out3514_out1 <= Logical_Operator_out2490_out1 XOR Logical_Operator_out2494_out1;

  Logical_Operator_out3515_out1 <= Logical_Operator_out2491_out1 XOR Logical_Operator_out2495_out1;

  Logical_Operator_out3516_out1 <= Logical_Operator_out2492_out1 XOR Logical_Operator_out2496_out1;

  Logical_Operator_out3517_out1 <= Logical_Operator_out1467_out1 XOR Logical_Operator_out1471_out1;

  Logical_Operator_out3518_out1 <= Logical_Operator_out1468_out1 XOR Logical_Operator_out1472_out1;

  Logical_Operator_out3519_out1 <= Logical_Operator_out444_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out3520_out1 <= in888 XOR in896;

  Logical_Operator_out3521_out1 <= Logical_Operator_out2497_out1 XOR Logical_Operator_out2501_out1;

  Logical_Operator_out3522_out1 <= Logical_Operator_out2498_out1 XOR Logical_Operator_out2502_out1;

  Logical_Operator_out3523_out1 <= Logical_Operator_out2499_out1 XOR Logical_Operator_out2503_out1;

  Logical_Operator_out3524_out1 <= Logical_Operator_out2500_out1 XOR Logical_Operator_out2504_out1;

  Logical_Operator_out3525_out1 <= Logical_Operator_out1475_out1 XOR Logical_Operator_out1479_out1;

  Logical_Operator_out3526_out1 <= Logical_Operator_out1476_out1 XOR Logical_Operator_out1480_out1;

  Logical_Operator_out3527_out1 <= Logical_Operator_out452_out1 XOR Logical_Operator_out456_out1;

  Logical_Operator_out3528_out1 <= in904 XOR in912;

  Logical_Operator_out3529_out1 <= Logical_Operator_out2505_out1 XOR Logical_Operator_out2509_out1;

  Logical_Operator_out3530_out1 <= Logical_Operator_out2506_out1 XOR Logical_Operator_out2510_out1;

  Logical_Operator_out3531_out1 <= Logical_Operator_out2507_out1 XOR Logical_Operator_out2511_out1;

  Logical_Operator_out3532_out1 <= Logical_Operator_out2508_out1 XOR Logical_Operator_out2512_out1;

  Logical_Operator_out3533_out1 <= Logical_Operator_out1483_out1 XOR Logical_Operator_out1487_out1;

  Logical_Operator_out3534_out1 <= Logical_Operator_out1484_out1 XOR Logical_Operator_out1488_out1;

  Logical_Operator_out3535_out1 <= Logical_Operator_out460_out1 XOR Logical_Operator_out464_out1;

  Logical_Operator_out3536_out1 <= in920 XOR in928;

  Logical_Operator_out3537_out1 <= Logical_Operator_out2513_out1 XOR Logical_Operator_out2517_out1;

  Logical_Operator_out3538_out1 <= Logical_Operator_out2514_out1 XOR Logical_Operator_out2518_out1;

  Logical_Operator_out3539_out1 <= Logical_Operator_out2515_out1 XOR Logical_Operator_out2519_out1;

  Logical_Operator_out3540_out1 <= Logical_Operator_out2516_out1 XOR Logical_Operator_out2520_out1;

  Logical_Operator_out3541_out1 <= Logical_Operator_out1491_out1 XOR Logical_Operator_out1495_out1;

  Logical_Operator_out3542_out1 <= Logical_Operator_out1492_out1 XOR Logical_Operator_out1496_out1;

  Logical_Operator_out3543_out1 <= Logical_Operator_out468_out1 XOR Logical_Operator_out472_out1;

  Logical_Operator_out3544_out1 <= in936 XOR in944;

  Logical_Operator_out3545_out1 <= Logical_Operator_out2521_out1 XOR Logical_Operator_out2525_out1;

  Logical_Operator_out3546_out1 <= Logical_Operator_out2522_out1 XOR Logical_Operator_out2526_out1;

  Logical_Operator_out3547_out1 <= Logical_Operator_out2523_out1 XOR Logical_Operator_out2527_out1;

  Logical_Operator_out3548_out1 <= Logical_Operator_out2524_out1 XOR Logical_Operator_out2528_out1;

  Logical_Operator_out3549_out1 <= Logical_Operator_out1499_out1 XOR Logical_Operator_out1503_out1;

  Logical_Operator_out3550_out1 <= Logical_Operator_out1500_out1 XOR Logical_Operator_out1504_out1;

  Logical_Operator_out3551_out1 <= Logical_Operator_out476_out1 XOR Logical_Operator_out480_out1;

  Logical_Operator_out3552_out1 <= in952 XOR in960;

  Logical_Operator_out3553_out1 <= Logical_Operator_out2529_out1 XOR Logical_Operator_out2533_out1;

  Logical_Operator_out3554_out1 <= Logical_Operator_out2530_out1 XOR Logical_Operator_out2534_out1;

  Logical_Operator_out3555_out1 <= Logical_Operator_out2531_out1 XOR Logical_Operator_out2535_out1;

  Logical_Operator_out3556_out1 <= Logical_Operator_out2532_out1 XOR Logical_Operator_out2536_out1;

  Logical_Operator_out3557_out1 <= Logical_Operator_out1507_out1 XOR Logical_Operator_out1511_out1;

  Logical_Operator_out3558_out1 <= Logical_Operator_out1508_out1 XOR Logical_Operator_out1512_out1;

  Logical_Operator_out3559_out1 <= Logical_Operator_out484_out1 XOR Logical_Operator_out488_out1;

  Logical_Operator_out3560_out1 <= in968 XOR in976;

  Logical_Operator_out3561_out1 <= Logical_Operator_out2537_out1 XOR Logical_Operator_out2541_out1;

  Logical_Operator_out3562_out1 <= Logical_Operator_out2538_out1 XOR Logical_Operator_out2542_out1;

  Logical_Operator_out3563_out1 <= Logical_Operator_out2539_out1 XOR Logical_Operator_out2543_out1;

  Logical_Operator_out3564_out1 <= Logical_Operator_out2540_out1 XOR Logical_Operator_out2544_out1;

  Logical_Operator_out3565_out1 <= Logical_Operator_out1515_out1 XOR Logical_Operator_out1519_out1;

  Logical_Operator_out3566_out1 <= Logical_Operator_out1516_out1 XOR Logical_Operator_out1520_out1;

  Logical_Operator_out3567_out1 <= Logical_Operator_out492_out1 XOR Logical_Operator_out496_out1;

  Logical_Operator_out3568_out1 <= in984 XOR in992;

  Logical_Operator_out3569_out1 <= Logical_Operator_out2545_out1 XOR Logical_Operator_out2549_out1;

  Logical_Operator_out3570_out1 <= Logical_Operator_out2546_out1 XOR Logical_Operator_out2550_out1;

  Logical_Operator_out3571_out1 <= Logical_Operator_out2547_out1 XOR Logical_Operator_out2551_out1;

  Logical_Operator_out3572_out1 <= Logical_Operator_out2548_out1 XOR Logical_Operator_out2552_out1;

  Logical_Operator_out3573_out1 <= Logical_Operator_out1523_out1 XOR Logical_Operator_out1527_out1;

  Logical_Operator_out3574_out1 <= Logical_Operator_out1524_out1 XOR Logical_Operator_out1528_out1;

  Logical_Operator_out3575_out1 <= Logical_Operator_out500_out1 XOR Logical_Operator_out504_out1;

  Logical_Operator_out3576_out1 <= in1000 XOR in1008;

  Logical_Operator_out3577_out1 <= Logical_Operator_out2553_out1 XOR Logical_Operator_out2557_out1;

  Logical_Operator_out3578_out1 <= Logical_Operator_out2554_out1 XOR Logical_Operator_out2558_out1;

  Logical_Operator_out3579_out1 <= Logical_Operator_out2555_out1 XOR Logical_Operator_out2559_out1;

  Logical_Operator_out3580_out1 <= Logical_Operator_out2556_out1 XOR Logical_Operator_out2560_out1;

  Logical_Operator_out3581_out1 <= Logical_Operator_out1531_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out3582_out1 <= Logical_Operator_out1532_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out3583_out1 <= Logical_Operator_out508_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out3584_out1 <= in1016 XOR in1024;

  Logical_Operator_out3585_out1 <= Logical_Operator_out2561_out1 XOR Logical_Operator_out2565_out1;

  Logical_Operator_out3586_out1 <= Logical_Operator_out2562_out1 XOR Logical_Operator_out2566_out1;

  Logical_Operator_out3587_out1 <= Logical_Operator_out2563_out1 XOR Logical_Operator_out2567_out1;

  Logical_Operator_out3588_out1 <= Logical_Operator_out2564_out1 XOR Logical_Operator_out2568_out1;

  Logical_Operator_out3589_out1 <= Logical_Operator_out1539_out1 XOR Logical_Operator_out1543_out1;

  Logical_Operator_out3590_out1 <= Logical_Operator_out1540_out1 XOR Logical_Operator_out1544_out1;

  Logical_Operator_out3591_out1 <= Logical_Operator_out516_out1 XOR Logical_Operator_out520_out1;

  Logical_Operator_out3592_out1 <= in1032 XOR in1040;

  Logical_Operator_out3593_out1 <= Logical_Operator_out2569_out1 XOR Logical_Operator_out2573_out1;

  Logical_Operator_out3594_out1 <= Logical_Operator_out2570_out1 XOR Logical_Operator_out2574_out1;

  Logical_Operator_out3595_out1 <= Logical_Operator_out2571_out1 XOR Logical_Operator_out2575_out1;

  Logical_Operator_out3596_out1 <= Logical_Operator_out2572_out1 XOR Logical_Operator_out2576_out1;

  Logical_Operator_out3597_out1 <= Logical_Operator_out1547_out1 XOR Logical_Operator_out1551_out1;

  Logical_Operator_out3598_out1 <= Logical_Operator_out1548_out1 XOR Logical_Operator_out1552_out1;

  Logical_Operator_out3599_out1 <= Logical_Operator_out524_out1 XOR Logical_Operator_out528_out1;

  Logical_Operator_out3600_out1 <= in1048 XOR in1056;

  Logical_Operator_out3601_out1 <= Logical_Operator_out2577_out1 XOR Logical_Operator_out2581_out1;

  Logical_Operator_out3602_out1 <= Logical_Operator_out2578_out1 XOR Logical_Operator_out2582_out1;

  Logical_Operator_out3603_out1 <= Logical_Operator_out2579_out1 XOR Logical_Operator_out2583_out1;

  Logical_Operator_out3604_out1 <= Logical_Operator_out2580_out1 XOR Logical_Operator_out2584_out1;

  Logical_Operator_out3605_out1 <= Logical_Operator_out1555_out1 XOR Logical_Operator_out1559_out1;

  Logical_Operator_out3606_out1 <= Logical_Operator_out1556_out1 XOR Logical_Operator_out1560_out1;

  Logical_Operator_out3607_out1 <= Logical_Operator_out532_out1 XOR Logical_Operator_out536_out1;

  Logical_Operator_out3608_out1 <= in1064 XOR in1072;

  Logical_Operator_out3609_out1 <= Logical_Operator_out2585_out1 XOR Logical_Operator_out2589_out1;

  Logical_Operator_out3610_out1 <= Logical_Operator_out2586_out1 XOR Logical_Operator_out2590_out1;

  Logical_Operator_out3611_out1 <= Logical_Operator_out2587_out1 XOR Logical_Operator_out2591_out1;

  Logical_Operator_out3612_out1 <= Logical_Operator_out2588_out1 XOR Logical_Operator_out2592_out1;

  Logical_Operator_out3613_out1 <= Logical_Operator_out1563_out1 XOR Logical_Operator_out1567_out1;

  Logical_Operator_out3614_out1 <= Logical_Operator_out1564_out1 XOR Logical_Operator_out1568_out1;

  Logical_Operator_out3615_out1 <= Logical_Operator_out540_out1 XOR Logical_Operator_out544_out1;

  Logical_Operator_out3616_out1 <= in1080 XOR in1088;

  Logical_Operator_out3617_out1 <= Logical_Operator_out2593_out1 XOR Logical_Operator_out2597_out1;

  Logical_Operator_out3618_out1 <= Logical_Operator_out2594_out1 XOR Logical_Operator_out2598_out1;

  Logical_Operator_out3619_out1 <= Logical_Operator_out2595_out1 XOR Logical_Operator_out2599_out1;

  Logical_Operator_out3620_out1 <= Logical_Operator_out2596_out1 XOR Logical_Operator_out2600_out1;

  Logical_Operator_out3621_out1 <= Logical_Operator_out1571_out1 XOR Logical_Operator_out1575_out1;

  Logical_Operator_out3622_out1 <= Logical_Operator_out1572_out1 XOR Logical_Operator_out1576_out1;

  Logical_Operator_out3623_out1 <= Logical_Operator_out548_out1 XOR Logical_Operator_out552_out1;

  Logical_Operator_out3624_out1 <= in1096 XOR in1104;

  Logical_Operator_out3625_out1 <= Logical_Operator_out2601_out1 XOR Logical_Operator_out2605_out1;

  Logical_Operator_out3626_out1 <= Logical_Operator_out2602_out1 XOR Logical_Operator_out2606_out1;

  Logical_Operator_out3627_out1 <= Logical_Operator_out2603_out1 XOR Logical_Operator_out2607_out1;

  Logical_Operator_out3628_out1 <= Logical_Operator_out2604_out1 XOR Logical_Operator_out2608_out1;

  Logical_Operator_out3629_out1 <= Logical_Operator_out1579_out1 XOR Logical_Operator_out1583_out1;

  Logical_Operator_out3630_out1 <= Logical_Operator_out1580_out1 XOR Logical_Operator_out1584_out1;

  Logical_Operator_out3631_out1 <= Logical_Operator_out556_out1 XOR Logical_Operator_out560_out1;

  Logical_Operator_out3632_out1 <= in1112 XOR in1120;

  Logical_Operator_out3633_out1 <= Logical_Operator_out2609_out1 XOR Logical_Operator_out2613_out1;

  Logical_Operator_out3634_out1 <= Logical_Operator_out2610_out1 XOR Logical_Operator_out2614_out1;

  Logical_Operator_out3635_out1 <= Logical_Operator_out2611_out1 XOR Logical_Operator_out2615_out1;

  Logical_Operator_out3636_out1 <= Logical_Operator_out2612_out1 XOR Logical_Operator_out2616_out1;

  Logical_Operator_out3637_out1 <= Logical_Operator_out1587_out1 XOR Logical_Operator_out1591_out1;

  Logical_Operator_out3638_out1 <= Logical_Operator_out1588_out1 XOR Logical_Operator_out1592_out1;

  Logical_Operator_out3639_out1 <= Logical_Operator_out564_out1 XOR Logical_Operator_out568_out1;

  Logical_Operator_out3640_out1 <= in1128 XOR in1136;

  Logical_Operator_out3641_out1 <= Logical_Operator_out2617_out1 XOR Logical_Operator_out2621_out1;

  Logical_Operator_out3642_out1 <= Logical_Operator_out2618_out1 XOR Logical_Operator_out2622_out1;

  Logical_Operator_out3643_out1 <= Logical_Operator_out2619_out1 XOR Logical_Operator_out2623_out1;

  Logical_Operator_out3644_out1 <= Logical_Operator_out2620_out1 XOR Logical_Operator_out2624_out1;

  Logical_Operator_out3645_out1 <= Logical_Operator_out1595_out1 XOR Logical_Operator_out1599_out1;

  Logical_Operator_out3646_out1 <= Logical_Operator_out1596_out1 XOR Logical_Operator_out1600_out1;

  Logical_Operator_out3647_out1 <= Logical_Operator_out572_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out3648_out1 <= in1144 XOR in1152;

  Logical_Operator_out3649_out1 <= Logical_Operator_out2625_out1 XOR Logical_Operator_out2629_out1;

  Logical_Operator_out3650_out1 <= Logical_Operator_out2626_out1 XOR Logical_Operator_out2630_out1;

  Logical_Operator_out3651_out1 <= Logical_Operator_out2627_out1 XOR Logical_Operator_out2631_out1;

  Logical_Operator_out3652_out1 <= Logical_Operator_out2628_out1 XOR Logical_Operator_out2632_out1;

  Logical_Operator_out3653_out1 <= Logical_Operator_out1603_out1 XOR Logical_Operator_out1607_out1;

  Logical_Operator_out3654_out1 <= Logical_Operator_out1604_out1 XOR Logical_Operator_out1608_out1;

  Logical_Operator_out3655_out1 <= Logical_Operator_out580_out1 XOR Logical_Operator_out584_out1;

  Logical_Operator_out3656_out1 <= in1160 XOR in1168;

  Logical_Operator_out3657_out1 <= Logical_Operator_out2633_out1 XOR Logical_Operator_out2637_out1;

  Logical_Operator_out3658_out1 <= Logical_Operator_out2634_out1 XOR Logical_Operator_out2638_out1;

  Logical_Operator_out3659_out1 <= Logical_Operator_out2635_out1 XOR Logical_Operator_out2639_out1;

  Logical_Operator_out3660_out1 <= Logical_Operator_out2636_out1 XOR Logical_Operator_out2640_out1;

  Logical_Operator_out3661_out1 <= Logical_Operator_out1611_out1 XOR Logical_Operator_out1615_out1;

  Logical_Operator_out3662_out1 <= Logical_Operator_out1612_out1 XOR Logical_Operator_out1616_out1;

  Logical_Operator_out3663_out1 <= Logical_Operator_out588_out1 XOR Logical_Operator_out592_out1;

  Logical_Operator_out3664_out1 <= in1176 XOR in1184;

  Logical_Operator_out3665_out1 <= Logical_Operator_out2641_out1 XOR Logical_Operator_out2645_out1;

  Logical_Operator_out3666_out1 <= Logical_Operator_out2642_out1 XOR Logical_Operator_out2646_out1;

  Logical_Operator_out3667_out1 <= Logical_Operator_out2643_out1 XOR Logical_Operator_out2647_out1;

  Logical_Operator_out3668_out1 <= Logical_Operator_out2644_out1 XOR Logical_Operator_out2648_out1;

  Logical_Operator_out3669_out1 <= Logical_Operator_out1619_out1 XOR Logical_Operator_out1623_out1;

  Logical_Operator_out3670_out1 <= Logical_Operator_out1620_out1 XOR Logical_Operator_out1624_out1;

  Logical_Operator_out3671_out1 <= Logical_Operator_out596_out1 XOR Logical_Operator_out600_out1;

  Logical_Operator_out3672_out1 <= in1192 XOR in1200;

  Logical_Operator_out3673_out1 <= Logical_Operator_out2649_out1 XOR Logical_Operator_out2653_out1;

  Logical_Operator_out3674_out1 <= Logical_Operator_out2650_out1 XOR Logical_Operator_out2654_out1;

  Logical_Operator_out3675_out1 <= Logical_Operator_out2651_out1 XOR Logical_Operator_out2655_out1;

  Logical_Operator_out3676_out1 <= Logical_Operator_out2652_out1 XOR Logical_Operator_out2656_out1;

  Logical_Operator_out3677_out1 <= Logical_Operator_out1627_out1 XOR Logical_Operator_out1631_out1;

  Logical_Operator_out3678_out1 <= Logical_Operator_out1628_out1 XOR Logical_Operator_out1632_out1;

  Logical_Operator_out3679_out1 <= Logical_Operator_out604_out1 XOR Logical_Operator_out608_out1;

  Logical_Operator_out3680_out1 <= in1208 XOR in1216;

  Logical_Operator_out3681_out1 <= Logical_Operator_out2657_out1 XOR Logical_Operator_out2661_out1;

  Logical_Operator_out3682_out1 <= Logical_Operator_out2658_out1 XOR Logical_Operator_out2662_out1;

  Logical_Operator_out3683_out1 <= Logical_Operator_out2659_out1 XOR Logical_Operator_out2663_out1;

  Logical_Operator_out3684_out1 <= Logical_Operator_out2660_out1 XOR Logical_Operator_out2664_out1;

  Logical_Operator_out3685_out1 <= Logical_Operator_out1635_out1 XOR Logical_Operator_out1639_out1;

  Logical_Operator_out3686_out1 <= Logical_Operator_out1636_out1 XOR Logical_Operator_out1640_out1;

  Logical_Operator_out3687_out1 <= Logical_Operator_out612_out1 XOR Logical_Operator_out616_out1;

  Logical_Operator_out3688_out1 <= in1224 XOR in1232;

  Logical_Operator_out3689_out1 <= Logical_Operator_out2665_out1 XOR Logical_Operator_out2669_out1;

  Logical_Operator_out3690_out1 <= Logical_Operator_out2666_out1 XOR Logical_Operator_out2670_out1;

  Logical_Operator_out3691_out1 <= Logical_Operator_out2667_out1 XOR Logical_Operator_out2671_out1;

  Logical_Operator_out3692_out1 <= Logical_Operator_out2668_out1 XOR Logical_Operator_out2672_out1;

  Logical_Operator_out3693_out1 <= Logical_Operator_out1643_out1 XOR Logical_Operator_out1647_out1;

  Logical_Operator_out3694_out1 <= Logical_Operator_out1644_out1 XOR Logical_Operator_out1648_out1;

  Logical_Operator_out3695_out1 <= Logical_Operator_out620_out1 XOR Logical_Operator_out624_out1;

  Logical_Operator_out3696_out1 <= in1240 XOR in1248;

  Logical_Operator_out3697_out1 <= Logical_Operator_out2673_out1 XOR Logical_Operator_out2677_out1;

  Logical_Operator_out3698_out1 <= Logical_Operator_out2674_out1 XOR Logical_Operator_out2678_out1;

  Logical_Operator_out3699_out1 <= Logical_Operator_out2675_out1 XOR Logical_Operator_out2679_out1;

  Logical_Operator_out3700_out1 <= Logical_Operator_out2676_out1 XOR Logical_Operator_out2680_out1;

  Logical_Operator_out3701_out1 <= Logical_Operator_out1651_out1 XOR Logical_Operator_out1655_out1;

  Logical_Operator_out3702_out1 <= Logical_Operator_out1652_out1 XOR Logical_Operator_out1656_out1;

  Logical_Operator_out3703_out1 <= Logical_Operator_out628_out1 XOR Logical_Operator_out632_out1;

  Logical_Operator_out3704_out1 <= in1256 XOR in1264;

  Logical_Operator_out3705_out1 <= Logical_Operator_out2681_out1 XOR Logical_Operator_out2685_out1;

  Logical_Operator_out3706_out1 <= Logical_Operator_out2682_out1 XOR Logical_Operator_out2686_out1;

  Logical_Operator_out3707_out1 <= Logical_Operator_out2683_out1 XOR Logical_Operator_out2687_out1;

  Logical_Operator_out3708_out1 <= Logical_Operator_out2684_out1 XOR Logical_Operator_out2688_out1;

  Logical_Operator_out3709_out1 <= Logical_Operator_out1659_out1 XOR Logical_Operator_out1663_out1;

  Logical_Operator_out3710_out1 <= Logical_Operator_out1660_out1 XOR Logical_Operator_out1664_out1;

  Logical_Operator_out3711_out1 <= Logical_Operator_out636_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out3712_out1 <= in1272 XOR in1280;

  Logical_Operator_out3713_out1 <= Logical_Operator_out2689_out1 XOR Logical_Operator_out2693_out1;

  Logical_Operator_out3714_out1 <= Logical_Operator_out2690_out1 XOR Logical_Operator_out2694_out1;

  Logical_Operator_out3715_out1 <= Logical_Operator_out2691_out1 XOR Logical_Operator_out2695_out1;

  Logical_Operator_out3716_out1 <= Logical_Operator_out2692_out1 XOR Logical_Operator_out2696_out1;

  Logical_Operator_out3717_out1 <= Logical_Operator_out1667_out1 XOR Logical_Operator_out1671_out1;

  Logical_Operator_out3718_out1 <= Logical_Operator_out1668_out1 XOR Logical_Operator_out1672_out1;

  Logical_Operator_out3719_out1 <= Logical_Operator_out644_out1 XOR Logical_Operator_out648_out1;

  Logical_Operator_out3720_out1 <= in1288 XOR in1296;

  Logical_Operator_out3721_out1 <= Logical_Operator_out2697_out1 XOR Logical_Operator_out2701_out1;

  Logical_Operator_out3722_out1 <= Logical_Operator_out2698_out1 XOR Logical_Operator_out2702_out1;

  Logical_Operator_out3723_out1 <= Logical_Operator_out2699_out1 XOR Logical_Operator_out2703_out1;

  Logical_Operator_out3724_out1 <= Logical_Operator_out2700_out1 XOR Logical_Operator_out2704_out1;

  Logical_Operator_out3725_out1 <= Logical_Operator_out1675_out1 XOR Logical_Operator_out1679_out1;

  Logical_Operator_out3726_out1 <= Logical_Operator_out1676_out1 XOR Logical_Operator_out1680_out1;

  Logical_Operator_out3727_out1 <= Logical_Operator_out652_out1 XOR Logical_Operator_out656_out1;

  Logical_Operator_out3728_out1 <= in1304 XOR in1312;

  Logical_Operator_out3729_out1 <= Logical_Operator_out2705_out1 XOR Logical_Operator_out2709_out1;

  Logical_Operator_out3730_out1 <= Logical_Operator_out2706_out1 XOR Logical_Operator_out2710_out1;

  Logical_Operator_out3731_out1 <= Logical_Operator_out2707_out1 XOR Logical_Operator_out2711_out1;

  Logical_Operator_out3732_out1 <= Logical_Operator_out2708_out1 XOR Logical_Operator_out2712_out1;

  Logical_Operator_out3733_out1 <= Logical_Operator_out1683_out1 XOR Logical_Operator_out1687_out1;

  Logical_Operator_out3734_out1 <= Logical_Operator_out1684_out1 XOR Logical_Operator_out1688_out1;

  Logical_Operator_out3735_out1 <= Logical_Operator_out660_out1 XOR Logical_Operator_out664_out1;

  Logical_Operator_out3736_out1 <= in1320 XOR in1328;

  Logical_Operator_out3737_out1 <= Logical_Operator_out2713_out1 XOR Logical_Operator_out2717_out1;

  Logical_Operator_out3738_out1 <= Logical_Operator_out2714_out1 XOR Logical_Operator_out2718_out1;

  Logical_Operator_out3739_out1 <= Logical_Operator_out2715_out1 XOR Logical_Operator_out2719_out1;

  Logical_Operator_out3740_out1 <= Logical_Operator_out2716_out1 XOR Logical_Operator_out2720_out1;

  Logical_Operator_out3741_out1 <= Logical_Operator_out1691_out1 XOR Logical_Operator_out1695_out1;

  Logical_Operator_out3742_out1 <= Logical_Operator_out1692_out1 XOR Logical_Operator_out1696_out1;

  Logical_Operator_out3743_out1 <= Logical_Operator_out668_out1 XOR Logical_Operator_out672_out1;

  Logical_Operator_out3744_out1 <= in1336 XOR in1344;

  Logical_Operator_out3745_out1 <= Logical_Operator_out2721_out1 XOR Logical_Operator_out2725_out1;

  Logical_Operator_out3746_out1 <= Logical_Operator_out2722_out1 XOR Logical_Operator_out2726_out1;

  Logical_Operator_out3747_out1 <= Logical_Operator_out2723_out1 XOR Logical_Operator_out2727_out1;

  Logical_Operator_out3748_out1 <= Logical_Operator_out2724_out1 XOR Logical_Operator_out2728_out1;

  Logical_Operator_out3749_out1 <= Logical_Operator_out1699_out1 XOR Logical_Operator_out1703_out1;

  Logical_Operator_out3750_out1 <= Logical_Operator_out1700_out1 XOR Logical_Operator_out1704_out1;

  Logical_Operator_out3751_out1 <= Logical_Operator_out676_out1 XOR Logical_Operator_out680_out1;

  Logical_Operator_out3752_out1 <= in1352 XOR in1360;

  Logical_Operator_out3753_out1 <= Logical_Operator_out2729_out1 XOR Logical_Operator_out2733_out1;

  Logical_Operator_out3754_out1 <= Logical_Operator_out2730_out1 XOR Logical_Operator_out2734_out1;

  Logical_Operator_out3755_out1 <= Logical_Operator_out2731_out1 XOR Logical_Operator_out2735_out1;

  Logical_Operator_out3756_out1 <= Logical_Operator_out2732_out1 XOR Logical_Operator_out2736_out1;

  Logical_Operator_out3757_out1 <= Logical_Operator_out1707_out1 XOR Logical_Operator_out1711_out1;

  Logical_Operator_out3758_out1 <= Logical_Operator_out1708_out1 XOR Logical_Operator_out1712_out1;

  Logical_Operator_out3759_out1 <= Logical_Operator_out684_out1 XOR Logical_Operator_out688_out1;

  Logical_Operator_out3760_out1 <= in1368 XOR in1376;

  Logical_Operator_out3761_out1 <= Logical_Operator_out2737_out1 XOR Logical_Operator_out2741_out1;

  Logical_Operator_out3762_out1 <= Logical_Operator_out2738_out1 XOR Logical_Operator_out2742_out1;

  Logical_Operator_out3763_out1 <= Logical_Operator_out2739_out1 XOR Logical_Operator_out2743_out1;

  Logical_Operator_out3764_out1 <= Logical_Operator_out2740_out1 XOR Logical_Operator_out2744_out1;

  Logical_Operator_out3765_out1 <= Logical_Operator_out1715_out1 XOR Logical_Operator_out1719_out1;

  Logical_Operator_out3766_out1 <= Logical_Operator_out1716_out1 XOR Logical_Operator_out1720_out1;

  Logical_Operator_out3767_out1 <= Logical_Operator_out692_out1 XOR Logical_Operator_out696_out1;

  Logical_Operator_out3768_out1 <= in1384 XOR in1392;

  Logical_Operator_out3769_out1 <= Logical_Operator_out2745_out1 XOR Logical_Operator_out2749_out1;

  Logical_Operator_out3770_out1 <= Logical_Operator_out2746_out1 XOR Logical_Operator_out2750_out1;

  Logical_Operator_out3771_out1 <= Logical_Operator_out2747_out1 XOR Logical_Operator_out2751_out1;

  Logical_Operator_out3772_out1 <= Logical_Operator_out2748_out1 XOR Logical_Operator_out2752_out1;

  Logical_Operator_out3773_out1 <= Logical_Operator_out1723_out1 XOR Logical_Operator_out1727_out1;

  Logical_Operator_out3774_out1 <= Logical_Operator_out1724_out1 XOR Logical_Operator_out1728_out1;

  Logical_Operator_out3775_out1 <= Logical_Operator_out700_out1 XOR Logical_Operator_out704_out1;

  Logical_Operator_out3776_out1 <= in1400 XOR in1408;

  Logical_Operator_out3777_out1 <= Logical_Operator_out2753_out1 XOR Logical_Operator_out2757_out1;

  Logical_Operator_out3778_out1 <= Logical_Operator_out2754_out1 XOR Logical_Operator_out2758_out1;

  Logical_Operator_out3779_out1 <= Logical_Operator_out2755_out1 XOR Logical_Operator_out2759_out1;

  Logical_Operator_out3780_out1 <= Logical_Operator_out2756_out1 XOR Logical_Operator_out2760_out1;

  Logical_Operator_out3781_out1 <= Logical_Operator_out1731_out1 XOR Logical_Operator_out1735_out1;

  Logical_Operator_out3782_out1 <= Logical_Operator_out1732_out1 XOR Logical_Operator_out1736_out1;

  Logical_Operator_out3783_out1 <= Logical_Operator_out708_out1 XOR Logical_Operator_out712_out1;

  Logical_Operator_out3784_out1 <= in1416 XOR in1424;

  Logical_Operator_out3785_out1 <= Logical_Operator_out2761_out1 XOR Logical_Operator_out2765_out1;

  Logical_Operator_out3786_out1 <= Logical_Operator_out2762_out1 XOR Logical_Operator_out2766_out1;

  Logical_Operator_out3787_out1 <= Logical_Operator_out2763_out1 XOR Logical_Operator_out2767_out1;

  Logical_Operator_out3788_out1 <= Logical_Operator_out2764_out1 XOR Logical_Operator_out2768_out1;

  Logical_Operator_out3789_out1 <= Logical_Operator_out1739_out1 XOR Logical_Operator_out1743_out1;

  Logical_Operator_out3790_out1 <= Logical_Operator_out1740_out1 XOR Logical_Operator_out1744_out1;

  Logical_Operator_out3791_out1 <= Logical_Operator_out716_out1 XOR Logical_Operator_out720_out1;

  Logical_Operator_out3792_out1 <= in1432 XOR in1440;

  Logical_Operator_out3793_out1 <= Logical_Operator_out2769_out1 XOR Logical_Operator_out2773_out1;

  Logical_Operator_out3794_out1 <= Logical_Operator_out2770_out1 XOR Logical_Operator_out2774_out1;

  Logical_Operator_out3795_out1 <= Logical_Operator_out2771_out1 XOR Logical_Operator_out2775_out1;

  Logical_Operator_out3796_out1 <= Logical_Operator_out2772_out1 XOR Logical_Operator_out2776_out1;

  Logical_Operator_out3797_out1 <= Logical_Operator_out1747_out1 XOR Logical_Operator_out1751_out1;

  Logical_Operator_out3798_out1 <= Logical_Operator_out1748_out1 XOR Logical_Operator_out1752_out1;

  Logical_Operator_out3799_out1 <= Logical_Operator_out724_out1 XOR Logical_Operator_out728_out1;

  Logical_Operator_out3800_out1 <= in1448 XOR in1456;

  Logical_Operator_out3801_out1 <= Logical_Operator_out2777_out1 XOR Logical_Operator_out2781_out1;

  Logical_Operator_out3802_out1 <= Logical_Operator_out2778_out1 XOR Logical_Operator_out2782_out1;

  Logical_Operator_out3803_out1 <= Logical_Operator_out2779_out1 XOR Logical_Operator_out2783_out1;

  Logical_Operator_out3804_out1 <= Logical_Operator_out2780_out1 XOR Logical_Operator_out2784_out1;

  Logical_Operator_out3805_out1 <= Logical_Operator_out1755_out1 XOR Logical_Operator_out1759_out1;

  Logical_Operator_out3806_out1 <= Logical_Operator_out1756_out1 XOR Logical_Operator_out1760_out1;

  Logical_Operator_out3807_out1 <= Logical_Operator_out732_out1 XOR Logical_Operator_out736_out1;

  Logical_Operator_out3808_out1 <= in1464 XOR in1472;

  Logical_Operator_out3809_out1 <= Logical_Operator_out2785_out1 XOR Logical_Operator_out2789_out1;

  Logical_Operator_out3810_out1 <= Logical_Operator_out2786_out1 XOR Logical_Operator_out2790_out1;

  Logical_Operator_out3811_out1 <= Logical_Operator_out2787_out1 XOR Logical_Operator_out2791_out1;

  Logical_Operator_out3812_out1 <= Logical_Operator_out2788_out1 XOR Logical_Operator_out2792_out1;

  Logical_Operator_out3813_out1 <= Logical_Operator_out1763_out1 XOR Logical_Operator_out1767_out1;

  Logical_Operator_out3814_out1 <= Logical_Operator_out1764_out1 XOR Logical_Operator_out1768_out1;

  Logical_Operator_out3815_out1 <= Logical_Operator_out740_out1 XOR Logical_Operator_out744_out1;

  Logical_Operator_out3816_out1 <= in1480 XOR in1488;

  Logical_Operator_out3817_out1 <= Logical_Operator_out2793_out1 XOR Logical_Operator_out2797_out1;

  Logical_Operator_out3818_out1 <= Logical_Operator_out2794_out1 XOR Logical_Operator_out2798_out1;

  Logical_Operator_out3819_out1 <= Logical_Operator_out2795_out1 XOR Logical_Operator_out2799_out1;

  Logical_Operator_out3820_out1 <= Logical_Operator_out2796_out1 XOR Logical_Operator_out2800_out1;

  Logical_Operator_out3821_out1 <= Logical_Operator_out1771_out1 XOR Logical_Operator_out1775_out1;

  Logical_Operator_out3822_out1 <= Logical_Operator_out1772_out1 XOR Logical_Operator_out1776_out1;

  Logical_Operator_out3823_out1 <= Logical_Operator_out748_out1 XOR Logical_Operator_out752_out1;

  Logical_Operator_out3824_out1 <= in1496 XOR in1504;

  Logical_Operator_out3825_out1 <= Logical_Operator_out2801_out1 XOR Logical_Operator_out2805_out1;

  Logical_Operator_out3826_out1 <= Logical_Operator_out2802_out1 XOR Logical_Operator_out2806_out1;

  Logical_Operator_out3827_out1 <= Logical_Operator_out2803_out1 XOR Logical_Operator_out2807_out1;

  Logical_Operator_out3828_out1 <= Logical_Operator_out2804_out1 XOR Logical_Operator_out2808_out1;

  Logical_Operator_out3829_out1 <= Logical_Operator_out1779_out1 XOR Logical_Operator_out1783_out1;

  Logical_Operator_out3830_out1 <= Logical_Operator_out1780_out1 XOR Logical_Operator_out1784_out1;

  Logical_Operator_out3831_out1 <= Logical_Operator_out756_out1 XOR Logical_Operator_out760_out1;

  Logical_Operator_out3832_out1 <= in1512 XOR in1520;

  Logical_Operator_out3833_out1 <= Logical_Operator_out2809_out1 XOR Logical_Operator_out2813_out1;

  Logical_Operator_out3834_out1 <= Logical_Operator_out2810_out1 XOR Logical_Operator_out2814_out1;

  Logical_Operator_out3835_out1 <= Logical_Operator_out2811_out1 XOR Logical_Operator_out2815_out1;

  Logical_Operator_out3836_out1 <= Logical_Operator_out2812_out1 XOR Logical_Operator_out2816_out1;

  Logical_Operator_out3837_out1 <= Logical_Operator_out1787_out1 XOR Logical_Operator_out1791_out1;

  Logical_Operator_out3838_out1 <= Logical_Operator_out1788_out1 XOR Logical_Operator_out1792_out1;

  Logical_Operator_out3839_out1 <= Logical_Operator_out764_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out3840_out1 <= in1528 XOR in1536;

  Logical_Operator_out3841_out1 <= Logical_Operator_out2817_out1 XOR Logical_Operator_out2821_out1;

  Logical_Operator_out3842_out1 <= Logical_Operator_out2818_out1 XOR Logical_Operator_out2822_out1;

  Logical_Operator_out3843_out1 <= Logical_Operator_out2819_out1 XOR Logical_Operator_out2823_out1;

  Logical_Operator_out3844_out1 <= Logical_Operator_out2820_out1 XOR Logical_Operator_out2824_out1;

  Logical_Operator_out3845_out1 <= Logical_Operator_out1795_out1 XOR Logical_Operator_out1799_out1;

  Logical_Operator_out3846_out1 <= Logical_Operator_out1796_out1 XOR Logical_Operator_out1800_out1;

  Logical_Operator_out3847_out1 <= Logical_Operator_out772_out1 XOR Logical_Operator_out776_out1;

  Logical_Operator_out3848_out1 <= in1544 XOR in1552;

  Logical_Operator_out3849_out1 <= Logical_Operator_out2825_out1 XOR Logical_Operator_out2829_out1;

  Logical_Operator_out3850_out1 <= Logical_Operator_out2826_out1 XOR Logical_Operator_out2830_out1;

  Logical_Operator_out3851_out1 <= Logical_Operator_out2827_out1 XOR Logical_Operator_out2831_out1;

  Logical_Operator_out3852_out1 <= Logical_Operator_out2828_out1 XOR Logical_Operator_out2832_out1;

  Logical_Operator_out3853_out1 <= Logical_Operator_out1803_out1 XOR Logical_Operator_out1807_out1;

  Logical_Operator_out3854_out1 <= Logical_Operator_out1804_out1 XOR Logical_Operator_out1808_out1;

  Logical_Operator_out3855_out1 <= Logical_Operator_out780_out1 XOR Logical_Operator_out784_out1;

  Logical_Operator_out3856_out1 <= in1560 XOR in1568;

  Logical_Operator_out3857_out1 <= Logical_Operator_out2833_out1 XOR Logical_Operator_out2837_out1;

  Logical_Operator_out3858_out1 <= Logical_Operator_out2834_out1 XOR Logical_Operator_out2838_out1;

  Logical_Operator_out3859_out1 <= Logical_Operator_out2835_out1 XOR Logical_Operator_out2839_out1;

  Logical_Operator_out3860_out1 <= Logical_Operator_out2836_out1 XOR Logical_Operator_out2840_out1;

  Logical_Operator_out3861_out1 <= Logical_Operator_out1811_out1 XOR Logical_Operator_out1815_out1;

  Logical_Operator_out3862_out1 <= Logical_Operator_out1812_out1 XOR Logical_Operator_out1816_out1;

  Logical_Operator_out3863_out1 <= Logical_Operator_out788_out1 XOR Logical_Operator_out792_out1;

  Logical_Operator_out3864_out1 <= in1576 XOR in1584;

  Logical_Operator_out3865_out1 <= Logical_Operator_out2841_out1 XOR Logical_Operator_out2845_out1;

  Logical_Operator_out3866_out1 <= Logical_Operator_out2842_out1 XOR Logical_Operator_out2846_out1;

  Logical_Operator_out3867_out1 <= Logical_Operator_out2843_out1 XOR Logical_Operator_out2847_out1;

  Logical_Operator_out3868_out1 <= Logical_Operator_out2844_out1 XOR Logical_Operator_out2848_out1;

  Logical_Operator_out3869_out1 <= Logical_Operator_out1819_out1 XOR Logical_Operator_out1823_out1;

  Logical_Operator_out3870_out1 <= Logical_Operator_out1820_out1 XOR Logical_Operator_out1824_out1;

  Logical_Operator_out3871_out1 <= Logical_Operator_out796_out1 XOR Logical_Operator_out800_out1;

  Logical_Operator_out3872_out1 <= in1592 XOR in1600;

  Logical_Operator_out3873_out1 <= Logical_Operator_out2849_out1 XOR Logical_Operator_out2853_out1;

  Logical_Operator_out3874_out1 <= Logical_Operator_out2850_out1 XOR Logical_Operator_out2854_out1;

  Logical_Operator_out3875_out1 <= Logical_Operator_out2851_out1 XOR Logical_Operator_out2855_out1;

  Logical_Operator_out3876_out1 <= Logical_Operator_out2852_out1 XOR Logical_Operator_out2856_out1;

  Logical_Operator_out3877_out1 <= Logical_Operator_out1827_out1 XOR Logical_Operator_out1831_out1;

  Logical_Operator_out3878_out1 <= Logical_Operator_out1828_out1 XOR Logical_Operator_out1832_out1;

  Logical_Operator_out3879_out1 <= Logical_Operator_out804_out1 XOR Logical_Operator_out808_out1;

  Logical_Operator_out3880_out1 <= in1608 XOR in1616;

  Logical_Operator_out3881_out1 <= Logical_Operator_out2857_out1 XOR Logical_Operator_out2861_out1;

  Logical_Operator_out3882_out1 <= Logical_Operator_out2858_out1 XOR Logical_Operator_out2862_out1;

  Logical_Operator_out3883_out1 <= Logical_Operator_out2859_out1 XOR Logical_Operator_out2863_out1;

  Logical_Operator_out3884_out1 <= Logical_Operator_out2860_out1 XOR Logical_Operator_out2864_out1;

  Logical_Operator_out3885_out1 <= Logical_Operator_out1835_out1 XOR Logical_Operator_out1839_out1;

  Logical_Operator_out3886_out1 <= Logical_Operator_out1836_out1 XOR Logical_Operator_out1840_out1;

  Logical_Operator_out3887_out1 <= Logical_Operator_out812_out1 XOR Logical_Operator_out816_out1;

  Logical_Operator_out3888_out1 <= in1624 XOR in1632;

  Logical_Operator_out3889_out1 <= Logical_Operator_out2865_out1 XOR Logical_Operator_out2869_out1;

  Logical_Operator_out3890_out1 <= Logical_Operator_out2866_out1 XOR Logical_Operator_out2870_out1;

  Logical_Operator_out3891_out1 <= Logical_Operator_out2867_out1 XOR Logical_Operator_out2871_out1;

  Logical_Operator_out3892_out1 <= Logical_Operator_out2868_out1 XOR Logical_Operator_out2872_out1;

  Logical_Operator_out3893_out1 <= Logical_Operator_out1843_out1 XOR Logical_Operator_out1847_out1;

  Logical_Operator_out3894_out1 <= Logical_Operator_out1844_out1 XOR Logical_Operator_out1848_out1;

  Logical_Operator_out3895_out1 <= Logical_Operator_out820_out1 XOR Logical_Operator_out824_out1;

  Logical_Operator_out3896_out1 <= in1640 XOR in1648;

  Logical_Operator_out3897_out1 <= Logical_Operator_out2873_out1 XOR Logical_Operator_out2877_out1;

  Logical_Operator_out3898_out1 <= Logical_Operator_out2874_out1 XOR Logical_Operator_out2878_out1;

  Logical_Operator_out3899_out1 <= Logical_Operator_out2875_out1 XOR Logical_Operator_out2879_out1;

  Logical_Operator_out3900_out1 <= Logical_Operator_out2876_out1 XOR Logical_Operator_out2880_out1;

  Logical_Operator_out3901_out1 <= Logical_Operator_out1851_out1 XOR Logical_Operator_out1855_out1;

  Logical_Operator_out3902_out1 <= Logical_Operator_out1852_out1 XOR Logical_Operator_out1856_out1;

  Logical_Operator_out3903_out1 <= Logical_Operator_out828_out1 XOR Logical_Operator_out832_out1;

  Logical_Operator_out3904_out1 <= in1656 XOR in1664;

  Logical_Operator_out3905_out1 <= Logical_Operator_out2881_out1 XOR Logical_Operator_out2885_out1;

  Logical_Operator_out3906_out1 <= Logical_Operator_out2882_out1 XOR Logical_Operator_out2886_out1;

  Logical_Operator_out3907_out1 <= Logical_Operator_out2883_out1 XOR Logical_Operator_out2887_out1;

  Logical_Operator_out3908_out1 <= Logical_Operator_out2884_out1 XOR Logical_Operator_out2888_out1;

  Logical_Operator_out3909_out1 <= Logical_Operator_out1859_out1 XOR Logical_Operator_out1863_out1;

  Logical_Operator_out3910_out1 <= Logical_Operator_out1860_out1 XOR Logical_Operator_out1864_out1;

  Logical_Operator_out3911_out1 <= Logical_Operator_out836_out1 XOR Logical_Operator_out840_out1;

  Logical_Operator_out3912_out1 <= in1672 XOR in1680;

  Logical_Operator_out3913_out1 <= Logical_Operator_out2889_out1 XOR Logical_Operator_out2893_out1;

  Logical_Operator_out3914_out1 <= Logical_Operator_out2890_out1 XOR Logical_Operator_out2894_out1;

  Logical_Operator_out3915_out1 <= Logical_Operator_out2891_out1 XOR Logical_Operator_out2895_out1;

  Logical_Operator_out3916_out1 <= Logical_Operator_out2892_out1 XOR Logical_Operator_out2896_out1;

  Logical_Operator_out3917_out1 <= Logical_Operator_out1867_out1 XOR Logical_Operator_out1871_out1;

  Logical_Operator_out3918_out1 <= Logical_Operator_out1868_out1 XOR Logical_Operator_out1872_out1;

  Logical_Operator_out3919_out1 <= Logical_Operator_out844_out1 XOR Logical_Operator_out848_out1;

  Logical_Operator_out3920_out1 <= in1688 XOR in1696;

  Logical_Operator_out3921_out1 <= Logical_Operator_out2897_out1 XOR Logical_Operator_out2901_out1;

  Logical_Operator_out3922_out1 <= Logical_Operator_out2898_out1 XOR Logical_Operator_out2902_out1;

  Logical_Operator_out3923_out1 <= Logical_Operator_out2899_out1 XOR Logical_Operator_out2903_out1;

  Logical_Operator_out3924_out1 <= Logical_Operator_out2900_out1 XOR Logical_Operator_out2904_out1;

  Logical_Operator_out3925_out1 <= Logical_Operator_out1875_out1 XOR Logical_Operator_out1879_out1;

  Logical_Operator_out3926_out1 <= Logical_Operator_out1876_out1 XOR Logical_Operator_out1880_out1;

  Logical_Operator_out3927_out1 <= Logical_Operator_out852_out1 XOR Logical_Operator_out856_out1;

  Logical_Operator_out3928_out1 <= in1704 XOR in1712;

  Logical_Operator_out3929_out1 <= Logical_Operator_out2905_out1 XOR Logical_Operator_out2909_out1;

  Logical_Operator_out3930_out1 <= Logical_Operator_out2906_out1 XOR Logical_Operator_out2910_out1;

  Logical_Operator_out3931_out1 <= Logical_Operator_out2907_out1 XOR Logical_Operator_out2911_out1;

  Logical_Operator_out3932_out1 <= Logical_Operator_out2908_out1 XOR Logical_Operator_out2912_out1;

  Logical_Operator_out3933_out1 <= Logical_Operator_out1883_out1 XOR Logical_Operator_out1887_out1;

  Logical_Operator_out3934_out1 <= Logical_Operator_out1884_out1 XOR Logical_Operator_out1888_out1;

  Logical_Operator_out3935_out1 <= Logical_Operator_out860_out1 XOR Logical_Operator_out864_out1;

  Logical_Operator_out3936_out1 <= in1720 XOR in1728;

  Logical_Operator_out3937_out1 <= Logical_Operator_out2913_out1 XOR Logical_Operator_out2917_out1;

  Logical_Operator_out3938_out1 <= Logical_Operator_out2914_out1 XOR Logical_Operator_out2918_out1;

  Logical_Operator_out3939_out1 <= Logical_Operator_out2915_out1 XOR Logical_Operator_out2919_out1;

  Logical_Operator_out3940_out1 <= Logical_Operator_out2916_out1 XOR Logical_Operator_out2920_out1;

  Logical_Operator_out3941_out1 <= Logical_Operator_out1891_out1 XOR Logical_Operator_out1895_out1;

  Logical_Operator_out3942_out1 <= Logical_Operator_out1892_out1 XOR Logical_Operator_out1896_out1;

  Logical_Operator_out3943_out1 <= Logical_Operator_out868_out1 XOR Logical_Operator_out872_out1;

  Logical_Operator_out3944_out1 <= in1736 XOR in1744;

  Logical_Operator_out3945_out1 <= Logical_Operator_out2921_out1 XOR Logical_Operator_out2925_out1;

  Logical_Operator_out3946_out1 <= Logical_Operator_out2922_out1 XOR Logical_Operator_out2926_out1;

  Logical_Operator_out3947_out1 <= Logical_Operator_out2923_out1 XOR Logical_Operator_out2927_out1;

  Logical_Operator_out3948_out1 <= Logical_Operator_out2924_out1 XOR Logical_Operator_out2928_out1;

  Logical_Operator_out3949_out1 <= Logical_Operator_out1899_out1 XOR Logical_Operator_out1903_out1;

  Logical_Operator_out3950_out1 <= Logical_Operator_out1900_out1 XOR Logical_Operator_out1904_out1;

  Logical_Operator_out3951_out1 <= Logical_Operator_out876_out1 XOR Logical_Operator_out880_out1;

  Logical_Operator_out3952_out1 <= in1752 XOR in1760;

  Logical_Operator_out3953_out1 <= Logical_Operator_out2929_out1 XOR Logical_Operator_out2933_out1;

  Logical_Operator_out3954_out1 <= Logical_Operator_out2930_out1 XOR Logical_Operator_out2934_out1;

  Logical_Operator_out3955_out1 <= Logical_Operator_out2931_out1 XOR Logical_Operator_out2935_out1;

  Logical_Operator_out3956_out1 <= Logical_Operator_out2932_out1 XOR Logical_Operator_out2936_out1;

  Logical_Operator_out3957_out1 <= Logical_Operator_out1907_out1 XOR Logical_Operator_out1911_out1;

  Logical_Operator_out3958_out1 <= Logical_Operator_out1908_out1 XOR Logical_Operator_out1912_out1;

  Logical_Operator_out3959_out1 <= Logical_Operator_out884_out1 XOR Logical_Operator_out888_out1;

  Logical_Operator_out3960_out1 <= in1768 XOR in1776;

  Logical_Operator_out3961_out1 <= Logical_Operator_out2937_out1 XOR Logical_Operator_out2941_out1;

  Logical_Operator_out3962_out1 <= Logical_Operator_out2938_out1 XOR Logical_Operator_out2942_out1;

  Logical_Operator_out3963_out1 <= Logical_Operator_out2939_out1 XOR Logical_Operator_out2943_out1;

  Logical_Operator_out3964_out1 <= Logical_Operator_out2940_out1 XOR Logical_Operator_out2944_out1;

  Logical_Operator_out3965_out1 <= Logical_Operator_out1915_out1 XOR Logical_Operator_out1919_out1;

  Logical_Operator_out3966_out1 <= Logical_Operator_out1916_out1 XOR Logical_Operator_out1920_out1;

  Logical_Operator_out3967_out1 <= Logical_Operator_out892_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out3968_out1 <= in1784 XOR in1792;

  Logical_Operator_out3969_out1 <= Logical_Operator_out2945_out1 XOR Logical_Operator_out2949_out1;

  Logical_Operator_out3970_out1 <= Logical_Operator_out2946_out1 XOR Logical_Operator_out2950_out1;

  Logical_Operator_out3971_out1 <= Logical_Operator_out2947_out1 XOR Logical_Operator_out2951_out1;

  Logical_Operator_out3972_out1 <= Logical_Operator_out2948_out1 XOR Logical_Operator_out2952_out1;

  Logical_Operator_out3973_out1 <= Logical_Operator_out1923_out1 XOR Logical_Operator_out1927_out1;

  Logical_Operator_out3974_out1 <= Logical_Operator_out1924_out1 XOR Logical_Operator_out1928_out1;

  Logical_Operator_out3975_out1 <= Logical_Operator_out900_out1 XOR Logical_Operator_out904_out1;

  Logical_Operator_out3976_out1 <= in1800 XOR in1808;

  Logical_Operator_out3977_out1 <= Logical_Operator_out2953_out1 XOR Logical_Operator_out2957_out1;

  Logical_Operator_out3978_out1 <= Logical_Operator_out2954_out1 XOR Logical_Operator_out2958_out1;

  Logical_Operator_out3979_out1 <= Logical_Operator_out2955_out1 XOR Logical_Operator_out2959_out1;

  Logical_Operator_out3980_out1 <= Logical_Operator_out2956_out1 XOR Logical_Operator_out2960_out1;

  Logical_Operator_out3981_out1 <= Logical_Operator_out1931_out1 XOR Logical_Operator_out1935_out1;

  Logical_Operator_out3982_out1 <= Logical_Operator_out1932_out1 XOR Logical_Operator_out1936_out1;

  Logical_Operator_out3983_out1 <= Logical_Operator_out908_out1 XOR Logical_Operator_out912_out1;

  Logical_Operator_out3984_out1 <= in1816 XOR in1824;

  Logical_Operator_out3985_out1 <= Logical_Operator_out2961_out1 XOR Logical_Operator_out2965_out1;

  Logical_Operator_out3986_out1 <= Logical_Operator_out2962_out1 XOR Logical_Operator_out2966_out1;

  Logical_Operator_out3987_out1 <= Logical_Operator_out2963_out1 XOR Logical_Operator_out2967_out1;

  Logical_Operator_out3988_out1 <= Logical_Operator_out2964_out1 XOR Logical_Operator_out2968_out1;

  Logical_Operator_out3989_out1 <= Logical_Operator_out1939_out1 XOR Logical_Operator_out1943_out1;

  Logical_Operator_out3990_out1 <= Logical_Operator_out1940_out1 XOR Logical_Operator_out1944_out1;

  Logical_Operator_out3991_out1 <= Logical_Operator_out916_out1 XOR Logical_Operator_out920_out1;

  Logical_Operator_out3992_out1 <= in1832 XOR in1840;

  Logical_Operator_out3993_out1 <= Logical_Operator_out2969_out1 XOR Logical_Operator_out2973_out1;

  Logical_Operator_out3994_out1 <= Logical_Operator_out2970_out1 XOR Logical_Operator_out2974_out1;

  Logical_Operator_out3995_out1 <= Logical_Operator_out2971_out1 XOR Logical_Operator_out2975_out1;

  Logical_Operator_out3996_out1 <= Logical_Operator_out2972_out1 XOR Logical_Operator_out2976_out1;

  Logical_Operator_out3997_out1 <= Logical_Operator_out1947_out1 XOR Logical_Operator_out1951_out1;

  Logical_Operator_out3998_out1 <= Logical_Operator_out1948_out1 XOR Logical_Operator_out1952_out1;

  Logical_Operator_out3999_out1 <= Logical_Operator_out924_out1 XOR Logical_Operator_out928_out1;

  Logical_Operator_out4000_out1 <= in1848 XOR in1856;

  Logical_Operator_out4001_out1 <= Logical_Operator_out2977_out1 XOR Logical_Operator_out2981_out1;

  Logical_Operator_out4002_out1 <= Logical_Operator_out2978_out1 XOR Logical_Operator_out2982_out1;

  Logical_Operator_out4003_out1 <= Logical_Operator_out2979_out1 XOR Logical_Operator_out2983_out1;

  Logical_Operator_out4004_out1 <= Logical_Operator_out2980_out1 XOR Logical_Operator_out2984_out1;

  Logical_Operator_out4005_out1 <= Logical_Operator_out1955_out1 XOR Logical_Operator_out1959_out1;

  Logical_Operator_out4006_out1 <= Logical_Operator_out1956_out1 XOR Logical_Operator_out1960_out1;

  Logical_Operator_out4007_out1 <= Logical_Operator_out932_out1 XOR Logical_Operator_out936_out1;

  Logical_Operator_out4008_out1 <= in1864 XOR in1872;

  Logical_Operator_out4009_out1 <= Logical_Operator_out2985_out1 XOR Logical_Operator_out2989_out1;

  Logical_Operator_out4010_out1 <= Logical_Operator_out2986_out1 XOR Logical_Operator_out2990_out1;

  Logical_Operator_out4011_out1 <= Logical_Operator_out2987_out1 XOR Logical_Operator_out2991_out1;

  Logical_Operator_out4012_out1 <= Logical_Operator_out2988_out1 XOR Logical_Operator_out2992_out1;

  Logical_Operator_out4013_out1 <= Logical_Operator_out1963_out1 XOR Logical_Operator_out1967_out1;

  Logical_Operator_out4014_out1 <= Logical_Operator_out1964_out1 XOR Logical_Operator_out1968_out1;

  Logical_Operator_out4015_out1 <= Logical_Operator_out940_out1 XOR Logical_Operator_out944_out1;

  Logical_Operator_out4016_out1 <= in1880 XOR in1888;

  Logical_Operator_out4017_out1 <= Logical_Operator_out2993_out1 XOR Logical_Operator_out2997_out1;

  Logical_Operator_out4018_out1 <= Logical_Operator_out2994_out1 XOR Logical_Operator_out2998_out1;

  Logical_Operator_out4019_out1 <= Logical_Operator_out2995_out1 XOR Logical_Operator_out2999_out1;

  Logical_Operator_out4020_out1 <= Logical_Operator_out2996_out1 XOR Logical_Operator_out3000_out1;

  Logical_Operator_out4021_out1 <= Logical_Operator_out1971_out1 XOR Logical_Operator_out1975_out1;

  Logical_Operator_out4022_out1 <= Logical_Operator_out1972_out1 XOR Logical_Operator_out1976_out1;

  Logical_Operator_out4023_out1 <= Logical_Operator_out948_out1 XOR Logical_Operator_out952_out1;

  Logical_Operator_out4024_out1 <= in1896 XOR in1904;

  Logical_Operator_out4025_out1 <= Logical_Operator_out3001_out1 XOR Logical_Operator_out3005_out1;

  Logical_Operator_out4026_out1 <= Logical_Operator_out3002_out1 XOR Logical_Operator_out3006_out1;

  Logical_Operator_out4027_out1 <= Logical_Operator_out3003_out1 XOR Logical_Operator_out3007_out1;

  Logical_Operator_out4028_out1 <= Logical_Operator_out3004_out1 XOR Logical_Operator_out3008_out1;

  Logical_Operator_out4029_out1 <= Logical_Operator_out1979_out1 XOR Logical_Operator_out1983_out1;

  Logical_Operator_out4030_out1 <= Logical_Operator_out1980_out1 XOR Logical_Operator_out1984_out1;

  Logical_Operator_out4031_out1 <= Logical_Operator_out956_out1 XOR Logical_Operator_out960_out1;

  Logical_Operator_out4032_out1 <= in1912 XOR in1920;

  Logical_Operator_out4033_out1 <= Logical_Operator_out3009_out1 XOR Logical_Operator_out3013_out1;

  Logical_Operator_out4034_out1 <= Logical_Operator_out3010_out1 XOR Logical_Operator_out3014_out1;

  Logical_Operator_out4035_out1 <= Logical_Operator_out3011_out1 XOR Logical_Operator_out3015_out1;

  Logical_Operator_out4036_out1 <= Logical_Operator_out3012_out1 XOR Logical_Operator_out3016_out1;

  Logical_Operator_out4037_out1 <= Logical_Operator_out1987_out1 XOR Logical_Operator_out1991_out1;

  Logical_Operator_out4038_out1 <= Logical_Operator_out1988_out1 XOR Logical_Operator_out1992_out1;

  Logical_Operator_out4039_out1 <= Logical_Operator_out964_out1 XOR Logical_Operator_out968_out1;

  Logical_Operator_out4040_out1 <= in1928 XOR in1936;

  Logical_Operator_out4041_out1 <= Logical_Operator_out3017_out1 XOR Logical_Operator_out3021_out1;

  Logical_Operator_out4042_out1 <= Logical_Operator_out3018_out1 XOR Logical_Operator_out3022_out1;

  Logical_Operator_out4043_out1 <= Logical_Operator_out3019_out1 XOR Logical_Operator_out3023_out1;

  Logical_Operator_out4044_out1 <= Logical_Operator_out3020_out1 XOR Logical_Operator_out3024_out1;

  Logical_Operator_out4045_out1 <= Logical_Operator_out1995_out1 XOR Logical_Operator_out1999_out1;

  Logical_Operator_out4046_out1 <= Logical_Operator_out1996_out1 XOR Logical_Operator_out2000_out1;

  Logical_Operator_out4047_out1 <= Logical_Operator_out972_out1 XOR Logical_Operator_out976_out1;

  Logical_Operator_out4048_out1 <= in1944 XOR in1952;

  Logical_Operator_out4049_out1 <= Logical_Operator_out3025_out1 XOR Logical_Operator_out3029_out1;

  Logical_Operator_out4050_out1 <= Logical_Operator_out3026_out1 XOR Logical_Operator_out3030_out1;

  Logical_Operator_out4051_out1 <= Logical_Operator_out3027_out1 XOR Logical_Operator_out3031_out1;

  Logical_Operator_out4052_out1 <= Logical_Operator_out3028_out1 XOR Logical_Operator_out3032_out1;

  Logical_Operator_out4053_out1 <= Logical_Operator_out2003_out1 XOR Logical_Operator_out2007_out1;

  Logical_Operator_out4054_out1 <= Logical_Operator_out2004_out1 XOR Logical_Operator_out2008_out1;

  Logical_Operator_out4055_out1 <= Logical_Operator_out980_out1 XOR Logical_Operator_out984_out1;

  Logical_Operator_out4056_out1 <= in1960 XOR in1968;

  Logical_Operator_out4057_out1 <= Logical_Operator_out3033_out1 XOR Logical_Operator_out3037_out1;

  Logical_Operator_out4058_out1 <= Logical_Operator_out3034_out1 XOR Logical_Operator_out3038_out1;

  Logical_Operator_out4059_out1 <= Logical_Operator_out3035_out1 XOR Logical_Operator_out3039_out1;

  Logical_Operator_out4060_out1 <= Logical_Operator_out3036_out1 XOR Logical_Operator_out3040_out1;

  Logical_Operator_out4061_out1 <= Logical_Operator_out2011_out1 XOR Logical_Operator_out2015_out1;

  Logical_Operator_out4062_out1 <= Logical_Operator_out2012_out1 XOR Logical_Operator_out2016_out1;

  Logical_Operator_out4063_out1 <= Logical_Operator_out988_out1 XOR Logical_Operator_out992_out1;

  Logical_Operator_out4064_out1 <= in1976 XOR in1984;

  Logical_Operator_out4065_out1 <= Logical_Operator_out3041_out1 XOR Logical_Operator_out3045_out1;

  Logical_Operator_out4066_out1 <= Logical_Operator_out3042_out1 XOR Logical_Operator_out3046_out1;

  Logical_Operator_out4067_out1 <= Logical_Operator_out3043_out1 XOR Logical_Operator_out3047_out1;

  Logical_Operator_out4068_out1 <= Logical_Operator_out3044_out1 XOR Logical_Operator_out3048_out1;

  Logical_Operator_out4069_out1 <= Logical_Operator_out2019_out1 XOR Logical_Operator_out2023_out1;

  Logical_Operator_out4070_out1 <= Logical_Operator_out2020_out1 XOR Logical_Operator_out2024_out1;

  Logical_Operator_out4071_out1 <= Logical_Operator_out996_out1 XOR Logical_Operator_out1000_out1;

  Logical_Operator_out4072_out1 <= in1992 XOR in2000;

  Logical_Operator_out4073_out1 <= Logical_Operator_out3049_out1 XOR Logical_Operator_out3053_out1;

  Logical_Operator_out4074_out1 <= Logical_Operator_out3050_out1 XOR Logical_Operator_out3054_out1;

  Logical_Operator_out4075_out1 <= Logical_Operator_out3051_out1 XOR Logical_Operator_out3055_out1;

  Logical_Operator_out4076_out1 <= Logical_Operator_out3052_out1 XOR Logical_Operator_out3056_out1;

  Logical_Operator_out4077_out1 <= Logical_Operator_out2027_out1 XOR Logical_Operator_out2031_out1;

  Logical_Operator_out4078_out1 <= Logical_Operator_out2028_out1 XOR Logical_Operator_out2032_out1;

  Logical_Operator_out4079_out1 <= Logical_Operator_out1004_out1 XOR Logical_Operator_out1008_out1;

  Logical_Operator_out4080_out1 <= in2008 XOR in2016;

  Logical_Operator_out4081_out1 <= Logical_Operator_out3057_out1 XOR Logical_Operator_out3061_out1;

  Logical_Operator_out4082_out1 <= Logical_Operator_out3058_out1 XOR Logical_Operator_out3062_out1;

  Logical_Operator_out4083_out1 <= Logical_Operator_out3059_out1 XOR Logical_Operator_out3063_out1;

  Logical_Operator_out4084_out1 <= Logical_Operator_out3060_out1 XOR Logical_Operator_out3064_out1;

  Logical_Operator_out4085_out1 <= Logical_Operator_out2035_out1 XOR Logical_Operator_out2039_out1;

  Logical_Operator_out4086_out1 <= Logical_Operator_out2036_out1 XOR Logical_Operator_out2040_out1;

  Logical_Operator_out4087_out1 <= Logical_Operator_out1012_out1 XOR Logical_Operator_out1016_out1;

  Logical_Operator_out4088_out1 <= in2024 XOR in2032;

  Logical_Operator_out4089_out1 <= Logical_Operator_out3065_out1 XOR Logical_Operator_out3069_out1;

  Logical_Operator_out4090_out1 <= Logical_Operator_out3066_out1 XOR Logical_Operator_out3070_out1;

  Logical_Operator_out4091_out1 <= Logical_Operator_out3067_out1 XOR Logical_Operator_out3071_out1;

  Logical_Operator_out4092_out1 <= Logical_Operator_out3068_out1 XOR Logical_Operator_out3072_out1;

  Logical_Operator_out4093_out1 <= Logical_Operator_out2043_out1 XOR Logical_Operator_out2047_out1;

  Logical_Operator_out4094_out1 <= Logical_Operator_out2044_out1 XOR Logical_Operator_out2048_out1;

  Logical_Operator_out4095_out1 <= Logical_Operator_out1020_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out4096_out1 <= in2040 XOR in2048;

  Logical_Operator_out4097_out1 <= Logical_Operator_out3073_out1 XOR Logical_Operator_out3081_out1;

  Logical_Operator_out4098_out1 <= Logical_Operator_out3074_out1 XOR Logical_Operator_out3082_out1;

  Logical_Operator_out4099_out1 <= Logical_Operator_out3075_out1 XOR Logical_Operator_out3083_out1;

  Logical_Operator_out4100_out1 <= Logical_Operator_out3076_out1 XOR Logical_Operator_out3084_out1;

  Logical_Operator_out4101_out1 <= Logical_Operator_out3077_out1 XOR Logical_Operator_out3085_out1;

  Logical_Operator_out4102_out1 <= Logical_Operator_out3078_out1 XOR Logical_Operator_out3086_out1;

  Logical_Operator_out4103_out1 <= Logical_Operator_out3079_out1 XOR Logical_Operator_out3087_out1;

  Logical_Operator_out4104_out1 <= Logical_Operator_out3080_out1 XOR Logical_Operator_out3088_out1;

  Logical_Operator_out4105_out1 <= Logical_Operator_out2053_out1 XOR Logical_Operator_out2061_out1;

  Logical_Operator_out4106_out1 <= Logical_Operator_out2054_out1 XOR Logical_Operator_out2062_out1;

  Logical_Operator_out4107_out1 <= Logical_Operator_out2055_out1 XOR Logical_Operator_out2063_out1;

  Logical_Operator_out4108_out1 <= Logical_Operator_out2056_out1 XOR Logical_Operator_out2064_out1;

  Logical_Operator_out4109_out1 <= Logical_Operator_out1031_out1 XOR Logical_Operator_out1039_out1;

  Logical_Operator_out4110_out1 <= Logical_Operator_out1032_out1 XOR Logical_Operator_out1040_out1;

  Logical_Operator_out4111_out1 <= Logical_Operator_out8_out1 XOR Logical_Operator_out16_out1;

  Logical_Operator_out4112_out1 <= in16 XOR in32;

  Logical_Operator_out4113_out1 <= Logical_Operator_out3089_out1 XOR Logical_Operator_out3097_out1;

  Logical_Operator_out4114_out1 <= Logical_Operator_out3090_out1 XOR Logical_Operator_out3098_out1;

  Logical_Operator_out4115_out1 <= Logical_Operator_out3091_out1 XOR Logical_Operator_out3099_out1;

  Logical_Operator_out4116_out1 <= Logical_Operator_out3092_out1 XOR Logical_Operator_out3100_out1;

  Logical_Operator_out4117_out1 <= Logical_Operator_out3093_out1 XOR Logical_Operator_out3101_out1;

  Logical_Operator_out4118_out1 <= Logical_Operator_out3094_out1 XOR Logical_Operator_out3102_out1;

  Logical_Operator_out4119_out1 <= Logical_Operator_out3095_out1 XOR Logical_Operator_out3103_out1;

  Logical_Operator_out4120_out1 <= Logical_Operator_out3096_out1 XOR Logical_Operator_out3104_out1;

  Logical_Operator_out4121_out1 <= Logical_Operator_out2069_out1 XOR Logical_Operator_out2077_out1;

  Logical_Operator_out4122_out1 <= Logical_Operator_out2070_out1 XOR Logical_Operator_out2078_out1;

  Logical_Operator_out4123_out1 <= Logical_Operator_out2071_out1 XOR Logical_Operator_out2079_out1;

  Logical_Operator_out4124_out1 <= Logical_Operator_out2072_out1 XOR Logical_Operator_out2080_out1;

  Logical_Operator_out4125_out1 <= Logical_Operator_out1047_out1 XOR Logical_Operator_out1055_out1;

  Logical_Operator_out4126_out1 <= Logical_Operator_out1048_out1 XOR Logical_Operator_out1056_out1;

  Logical_Operator_out4127_out1 <= Logical_Operator_out24_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out4128_out1 <= in48 XOR in64;

  Logical_Operator_out4129_out1 <= Logical_Operator_out3105_out1 XOR Logical_Operator_out3113_out1;

  Logical_Operator_out4130_out1 <= Logical_Operator_out3106_out1 XOR Logical_Operator_out3114_out1;

  Logical_Operator_out4131_out1 <= Logical_Operator_out3107_out1 XOR Logical_Operator_out3115_out1;

  Logical_Operator_out4132_out1 <= Logical_Operator_out3108_out1 XOR Logical_Operator_out3116_out1;

  Logical_Operator_out4133_out1 <= Logical_Operator_out3109_out1 XOR Logical_Operator_out3117_out1;

  Logical_Operator_out4134_out1 <= Logical_Operator_out3110_out1 XOR Logical_Operator_out3118_out1;

  Logical_Operator_out4135_out1 <= Logical_Operator_out3111_out1 XOR Logical_Operator_out3119_out1;

  Logical_Operator_out4136_out1 <= Logical_Operator_out3112_out1 XOR Logical_Operator_out3120_out1;

  Logical_Operator_out4137_out1 <= Logical_Operator_out2085_out1 XOR Logical_Operator_out2093_out1;

  Logical_Operator_out4138_out1 <= Logical_Operator_out2086_out1 XOR Logical_Operator_out2094_out1;

  Logical_Operator_out4139_out1 <= Logical_Operator_out2087_out1 XOR Logical_Operator_out2095_out1;

  Logical_Operator_out4140_out1 <= Logical_Operator_out2088_out1 XOR Logical_Operator_out2096_out1;

  Logical_Operator_out4141_out1 <= Logical_Operator_out1063_out1 XOR Logical_Operator_out1071_out1;

  Logical_Operator_out4142_out1 <= Logical_Operator_out1064_out1 XOR Logical_Operator_out1072_out1;

  Logical_Operator_out4143_out1 <= Logical_Operator_out40_out1 XOR Logical_Operator_out48_out1;

  Logical_Operator_out4144_out1 <= in80 XOR in96;

  Logical_Operator_out4145_out1 <= Logical_Operator_out3121_out1 XOR Logical_Operator_out3129_out1;

  Logical_Operator_out4146_out1 <= Logical_Operator_out3122_out1 XOR Logical_Operator_out3130_out1;

  Logical_Operator_out4147_out1 <= Logical_Operator_out3123_out1 XOR Logical_Operator_out3131_out1;

  Logical_Operator_out4148_out1 <= Logical_Operator_out3124_out1 XOR Logical_Operator_out3132_out1;

  Logical_Operator_out4149_out1 <= Logical_Operator_out3125_out1 XOR Logical_Operator_out3133_out1;

  Logical_Operator_out4150_out1 <= Logical_Operator_out3126_out1 XOR Logical_Operator_out3134_out1;

  Logical_Operator_out4151_out1 <= Logical_Operator_out3127_out1 XOR Logical_Operator_out3135_out1;

  Logical_Operator_out4152_out1 <= Logical_Operator_out3128_out1 XOR Logical_Operator_out3136_out1;

  Logical_Operator_out4153_out1 <= Logical_Operator_out2101_out1 XOR Logical_Operator_out2109_out1;

  Logical_Operator_out4154_out1 <= Logical_Operator_out2102_out1 XOR Logical_Operator_out2110_out1;

  Logical_Operator_out4155_out1 <= Logical_Operator_out2103_out1 XOR Logical_Operator_out2111_out1;

  Logical_Operator_out4156_out1 <= Logical_Operator_out2104_out1 XOR Logical_Operator_out2112_out1;

  Logical_Operator_out4157_out1 <= Logical_Operator_out1079_out1 XOR Logical_Operator_out1087_out1;

  Logical_Operator_out4158_out1 <= Logical_Operator_out1080_out1 XOR Logical_Operator_out1088_out1;

  Logical_Operator_out4159_out1 <= Logical_Operator_out56_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out4160_out1 <= in112 XOR in128;

  Logical_Operator_out4161_out1 <= Logical_Operator_out3137_out1 XOR Logical_Operator_out3145_out1;

  Logical_Operator_out4162_out1 <= Logical_Operator_out3138_out1 XOR Logical_Operator_out3146_out1;

  Logical_Operator_out4163_out1 <= Logical_Operator_out3139_out1 XOR Logical_Operator_out3147_out1;

  Logical_Operator_out4164_out1 <= Logical_Operator_out3140_out1 XOR Logical_Operator_out3148_out1;

  Logical_Operator_out4165_out1 <= Logical_Operator_out3141_out1 XOR Logical_Operator_out3149_out1;

  Logical_Operator_out4166_out1 <= Logical_Operator_out3142_out1 XOR Logical_Operator_out3150_out1;

  Logical_Operator_out4167_out1 <= Logical_Operator_out3143_out1 XOR Logical_Operator_out3151_out1;

  Logical_Operator_out4168_out1 <= Logical_Operator_out3144_out1 XOR Logical_Operator_out3152_out1;

  Logical_Operator_out4169_out1 <= Logical_Operator_out2117_out1 XOR Logical_Operator_out2125_out1;

  Logical_Operator_out4170_out1 <= Logical_Operator_out2118_out1 XOR Logical_Operator_out2126_out1;

  Logical_Operator_out4171_out1 <= Logical_Operator_out2119_out1 XOR Logical_Operator_out2127_out1;

  Logical_Operator_out4172_out1 <= Logical_Operator_out2120_out1 XOR Logical_Operator_out2128_out1;

  Logical_Operator_out4173_out1 <= Logical_Operator_out1095_out1 XOR Logical_Operator_out1103_out1;

  Logical_Operator_out4174_out1 <= Logical_Operator_out1096_out1 XOR Logical_Operator_out1104_out1;

  Logical_Operator_out4175_out1 <= Logical_Operator_out72_out1 XOR Logical_Operator_out80_out1;

  Logical_Operator_out4176_out1 <= in144 XOR in160;

  Logical_Operator_out4177_out1 <= Logical_Operator_out3153_out1 XOR Logical_Operator_out3161_out1;

  Logical_Operator_out4178_out1 <= Logical_Operator_out3154_out1 XOR Logical_Operator_out3162_out1;

  Logical_Operator_out4179_out1 <= Logical_Operator_out3155_out1 XOR Logical_Operator_out3163_out1;

  Logical_Operator_out4180_out1 <= Logical_Operator_out3156_out1 XOR Logical_Operator_out3164_out1;

  Logical_Operator_out4181_out1 <= Logical_Operator_out3157_out1 XOR Logical_Operator_out3165_out1;

  Logical_Operator_out4182_out1 <= Logical_Operator_out3158_out1 XOR Logical_Operator_out3166_out1;

  Logical_Operator_out4183_out1 <= Logical_Operator_out3159_out1 XOR Logical_Operator_out3167_out1;

  Logical_Operator_out4184_out1 <= Logical_Operator_out3160_out1 XOR Logical_Operator_out3168_out1;

  Logical_Operator_out4185_out1 <= Logical_Operator_out2133_out1 XOR Logical_Operator_out2141_out1;

  Logical_Operator_out4186_out1 <= Logical_Operator_out2134_out1 XOR Logical_Operator_out2142_out1;

  Logical_Operator_out4187_out1 <= Logical_Operator_out2135_out1 XOR Logical_Operator_out2143_out1;

  Logical_Operator_out4188_out1 <= Logical_Operator_out2136_out1 XOR Logical_Operator_out2144_out1;

  Logical_Operator_out4189_out1 <= Logical_Operator_out1111_out1 XOR Logical_Operator_out1119_out1;

  Logical_Operator_out4190_out1 <= Logical_Operator_out1112_out1 XOR Logical_Operator_out1120_out1;

  Logical_Operator_out4191_out1 <= Logical_Operator_out88_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out4192_out1 <= in176 XOR in192;

  Logical_Operator_out4193_out1 <= Logical_Operator_out3169_out1 XOR Logical_Operator_out3177_out1;

  Logical_Operator_out4194_out1 <= Logical_Operator_out3170_out1 XOR Logical_Operator_out3178_out1;

  Logical_Operator_out4195_out1 <= Logical_Operator_out3171_out1 XOR Logical_Operator_out3179_out1;

  Logical_Operator_out4196_out1 <= Logical_Operator_out3172_out1 XOR Logical_Operator_out3180_out1;

  Logical_Operator_out4197_out1 <= Logical_Operator_out3173_out1 XOR Logical_Operator_out3181_out1;

  Logical_Operator_out4198_out1 <= Logical_Operator_out3174_out1 XOR Logical_Operator_out3182_out1;

  Logical_Operator_out4199_out1 <= Logical_Operator_out3175_out1 XOR Logical_Operator_out3183_out1;

  Logical_Operator_out4200_out1 <= Logical_Operator_out3176_out1 XOR Logical_Operator_out3184_out1;

  Logical_Operator_out4201_out1 <= Logical_Operator_out2149_out1 XOR Logical_Operator_out2157_out1;

  Logical_Operator_out4202_out1 <= Logical_Operator_out2150_out1 XOR Logical_Operator_out2158_out1;

  Logical_Operator_out4203_out1 <= Logical_Operator_out2151_out1 XOR Logical_Operator_out2159_out1;

  Logical_Operator_out4204_out1 <= Logical_Operator_out2152_out1 XOR Logical_Operator_out2160_out1;

  Logical_Operator_out4205_out1 <= Logical_Operator_out1127_out1 XOR Logical_Operator_out1135_out1;

  Logical_Operator_out4206_out1 <= Logical_Operator_out1128_out1 XOR Logical_Operator_out1136_out1;

  Logical_Operator_out4207_out1 <= Logical_Operator_out104_out1 XOR Logical_Operator_out112_out1;

  Logical_Operator_out4208_out1 <= in208 XOR in224;

  Logical_Operator_out4209_out1 <= Logical_Operator_out3185_out1 XOR Logical_Operator_out3193_out1;

  Logical_Operator_out4210_out1 <= Logical_Operator_out3186_out1 XOR Logical_Operator_out3194_out1;

  Logical_Operator_out4211_out1 <= Logical_Operator_out3187_out1 XOR Logical_Operator_out3195_out1;

  Logical_Operator_out4212_out1 <= Logical_Operator_out3188_out1 XOR Logical_Operator_out3196_out1;

  Logical_Operator_out4213_out1 <= Logical_Operator_out3189_out1 XOR Logical_Operator_out3197_out1;

  Logical_Operator_out4214_out1 <= Logical_Operator_out3190_out1 XOR Logical_Operator_out3198_out1;

  Logical_Operator_out4215_out1 <= Logical_Operator_out3191_out1 XOR Logical_Operator_out3199_out1;

  Logical_Operator_out4216_out1 <= Logical_Operator_out3192_out1 XOR Logical_Operator_out3200_out1;

  Logical_Operator_out4217_out1 <= Logical_Operator_out2165_out1 XOR Logical_Operator_out2173_out1;

  Logical_Operator_out4218_out1 <= Logical_Operator_out2166_out1 XOR Logical_Operator_out2174_out1;

  Logical_Operator_out4219_out1 <= Logical_Operator_out2167_out1 XOR Logical_Operator_out2175_out1;

  Logical_Operator_out4220_out1 <= Logical_Operator_out2168_out1 XOR Logical_Operator_out2176_out1;

  Logical_Operator_out4221_out1 <= Logical_Operator_out1143_out1 XOR Logical_Operator_out1151_out1;

  Logical_Operator_out4222_out1 <= Logical_Operator_out1144_out1 XOR Logical_Operator_out1152_out1;

  Logical_Operator_out4223_out1 <= Logical_Operator_out120_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out4224_out1 <= in240 XOR in256;

  Logical_Operator_out4225_out1 <= Logical_Operator_out3201_out1 XOR Logical_Operator_out3209_out1;

  Logical_Operator_out4226_out1 <= Logical_Operator_out3202_out1 XOR Logical_Operator_out3210_out1;

  Logical_Operator_out4227_out1 <= Logical_Operator_out3203_out1 XOR Logical_Operator_out3211_out1;

  Logical_Operator_out4228_out1 <= Logical_Operator_out3204_out1 XOR Logical_Operator_out3212_out1;

  Logical_Operator_out4229_out1 <= Logical_Operator_out3205_out1 XOR Logical_Operator_out3213_out1;

  Logical_Operator_out4230_out1 <= Logical_Operator_out3206_out1 XOR Logical_Operator_out3214_out1;

  Logical_Operator_out4231_out1 <= Logical_Operator_out3207_out1 XOR Logical_Operator_out3215_out1;

  Logical_Operator_out4232_out1 <= Logical_Operator_out3208_out1 XOR Logical_Operator_out3216_out1;

  Logical_Operator_out4233_out1 <= Logical_Operator_out2181_out1 XOR Logical_Operator_out2189_out1;

  Logical_Operator_out4234_out1 <= Logical_Operator_out2182_out1 XOR Logical_Operator_out2190_out1;

  Logical_Operator_out4235_out1 <= Logical_Operator_out2183_out1 XOR Logical_Operator_out2191_out1;

  Logical_Operator_out4236_out1 <= Logical_Operator_out2184_out1 XOR Logical_Operator_out2192_out1;

  Logical_Operator_out4237_out1 <= Logical_Operator_out1159_out1 XOR Logical_Operator_out1167_out1;

  Logical_Operator_out4238_out1 <= Logical_Operator_out1160_out1 XOR Logical_Operator_out1168_out1;

  Logical_Operator_out4239_out1 <= Logical_Operator_out136_out1 XOR Logical_Operator_out144_out1;

  Logical_Operator_out4240_out1 <= in272 XOR in288;

  Logical_Operator_out4241_out1 <= Logical_Operator_out3217_out1 XOR Logical_Operator_out3225_out1;

  Logical_Operator_out4242_out1 <= Logical_Operator_out3218_out1 XOR Logical_Operator_out3226_out1;

  Logical_Operator_out4243_out1 <= Logical_Operator_out3219_out1 XOR Logical_Operator_out3227_out1;

  Logical_Operator_out4244_out1 <= Logical_Operator_out3220_out1 XOR Logical_Operator_out3228_out1;

  Logical_Operator_out4245_out1 <= Logical_Operator_out3221_out1 XOR Logical_Operator_out3229_out1;

  Logical_Operator_out4246_out1 <= Logical_Operator_out3222_out1 XOR Logical_Operator_out3230_out1;

  Logical_Operator_out4247_out1 <= Logical_Operator_out3223_out1 XOR Logical_Operator_out3231_out1;

  Logical_Operator_out4248_out1 <= Logical_Operator_out3224_out1 XOR Logical_Operator_out3232_out1;

  Logical_Operator_out4249_out1 <= Logical_Operator_out2197_out1 XOR Logical_Operator_out2205_out1;

  Logical_Operator_out4250_out1 <= Logical_Operator_out2198_out1 XOR Logical_Operator_out2206_out1;

  Logical_Operator_out4251_out1 <= Logical_Operator_out2199_out1 XOR Logical_Operator_out2207_out1;

  Logical_Operator_out4252_out1 <= Logical_Operator_out2200_out1 XOR Logical_Operator_out2208_out1;

  Logical_Operator_out4253_out1 <= Logical_Operator_out1175_out1 XOR Logical_Operator_out1183_out1;

  Logical_Operator_out4254_out1 <= Logical_Operator_out1176_out1 XOR Logical_Operator_out1184_out1;

  Logical_Operator_out4255_out1 <= Logical_Operator_out152_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out4256_out1 <= in304 XOR in320;

  Logical_Operator_out4257_out1 <= Logical_Operator_out3233_out1 XOR Logical_Operator_out3241_out1;

  Logical_Operator_out4258_out1 <= Logical_Operator_out3234_out1 XOR Logical_Operator_out3242_out1;

  Logical_Operator_out4259_out1 <= Logical_Operator_out3235_out1 XOR Logical_Operator_out3243_out1;

  Logical_Operator_out4260_out1 <= Logical_Operator_out3236_out1 XOR Logical_Operator_out3244_out1;

  Logical_Operator_out4261_out1 <= Logical_Operator_out3237_out1 XOR Logical_Operator_out3245_out1;

  Logical_Operator_out4262_out1 <= Logical_Operator_out3238_out1 XOR Logical_Operator_out3246_out1;

  Logical_Operator_out4263_out1 <= Logical_Operator_out3239_out1 XOR Logical_Operator_out3247_out1;

  Logical_Operator_out4264_out1 <= Logical_Operator_out3240_out1 XOR Logical_Operator_out3248_out1;

  Logical_Operator_out4265_out1 <= Logical_Operator_out2213_out1 XOR Logical_Operator_out2221_out1;

  Logical_Operator_out4266_out1 <= Logical_Operator_out2214_out1 XOR Logical_Operator_out2222_out1;

  Logical_Operator_out4267_out1 <= Logical_Operator_out2215_out1 XOR Logical_Operator_out2223_out1;

  Logical_Operator_out4268_out1 <= Logical_Operator_out2216_out1 XOR Logical_Operator_out2224_out1;

  Logical_Operator_out4269_out1 <= Logical_Operator_out1191_out1 XOR Logical_Operator_out1199_out1;

  Logical_Operator_out4270_out1 <= Logical_Operator_out1192_out1 XOR Logical_Operator_out1200_out1;

  Logical_Operator_out4271_out1 <= Logical_Operator_out168_out1 XOR Logical_Operator_out176_out1;

  Logical_Operator_out4272_out1 <= in336 XOR in352;

  Logical_Operator_out4273_out1 <= Logical_Operator_out3249_out1 XOR Logical_Operator_out3257_out1;

  Logical_Operator_out4274_out1 <= Logical_Operator_out3250_out1 XOR Logical_Operator_out3258_out1;

  Logical_Operator_out4275_out1 <= Logical_Operator_out3251_out1 XOR Logical_Operator_out3259_out1;

  Logical_Operator_out4276_out1 <= Logical_Operator_out3252_out1 XOR Logical_Operator_out3260_out1;

  Logical_Operator_out4277_out1 <= Logical_Operator_out3253_out1 XOR Logical_Operator_out3261_out1;

  Logical_Operator_out4278_out1 <= Logical_Operator_out3254_out1 XOR Logical_Operator_out3262_out1;

  Logical_Operator_out4279_out1 <= Logical_Operator_out3255_out1 XOR Logical_Operator_out3263_out1;

  Logical_Operator_out4280_out1 <= Logical_Operator_out3256_out1 XOR Logical_Operator_out3264_out1;

  Logical_Operator_out4281_out1 <= Logical_Operator_out2229_out1 XOR Logical_Operator_out2237_out1;

  Logical_Operator_out4282_out1 <= Logical_Operator_out2230_out1 XOR Logical_Operator_out2238_out1;

  Logical_Operator_out4283_out1 <= Logical_Operator_out2231_out1 XOR Logical_Operator_out2239_out1;

  Logical_Operator_out4284_out1 <= Logical_Operator_out2232_out1 XOR Logical_Operator_out2240_out1;

  Logical_Operator_out4285_out1 <= Logical_Operator_out1207_out1 XOR Logical_Operator_out1215_out1;

  Logical_Operator_out4286_out1 <= Logical_Operator_out1208_out1 XOR Logical_Operator_out1216_out1;

  Logical_Operator_out4287_out1 <= Logical_Operator_out184_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out4288_out1 <= in368 XOR in384;

  Logical_Operator_out4289_out1 <= Logical_Operator_out3265_out1 XOR Logical_Operator_out3273_out1;

  Logical_Operator_out4290_out1 <= Logical_Operator_out3266_out1 XOR Logical_Operator_out3274_out1;

  Logical_Operator_out4291_out1 <= Logical_Operator_out3267_out1 XOR Logical_Operator_out3275_out1;

  Logical_Operator_out4292_out1 <= Logical_Operator_out3268_out1 XOR Logical_Operator_out3276_out1;

  Logical_Operator_out4293_out1 <= Logical_Operator_out3269_out1 XOR Logical_Operator_out3277_out1;

  Logical_Operator_out4294_out1 <= Logical_Operator_out3270_out1 XOR Logical_Operator_out3278_out1;

  Logical_Operator_out4295_out1 <= Logical_Operator_out3271_out1 XOR Logical_Operator_out3279_out1;

  Logical_Operator_out4296_out1 <= Logical_Operator_out3272_out1 XOR Logical_Operator_out3280_out1;

  Logical_Operator_out4297_out1 <= Logical_Operator_out2245_out1 XOR Logical_Operator_out2253_out1;

  Logical_Operator_out4298_out1 <= Logical_Operator_out2246_out1 XOR Logical_Operator_out2254_out1;

  Logical_Operator_out4299_out1 <= Logical_Operator_out2247_out1 XOR Logical_Operator_out2255_out1;

  Logical_Operator_out4300_out1 <= Logical_Operator_out2248_out1 XOR Logical_Operator_out2256_out1;

  Logical_Operator_out4301_out1 <= Logical_Operator_out1223_out1 XOR Logical_Operator_out1231_out1;

  Logical_Operator_out4302_out1 <= Logical_Operator_out1224_out1 XOR Logical_Operator_out1232_out1;

  Logical_Operator_out4303_out1 <= Logical_Operator_out200_out1 XOR Logical_Operator_out208_out1;

  Logical_Operator_out4304_out1 <= in400 XOR in416;

  Logical_Operator_out4305_out1 <= Logical_Operator_out3281_out1 XOR Logical_Operator_out3289_out1;

  Logical_Operator_out4306_out1 <= Logical_Operator_out3282_out1 XOR Logical_Operator_out3290_out1;

  Logical_Operator_out4307_out1 <= Logical_Operator_out3283_out1 XOR Logical_Operator_out3291_out1;

  Logical_Operator_out4308_out1 <= Logical_Operator_out3284_out1 XOR Logical_Operator_out3292_out1;

  Logical_Operator_out4309_out1 <= Logical_Operator_out3285_out1 XOR Logical_Operator_out3293_out1;

  Logical_Operator_out4310_out1 <= Logical_Operator_out3286_out1 XOR Logical_Operator_out3294_out1;

  Logical_Operator_out4311_out1 <= Logical_Operator_out3287_out1 XOR Logical_Operator_out3295_out1;

  Logical_Operator_out4312_out1 <= Logical_Operator_out3288_out1 XOR Logical_Operator_out3296_out1;

  Logical_Operator_out4313_out1 <= Logical_Operator_out2261_out1 XOR Logical_Operator_out2269_out1;

  Logical_Operator_out4314_out1 <= Logical_Operator_out2262_out1 XOR Logical_Operator_out2270_out1;

  Logical_Operator_out4315_out1 <= Logical_Operator_out2263_out1 XOR Logical_Operator_out2271_out1;

  Logical_Operator_out4316_out1 <= Logical_Operator_out2264_out1 XOR Logical_Operator_out2272_out1;

  Logical_Operator_out4317_out1 <= Logical_Operator_out1239_out1 XOR Logical_Operator_out1247_out1;

  Logical_Operator_out4318_out1 <= Logical_Operator_out1240_out1 XOR Logical_Operator_out1248_out1;

  Logical_Operator_out4319_out1 <= Logical_Operator_out216_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out4320_out1 <= in432 XOR in448;

  Logical_Operator_out4321_out1 <= Logical_Operator_out3297_out1 XOR Logical_Operator_out3305_out1;

  Logical_Operator_out4322_out1 <= Logical_Operator_out3298_out1 XOR Logical_Operator_out3306_out1;

  Logical_Operator_out4323_out1 <= Logical_Operator_out3299_out1 XOR Logical_Operator_out3307_out1;

  Logical_Operator_out4324_out1 <= Logical_Operator_out3300_out1 XOR Logical_Operator_out3308_out1;

  Logical_Operator_out4325_out1 <= Logical_Operator_out3301_out1 XOR Logical_Operator_out3309_out1;

  Logical_Operator_out4326_out1 <= Logical_Operator_out3302_out1 XOR Logical_Operator_out3310_out1;

  Logical_Operator_out4327_out1 <= Logical_Operator_out3303_out1 XOR Logical_Operator_out3311_out1;

  Logical_Operator_out4328_out1 <= Logical_Operator_out3304_out1 XOR Logical_Operator_out3312_out1;

  Logical_Operator_out4329_out1 <= Logical_Operator_out2277_out1 XOR Logical_Operator_out2285_out1;

  Logical_Operator_out4330_out1 <= Logical_Operator_out2278_out1 XOR Logical_Operator_out2286_out1;

  Logical_Operator_out4331_out1 <= Logical_Operator_out2279_out1 XOR Logical_Operator_out2287_out1;

  Logical_Operator_out4332_out1 <= Logical_Operator_out2280_out1 XOR Logical_Operator_out2288_out1;

  Logical_Operator_out4333_out1 <= Logical_Operator_out1255_out1 XOR Logical_Operator_out1263_out1;

  Logical_Operator_out4334_out1 <= Logical_Operator_out1256_out1 XOR Logical_Operator_out1264_out1;

  Logical_Operator_out4335_out1 <= Logical_Operator_out232_out1 XOR Logical_Operator_out240_out1;

  Logical_Operator_out4336_out1 <= in464 XOR in480;

  Logical_Operator_out4337_out1 <= Logical_Operator_out3313_out1 XOR Logical_Operator_out3321_out1;

  Logical_Operator_out4338_out1 <= Logical_Operator_out3314_out1 XOR Logical_Operator_out3322_out1;

  Logical_Operator_out4339_out1 <= Logical_Operator_out3315_out1 XOR Logical_Operator_out3323_out1;

  Logical_Operator_out4340_out1 <= Logical_Operator_out3316_out1 XOR Logical_Operator_out3324_out1;

  Logical_Operator_out4341_out1 <= Logical_Operator_out3317_out1 XOR Logical_Operator_out3325_out1;

  Logical_Operator_out4342_out1 <= Logical_Operator_out3318_out1 XOR Logical_Operator_out3326_out1;

  Logical_Operator_out4343_out1 <= Logical_Operator_out3319_out1 XOR Logical_Operator_out3327_out1;

  Logical_Operator_out4344_out1 <= Logical_Operator_out3320_out1 XOR Logical_Operator_out3328_out1;

  Logical_Operator_out4345_out1 <= Logical_Operator_out2293_out1 XOR Logical_Operator_out2301_out1;

  Logical_Operator_out4346_out1 <= Logical_Operator_out2294_out1 XOR Logical_Operator_out2302_out1;

  Logical_Operator_out4347_out1 <= Logical_Operator_out2295_out1 XOR Logical_Operator_out2303_out1;

  Logical_Operator_out4348_out1 <= Logical_Operator_out2296_out1 XOR Logical_Operator_out2304_out1;

  Logical_Operator_out4349_out1 <= Logical_Operator_out1271_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out4350_out1 <= Logical_Operator_out1272_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out4351_out1 <= Logical_Operator_out248_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out4352_out1 <= in496 XOR in512;

  Logical_Operator_out4353_out1 <= Logical_Operator_out3329_out1 XOR Logical_Operator_out3337_out1;

  Logical_Operator_out4354_out1 <= Logical_Operator_out3330_out1 XOR Logical_Operator_out3338_out1;

  Logical_Operator_out4355_out1 <= Logical_Operator_out3331_out1 XOR Logical_Operator_out3339_out1;

  Logical_Operator_out4356_out1 <= Logical_Operator_out3332_out1 XOR Logical_Operator_out3340_out1;

  Logical_Operator_out4357_out1 <= Logical_Operator_out3333_out1 XOR Logical_Operator_out3341_out1;

  Logical_Operator_out4358_out1 <= Logical_Operator_out3334_out1 XOR Logical_Operator_out3342_out1;

  Logical_Operator_out4359_out1 <= Logical_Operator_out3335_out1 XOR Logical_Operator_out3343_out1;

  Logical_Operator_out4360_out1 <= Logical_Operator_out3336_out1 XOR Logical_Operator_out3344_out1;

  Logical_Operator_out4361_out1 <= Logical_Operator_out2309_out1 XOR Logical_Operator_out2317_out1;

  Logical_Operator_out4362_out1 <= Logical_Operator_out2310_out1 XOR Logical_Operator_out2318_out1;

  Logical_Operator_out4363_out1 <= Logical_Operator_out2311_out1 XOR Logical_Operator_out2319_out1;

  Logical_Operator_out4364_out1 <= Logical_Operator_out2312_out1 XOR Logical_Operator_out2320_out1;

  Logical_Operator_out4365_out1 <= Logical_Operator_out1287_out1 XOR Logical_Operator_out1295_out1;

  Logical_Operator_out4366_out1 <= Logical_Operator_out1288_out1 XOR Logical_Operator_out1296_out1;

  Logical_Operator_out4367_out1 <= Logical_Operator_out264_out1 XOR Logical_Operator_out272_out1;

  Logical_Operator_out4368_out1 <= in528 XOR in544;

  Logical_Operator_out4369_out1 <= Logical_Operator_out3345_out1 XOR Logical_Operator_out3353_out1;

  Logical_Operator_out4370_out1 <= Logical_Operator_out3346_out1 XOR Logical_Operator_out3354_out1;

  Logical_Operator_out4371_out1 <= Logical_Operator_out3347_out1 XOR Logical_Operator_out3355_out1;

  Logical_Operator_out4372_out1 <= Logical_Operator_out3348_out1 XOR Logical_Operator_out3356_out1;

  Logical_Operator_out4373_out1 <= Logical_Operator_out3349_out1 XOR Logical_Operator_out3357_out1;

  Logical_Operator_out4374_out1 <= Logical_Operator_out3350_out1 XOR Logical_Operator_out3358_out1;

  Logical_Operator_out4375_out1 <= Logical_Operator_out3351_out1 XOR Logical_Operator_out3359_out1;

  Logical_Operator_out4376_out1 <= Logical_Operator_out3352_out1 XOR Logical_Operator_out3360_out1;

  Logical_Operator_out4377_out1 <= Logical_Operator_out2325_out1 XOR Logical_Operator_out2333_out1;

  Logical_Operator_out4378_out1 <= Logical_Operator_out2326_out1 XOR Logical_Operator_out2334_out1;

  Logical_Operator_out4379_out1 <= Logical_Operator_out2327_out1 XOR Logical_Operator_out2335_out1;

  Logical_Operator_out4380_out1 <= Logical_Operator_out2328_out1 XOR Logical_Operator_out2336_out1;

  Logical_Operator_out4381_out1 <= Logical_Operator_out1303_out1 XOR Logical_Operator_out1311_out1;

  Logical_Operator_out4382_out1 <= Logical_Operator_out1304_out1 XOR Logical_Operator_out1312_out1;

  Logical_Operator_out4383_out1 <= Logical_Operator_out280_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out4384_out1 <= in560 XOR in576;

  Logical_Operator_out4385_out1 <= Logical_Operator_out3361_out1 XOR Logical_Operator_out3369_out1;

  Logical_Operator_out4386_out1 <= Logical_Operator_out3362_out1 XOR Logical_Operator_out3370_out1;

  Logical_Operator_out4387_out1 <= Logical_Operator_out3363_out1 XOR Logical_Operator_out3371_out1;

  Logical_Operator_out4388_out1 <= Logical_Operator_out3364_out1 XOR Logical_Operator_out3372_out1;

  Logical_Operator_out4389_out1 <= Logical_Operator_out3365_out1 XOR Logical_Operator_out3373_out1;

  Logical_Operator_out4390_out1 <= Logical_Operator_out3366_out1 XOR Logical_Operator_out3374_out1;

  Logical_Operator_out4391_out1 <= Logical_Operator_out3367_out1 XOR Logical_Operator_out3375_out1;

  Logical_Operator_out4392_out1 <= Logical_Operator_out3368_out1 XOR Logical_Operator_out3376_out1;

  Logical_Operator_out4393_out1 <= Logical_Operator_out2341_out1 XOR Logical_Operator_out2349_out1;

  Logical_Operator_out4394_out1 <= Logical_Operator_out2342_out1 XOR Logical_Operator_out2350_out1;

  Logical_Operator_out4395_out1 <= Logical_Operator_out2343_out1 XOR Logical_Operator_out2351_out1;

  Logical_Operator_out4396_out1 <= Logical_Operator_out2344_out1 XOR Logical_Operator_out2352_out1;

  Logical_Operator_out4397_out1 <= Logical_Operator_out1319_out1 XOR Logical_Operator_out1327_out1;

  Logical_Operator_out4398_out1 <= Logical_Operator_out1320_out1 XOR Logical_Operator_out1328_out1;

  Logical_Operator_out4399_out1 <= Logical_Operator_out296_out1 XOR Logical_Operator_out304_out1;

  Logical_Operator_out4400_out1 <= in592 XOR in608;

  Logical_Operator_out4401_out1 <= Logical_Operator_out3377_out1 XOR Logical_Operator_out3385_out1;

  Logical_Operator_out4402_out1 <= Logical_Operator_out3378_out1 XOR Logical_Operator_out3386_out1;

  Logical_Operator_out4403_out1 <= Logical_Operator_out3379_out1 XOR Logical_Operator_out3387_out1;

  Logical_Operator_out4404_out1 <= Logical_Operator_out3380_out1 XOR Logical_Operator_out3388_out1;

  Logical_Operator_out4405_out1 <= Logical_Operator_out3381_out1 XOR Logical_Operator_out3389_out1;

  Logical_Operator_out4406_out1 <= Logical_Operator_out3382_out1 XOR Logical_Operator_out3390_out1;

  Logical_Operator_out4407_out1 <= Logical_Operator_out3383_out1 XOR Logical_Operator_out3391_out1;

  Logical_Operator_out4408_out1 <= Logical_Operator_out3384_out1 XOR Logical_Operator_out3392_out1;

  Logical_Operator_out4409_out1 <= Logical_Operator_out2357_out1 XOR Logical_Operator_out2365_out1;

  Logical_Operator_out4410_out1 <= Logical_Operator_out2358_out1 XOR Logical_Operator_out2366_out1;

  Logical_Operator_out4411_out1 <= Logical_Operator_out2359_out1 XOR Logical_Operator_out2367_out1;

  Logical_Operator_out4412_out1 <= Logical_Operator_out2360_out1 XOR Logical_Operator_out2368_out1;

  Logical_Operator_out4413_out1 <= Logical_Operator_out1335_out1 XOR Logical_Operator_out1343_out1;

  Logical_Operator_out4414_out1 <= Logical_Operator_out1336_out1 XOR Logical_Operator_out1344_out1;

  Logical_Operator_out4415_out1 <= Logical_Operator_out312_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out4416_out1 <= in624 XOR in640;

  Logical_Operator_out4417_out1 <= Logical_Operator_out3393_out1 XOR Logical_Operator_out3401_out1;

  Logical_Operator_out4418_out1 <= Logical_Operator_out3394_out1 XOR Logical_Operator_out3402_out1;

  Logical_Operator_out4419_out1 <= Logical_Operator_out3395_out1 XOR Logical_Operator_out3403_out1;

  Logical_Operator_out4420_out1 <= Logical_Operator_out3396_out1 XOR Logical_Operator_out3404_out1;

  Logical_Operator_out4421_out1 <= Logical_Operator_out3397_out1 XOR Logical_Operator_out3405_out1;

  Logical_Operator_out4422_out1 <= Logical_Operator_out3398_out1 XOR Logical_Operator_out3406_out1;

  Logical_Operator_out4423_out1 <= Logical_Operator_out3399_out1 XOR Logical_Operator_out3407_out1;

  Logical_Operator_out4424_out1 <= Logical_Operator_out3400_out1 XOR Logical_Operator_out3408_out1;

  Logical_Operator_out4425_out1 <= Logical_Operator_out2373_out1 XOR Logical_Operator_out2381_out1;

  Logical_Operator_out4426_out1 <= Logical_Operator_out2374_out1 XOR Logical_Operator_out2382_out1;

  Logical_Operator_out4427_out1 <= Logical_Operator_out2375_out1 XOR Logical_Operator_out2383_out1;

  Logical_Operator_out4428_out1 <= Logical_Operator_out2376_out1 XOR Logical_Operator_out2384_out1;

  Logical_Operator_out4429_out1 <= Logical_Operator_out1351_out1 XOR Logical_Operator_out1359_out1;

  Logical_Operator_out4430_out1 <= Logical_Operator_out1352_out1 XOR Logical_Operator_out1360_out1;

  Logical_Operator_out4431_out1 <= Logical_Operator_out328_out1 XOR Logical_Operator_out336_out1;

  Logical_Operator_out4432_out1 <= in656 XOR in672;

  Logical_Operator_out4433_out1 <= Logical_Operator_out3409_out1 XOR Logical_Operator_out3417_out1;

  Logical_Operator_out4434_out1 <= Logical_Operator_out3410_out1 XOR Logical_Operator_out3418_out1;

  Logical_Operator_out4435_out1 <= Logical_Operator_out3411_out1 XOR Logical_Operator_out3419_out1;

  Logical_Operator_out4436_out1 <= Logical_Operator_out3412_out1 XOR Logical_Operator_out3420_out1;

  Logical_Operator_out4437_out1 <= Logical_Operator_out3413_out1 XOR Logical_Operator_out3421_out1;

  Logical_Operator_out4438_out1 <= Logical_Operator_out3414_out1 XOR Logical_Operator_out3422_out1;

  Logical_Operator_out4439_out1 <= Logical_Operator_out3415_out1 XOR Logical_Operator_out3423_out1;

  Logical_Operator_out4440_out1 <= Logical_Operator_out3416_out1 XOR Logical_Operator_out3424_out1;

  Logical_Operator_out4441_out1 <= Logical_Operator_out2389_out1 XOR Logical_Operator_out2397_out1;

  Logical_Operator_out4442_out1 <= Logical_Operator_out2390_out1 XOR Logical_Operator_out2398_out1;

  Logical_Operator_out4443_out1 <= Logical_Operator_out2391_out1 XOR Logical_Operator_out2399_out1;

  Logical_Operator_out4444_out1 <= Logical_Operator_out2392_out1 XOR Logical_Operator_out2400_out1;

  Logical_Operator_out4445_out1 <= Logical_Operator_out1367_out1 XOR Logical_Operator_out1375_out1;

  Logical_Operator_out4446_out1 <= Logical_Operator_out1368_out1 XOR Logical_Operator_out1376_out1;

  Logical_Operator_out4447_out1 <= Logical_Operator_out344_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out4448_out1 <= in688 XOR in704;

  Logical_Operator_out4449_out1 <= Logical_Operator_out3425_out1 XOR Logical_Operator_out3433_out1;

  Logical_Operator_out4450_out1 <= Logical_Operator_out3426_out1 XOR Logical_Operator_out3434_out1;

  Logical_Operator_out4451_out1 <= Logical_Operator_out3427_out1 XOR Logical_Operator_out3435_out1;

  Logical_Operator_out4452_out1 <= Logical_Operator_out3428_out1 XOR Logical_Operator_out3436_out1;

  Logical_Operator_out4453_out1 <= Logical_Operator_out3429_out1 XOR Logical_Operator_out3437_out1;

  Logical_Operator_out4454_out1 <= Logical_Operator_out3430_out1 XOR Logical_Operator_out3438_out1;

  Logical_Operator_out4455_out1 <= Logical_Operator_out3431_out1 XOR Logical_Operator_out3439_out1;

  Logical_Operator_out4456_out1 <= Logical_Operator_out3432_out1 XOR Logical_Operator_out3440_out1;

  Logical_Operator_out4457_out1 <= Logical_Operator_out2405_out1 XOR Logical_Operator_out2413_out1;

  Logical_Operator_out4458_out1 <= Logical_Operator_out2406_out1 XOR Logical_Operator_out2414_out1;

  Logical_Operator_out4459_out1 <= Logical_Operator_out2407_out1 XOR Logical_Operator_out2415_out1;

  Logical_Operator_out4460_out1 <= Logical_Operator_out2408_out1 XOR Logical_Operator_out2416_out1;

  Logical_Operator_out4461_out1 <= Logical_Operator_out1383_out1 XOR Logical_Operator_out1391_out1;

  Logical_Operator_out4462_out1 <= Logical_Operator_out1384_out1 XOR Logical_Operator_out1392_out1;

  Logical_Operator_out4463_out1 <= Logical_Operator_out360_out1 XOR Logical_Operator_out368_out1;

  Logical_Operator_out4464_out1 <= in720 XOR in736;

  Logical_Operator_out4465_out1 <= Logical_Operator_out3441_out1 XOR Logical_Operator_out3449_out1;

  Logical_Operator_out4466_out1 <= Logical_Operator_out3442_out1 XOR Logical_Operator_out3450_out1;

  Logical_Operator_out4467_out1 <= Logical_Operator_out3443_out1 XOR Logical_Operator_out3451_out1;

  Logical_Operator_out4468_out1 <= Logical_Operator_out3444_out1 XOR Logical_Operator_out3452_out1;

  Logical_Operator_out4469_out1 <= Logical_Operator_out3445_out1 XOR Logical_Operator_out3453_out1;

  Logical_Operator_out4470_out1 <= Logical_Operator_out3446_out1 XOR Logical_Operator_out3454_out1;

  Logical_Operator_out4471_out1 <= Logical_Operator_out3447_out1 XOR Logical_Operator_out3455_out1;

  Logical_Operator_out4472_out1 <= Logical_Operator_out3448_out1 XOR Logical_Operator_out3456_out1;

  Logical_Operator_out4473_out1 <= Logical_Operator_out2421_out1 XOR Logical_Operator_out2429_out1;

  Logical_Operator_out4474_out1 <= Logical_Operator_out2422_out1 XOR Logical_Operator_out2430_out1;

  Logical_Operator_out4475_out1 <= Logical_Operator_out2423_out1 XOR Logical_Operator_out2431_out1;

  Logical_Operator_out4476_out1 <= Logical_Operator_out2424_out1 XOR Logical_Operator_out2432_out1;

  Logical_Operator_out4477_out1 <= Logical_Operator_out1399_out1 XOR Logical_Operator_out1407_out1;

  Logical_Operator_out4478_out1 <= Logical_Operator_out1400_out1 XOR Logical_Operator_out1408_out1;

  Logical_Operator_out4479_out1 <= Logical_Operator_out376_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out4480_out1 <= in752 XOR in768;

  Logical_Operator_out4481_out1 <= Logical_Operator_out3457_out1 XOR Logical_Operator_out3465_out1;

  Logical_Operator_out4482_out1 <= Logical_Operator_out3458_out1 XOR Logical_Operator_out3466_out1;

  Logical_Operator_out4483_out1 <= Logical_Operator_out3459_out1 XOR Logical_Operator_out3467_out1;

  Logical_Operator_out4484_out1 <= Logical_Operator_out3460_out1 XOR Logical_Operator_out3468_out1;

  Logical_Operator_out4485_out1 <= Logical_Operator_out3461_out1 XOR Logical_Operator_out3469_out1;

  Logical_Operator_out4486_out1 <= Logical_Operator_out3462_out1 XOR Logical_Operator_out3470_out1;

  Logical_Operator_out4487_out1 <= Logical_Operator_out3463_out1 XOR Logical_Operator_out3471_out1;

  Logical_Operator_out4488_out1 <= Logical_Operator_out3464_out1 XOR Logical_Operator_out3472_out1;

  Logical_Operator_out4489_out1 <= Logical_Operator_out2437_out1 XOR Logical_Operator_out2445_out1;

  Logical_Operator_out4490_out1 <= Logical_Operator_out2438_out1 XOR Logical_Operator_out2446_out1;

  Logical_Operator_out4491_out1 <= Logical_Operator_out2439_out1 XOR Logical_Operator_out2447_out1;

  Logical_Operator_out4492_out1 <= Logical_Operator_out2440_out1 XOR Logical_Operator_out2448_out1;

  Logical_Operator_out4493_out1 <= Logical_Operator_out1415_out1 XOR Logical_Operator_out1423_out1;

  Logical_Operator_out4494_out1 <= Logical_Operator_out1416_out1 XOR Logical_Operator_out1424_out1;

  Logical_Operator_out4495_out1 <= Logical_Operator_out392_out1 XOR Logical_Operator_out400_out1;

  Logical_Operator_out4496_out1 <= in784 XOR in800;

  Logical_Operator_out4497_out1 <= Logical_Operator_out3473_out1 XOR Logical_Operator_out3481_out1;

  Logical_Operator_out4498_out1 <= Logical_Operator_out3474_out1 XOR Logical_Operator_out3482_out1;

  Logical_Operator_out4499_out1 <= Logical_Operator_out3475_out1 XOR Logical_Operator_out3483_out1;

  Logical_Operator_out4500_out1 <= Logical_Operator_out3476_out1 XOR Logical_Operator_out3484_out1;

  Logical_Operator_out4501_out1 <= Logical_Operator_out3477_out1 XOR Logical_Operator_out3485_out1;

  Logical_Operator_out4502_out1 <= Logical_Operator_out3478_out1 XOR Logical_Operator_out3486_out1;

  Logical_Operator_out4503_out1 <= Logical_Operator_out3479_out1 XOR Logical_Operator_out3487_out1;

  Logical_Operator_out4504_out1 <= Logical_Operator_out3480_out1 XOR Logical_Operator_out3488_out1;

  Logical_Operator_out4505_out1 <= Logical_Operator_out2453_out1 XOR Logical_Operator_out2461_out1;

  Logical_Operator_out4506_out1 <= Logical_Operator_out2454_out1 XOR Logical_Operator_out2462_out1;

  Logical_Operator_out4507_out1 <= Logical_Operator_out2455_out1 XOR Logical_Operator_out2463_out1;

  Logical_Operator_out4508_out1 <= Logical_Operator_out2456_out1 XOR Logical_Operator_out2464_out1;

  Logical_Operator_out4509_out1 <= Logical_Operator_out1431_out1 XOR Logical_Operator_out1439_out1;

  Logical_Operator_out4510_out1 <= Logical_Operator_out1432_out1 XOR Logical_Operator_out1440_out1;

  Logical_Operator_out4511_out1 <= Logical_Operator_out408_out1 XOR Logical_Operator_out416_out1;

  Logical_Operator_out4512_out1 <= in816 XOR in832;

  Logical_Operator_out4513_out1 <= Logical_Operator_out3489_out1 XOR Logical_Operator_out3497_out1;

  Logical_Operator_out4514_out1 <= Logical_Operator_out3490_out1 XOR Logical_Operator_out3498_out1;

  Logical_Operator_out4515_out1 <= Logical_Operator_out3491_out1 XOR Logical_Operator_out3499_out1;

  Logical_Operator_out4516_out1 <= Logical_Operator_out3492_out1 XOR Logical_Operator_out3500_out1;

  Logical_Operator_out4517_out1 <= Logical_Operator_out3493_out1 XOR Logical_Operator_out3501_out1;

  Logical_Operator_out4518_out1 <= Logical_Operator_out3494_out1 XOR Logical_Operator_out3502_out1;

  Logical_Operator_out4519_out1 <= Logical_Operator_out3495_out1 XOR Logical_Operator_out3503_out1;

  Logical_Operator_out4520_out1 <= Logical_Operator_out3496_out1 XOR Logical_Operator_out3504_out1;

  Logical_Operator_out4521_out1 <= Logical_Operator_out2469_out1 XOR Logical_Operator_out2477_out1;

  Logical_Operator_out4522_out1 <= Logical_Operator_out2470_out1 XOR Logical_Operator_out2478_out1;

  Logical_Operator_out4523_out1 <= Logical_Operator_out2471_out1 XOR Logical_Operator_out2479_out1;

  Logical_Operator_out4524_out1 <= Logical_Operator_out2472_out1 XOR Logical_Operator_out2480_out1;

  Logical_Operator_out4525_out1 <= Logical_Operator_out1447_out1 XOR Logical_Operator_out1455_out1;

  Logical_Operator_out4526_out1 <= Logical_Operator_out1448_out1 XOR Logical_Operator_out1456_out1;

  Logical_Operator_out4527_out1 <= Logical_Operator_out424_out1 XOR Logical_Operator_out432_out1;

  Logical_Operator_out4528_out1 <= in848 XOR in864;

  Logical_Operator_out4529_out1 <= Logical_Operator_out3505_out1 XOR Logical_Operator_out3513_out1;

  Logical_Operator_out4530_out1 <= Logical_Operator_out3506_out1 XOR Logical_Operator_out3514_out1;

  Logical_Operator_out4531_out1 <= Logical_Operator_out3507_out1 XOR Logical_Operator_out3515_out1;

  Logical_Operator_out4532_out1 <= Logical_Operator_out3508_out1 XOR Logical_Operator_out3516_out1;

  Logical_Operator_out4533_out1 <= Logical_Operator_out3509_out1 XOR Logical_Operator_out3517_out1;

  Logical_Operator_out4534_out1 <= Logical_Operator_out3510_out1 XOR Logical_Operator_out3518_out1;

  Logical_Operator_out4535_out1 <= Logical_Operator_out3511_out1 XOR Logical_Operator_out3519_out1;

  Logical_Operator_out4536_out1 <= Logical_Operator_out3512_out1 XOR Logical_Operator_out3520_out1;

  Logical_Operator_out4537_out1 <= Logical_Operator_out2485_out1 XOR Logical_Operator_out2493_out1;

  Logical_Operator_out4538_out1 <= Logical_Operator_out2486_out1 XOR Logical_Operator_out2494_out1;

  Logical_Operator_out4539_out1 <= Logical_Operator_out2487_out1 XOR Logical_Operator_out2495_out1;

  Logical_Operator_out4540_out1 <= Logical_Operator_out2488_out1 XOR Logical_Operator_out2496_out1;

  Logical_Operator_out4541_out1 <= Logical_Operator_out1463_out1 XOR Logical_Operator_out1471_out1;

  Logical_Operator_out4542_out1 <= Logical_Operator_out1464_out1 XOR Logical_Operator_out1472_out1;

  Logical_Operator_out4543_out1 <= Logical_Operator_out440_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out4544_out1 <= in880 XOR in896;

  Logical_Operator_out4545_out1 <= Logical_Operator_out3521_out1 XOR Logical_Operator_out3529_out1;

  Logical_Operator_out4546_out1 <= Logical_Operator_out3522_out1 XOR Logical_Operator_out3530_out1;

  Logical_Operator_out4547_out1 <= Logical_Operator_out3523_out1 XOR Logical_Operator_out3531_out1;

  Logical_Operator_out4548_out1 <= Logical_Operator_out3524_out1 XOR Logical_Operator_out3532_out1;

  Logical_Operator_out4549_out1 <= Logical_Operator_out3525_out1 XOR Logical_Operator_out3533_out1;

  Logical_Operator_out4550_out1 <= Logical_Operator_out3526_out1 XOR Logical_Operator_out3534_out1;

  Logical_Operator_out4551_out1 <= Logical_Operator_out3527_out1 XOR Logical_Operator_out3535_out1;

  Logical_Operator_out4552_out1 <= Logical_Operator_out3528_out1 XOR Logical_Operator_out3536_out1;

  Logical_Operator_out4553_out1 <= Logical_Operator_out2501_out1 XOR Logical_Operator_out2509_out1;

  Logical_Operator_out4554_out1 <= Logical_Operator_out2502_out1 XOR Logical_Operator_out2510_out1;

  Logical_Operator_out4555_out1 <= Logical_Operator_out2503_out1 XOR Logical_Operator_out2511_out1;

  Logical_Operator_out4556_out1 <= Logical_Operator_out2504_out1 XOR Logical_Operator_out2512_out1;

  Logical_Operator_out4557_out1 <= Logical_Operator_out1479_out1 XOR Logical_Operator_out1487_out1;

  Logical_Operator_out4558_out1 <= Logical_Operator_out1480_out1 XOR Logical_Operator_out1488_out1;

  Logical_Operator_out4559_out1 <= Logical_Operator_out456_out1 XOR Logical_Operator_out464_out1;

  Logical_Operator_out4560_out1 <= in912 XOR in928;

  Logical_Operator_out4561_out1 <= Logical_Operator_out3537_out1 XOR Logical_Operator_out3545_out1;

  Logical_Operator_out4562_out1 <= Logical_Operator_out3538_out1 XOR Logical_Operator_out3546_out1;

  Logical_Operator_out4563_out1 <= Logical_Operator_out3539_out1 XOR Logical_Operator_out3547_out1;

  Logical_Operator_out4564_out1 <= Logical_Operator_out3540_out1 XOR Logical_Operator_out3548_out1;

  Logical_Operator_out4565_out1 <= Logical_Operator_out3541_out1 XOR Logical_Operator_out3549_out1;

  Logical_Operator_out4566_out1 <= Logical_Operator_out3542_out1 XOR Logical_Operator_out3550_out1;

  Logical_Operator_out4567_out1 <= Logical_Operator_out3543_out1 XOR Logical_Operator_out3551_out1;

  Logical_Operator_out4568_out1 <= Logical_Operator_out3544_out1 XOR Logical_Operator_out3552_out1;

  Logical_Operator_out4569_out1 <= Logical_Operator_out2517_out1 XOR Logical_Operator_out2525_out1;

  Logical_Operator_out4570_out1 <= Logical_Operator_out2518_out1 XOR Logical_Operator_out2526_out1;

  Logical_Operator_out4571_out1 <= Logical_Operator_out2519_out1 XOR Logical_Operator_out2527_out1;

  Logical_Operator_out4572_out1 <= Logical_Operator_out2520_out1 XOR Logical_Operator_out2528_out1;

  Logical_Operator_out4573_out1 <= Logical_Operator_out1495_out1 XOR Logical_Operator_out1503_out1;

  Logical_Operator_out4574_out1 <= Logical_Operator_out1496_out1 XOR Logical_Operator_out1504_out1;

  Logical_Operator_out4575_out1 <= Logical_Operator_out472_out1 XOR Logical_Operator_out480_out1;

  Logical_Operator_out4576_out1 <= in944 XOR in960;

  Logical_Operator_out4577_out1 <= Logical_Operator_out3553_out1 XOR Logical_Operator_out3561_out1;

  Logical_Operator_out4578_out1 <= Logical_Operator_out3554_out1 XOR Logical_Operator_out3562_out1;

  Logical_Operator_out4579_out1 <= Logical_Operator_out3555_out1 XOR Logical_Operator_out3563_out1;

  Logical_Operator_out4580_out1 <= Logical_Operator_out3556_out1 XOR Logical_Operator_out3564_out1;

  Logical_Operator_out4581_out1 <= Logical_Operator_out3557_out1 XOR Logical_Operator_out3565_out1;

  Logical_Operator_out4582_out1 <= Logical_Operator_out3558_out1 XOR Logical_Operator_out3566_out1;

  Logical_Operator_out4583_out1 <= Logical_Operator_out3559_out1 XOR Logical_Operator_out3567_out1;

  Logical_Operator_out4584_out1 <= Logical_Operator_out3560_out1 XOR Logical_Operator_out3568_out1;

  Logical_Operator_out4585_out1 <= Logical_Operator_out2533_out1 XOR Logical_Operator_out2541_out1;

  Logical_Operator_out4586_out1 <= Logical_Operator_out2534_out1 XOR Logical_Operator_out2542_out1;

  Logical_Operator_out4587_out1 <= Logical_Operator_out2535_out1 XOR Logical_Operator_out2543_out1;

  Logical_Operator_out4588_out1 <= Logical_Operator_out2536_out1 XOR Logical_Operator_out2544_out1;

  Logical_Operator_out4589_out1 <= Logical_Operator_out1511_out1 XOR Logical_Operator_out1519_out1;

  Logical_Operator_out4590_out1 <= Logical_Operator_out1512_out1 XOR Logical_Operator_out1520_out1;

  Logical_Operator_out4591_out1 <= Logical_Operator_out488_out1 XOR Logical_Operator_out496_out1;

  Logical_Operator_out4592_out1 <= in976 XOR in992;

  Logical_Operator_out4593_out1 <= Logical_Operator_out3569_out1 XOR Logical_Operator_out3577_out1;

  Logical_Operator_out4594_out1 <= Logical_Operator_out3570_out1 XOR Logical_Operator_out3578_out1;

  Logical_Operator_out4595_out1 <= Logical_Operator_out3571_out1 XOR Logical_Operator_out3579_out1;

  Logical_Operator_out4596_out1 <= Logical_Operator_out3572_out1 XOR Logical_Operator_out3580_out1;

  Logical_Operator_out4597_out1 <= Logical_Operator_out3573_out1 XOR Logical_Operator_out3581_out1;

  Logical_Operator_out4598_out1 <= Logical_Operator_out3574_out1 XOR Logical_Operator_out3582_out1;

  Logical_Operator_out4599_out1 <= Logical_Operator_out3575_out1 XOR Logical_Operator_out3583_out1;

  Logical_Operator_out4600_out1 <= Logical_Operator_out3576_out1 XOR Logical_Operator_out3584_out1;

  Logical_Operator_out4601_out1 <= Logical_Operator_out2549_out1 XOR Logical_Operator_out2557_out1;

  Logical_Operator_out4602_out1 <= Logical_Operator_out2550_out1 XOR Logical_Operator_out2558_out1;

  Logical_Operator_out4603_out1 <= Logical_Operator_out2551_out1 XOR Logical_Operator_out2559_out1;

  Logical_Operator_out4604_out1 <= Logical_Operator_out2552_out1 XOR Logical_Operator_out2560_out1;

  Logical_Operator_out4605_out1 <= Logical_Operator_out1527_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out4606_out1 <= Logical_Operator_out1528_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out4607_out1 <= Logical_Operator_out504_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out4608_out1 <= in1008 XOR in1024;

  Logical_Operator_out4609_out1 <= Logical_Operator_out3585_out1 XOR Logical_Operator_out3593_out1;

  Logical_Operator_out4610_out1 <= Logical_Operator_out3586_out1 XOR Logical_Operator_out3594_out1;

  Logical_Operator_out4611_out1 <= Logical_Operator_out3587_out1 XOR Logical_Operator_out3595_out1;

  Logical_Operator_out4612_out1 <= Logical_Operator_out3588_out1 XOR Logical_Operator_out3596_out1;

  Logical_Operator_out4613_out1 <= Logical_Operator_out3589_out1 XOR Logical_Operator_out3597_out1;

  Logical_Operator_out4614_out1 <= Logical_Operator_out3590_out1 XOR Logical_Operator_out3598_out1;

  Logical_Operator_out4615_out1 <= Logical_Operator_out3591_out1 XOR Logical_Operator_out3599_out1;

  Logical_Operator_out4616_out1 <= Logical_Operator_out3592_out1 XOR Logical_Operator_out3600_out1;

  Logical_Operator_out4617_out1 <= Logical_Operator_out2565_out1 XOR Logical_Operator_out2573_out1;

  Logical_Operator_out4618_out1 <= Logical_Operator_out2566_out1 XOR Logical_Operator_out2574_out1;

  Logical_Operator_out4619_out1 <= Logical_Operator_out2567_out1 XOR Logical_Operator_out2575_out1;

  Logical_Operator_out4620_out1 <= Logical_Operator_out2568_out1 XOR Logical_Operator_out2576_out1;

  Logical_Operator_out4621_out1 <= Logical_Operator_out1543_out1 XOR Logical_Operator_out1551_out1;

  Logical_Operator_out4622_out1 <= Logical_Operator_out1544_out1 XOR Logical_Operator_out1552_out1;

  Logical_Operator_out4623_out1 <= Logical_Operator_out520_out1 XOR Logical_Operator_out528_out1;

  Logical_Operator_out4624_out1 <= in1040 XOR in1056;

  Logical_Operator_out4625_out1 <= Logical_Operator_out3601_out1 XOR Logical_Operator_out3609_out1;

  Logical_Operator_out4626_out1 <= Logical_Operator_out3602_out1 XOR Logical_Operator_out3610_out1;

  Logical_Operator_out4627_out1 <= Logical_Operator_out3603_out1 XOR Logical_Operator_out3611_out1;

  Logical_Operator_out4628_out1 <= Logical_Operator_out3604_out1 XOR Logical_Operator_out3612_out1;

  Logical_Operator_out4629_out1 <= Logical_Operator_out3605_out1 XOR Logical_Operator_out3613_out1;

  Logical_Operator_out4630_out1 <= Logical_Operator_out3606_out1 XOR Logical_Operator_out3614_out1;

  Logical_Operator_out4631_out1 <= Logical_Operator_out3607_out1 XOR Logical_Operator_out3615_out1;

  Logical_Operator_out4632_out1 <= Logical_Operator_out3608_out1 XOR Logical_Operator_out3616_out1;

  Logical_Operator_out4633_out1 <= Logical_Operator_out2581_out1 XOR Logical_Operator_out2589_out1;

  Logical_Operator_out4634_out1 <= Logical_Operator_out2582_out1 XOR Logical_Operator_out2590_out1;

  Logical_Operator_out4635_out1 <= Logical_Operator_out2583_out1 XOR Logical_Operator_out2591_out1;

  Logical_Operator_out4636_out1 <= Logical_Operator_out2584_out1 XOR Logical_Operator_out2592_out1;

  Logical_Operator_out4637_out1 <= Logical_Operator_out1559_out1 XOR Logical_Operator_out1567_out1;

  Logical_Operator_out4638_out1 <= Logical_Operator_out1560_out1 XOR Logical_Operator_out1568_out1;

  Logical_Operator_out4639_out1 <= Logical_Operator_out536_out1 XOR Logical_Operator_out544_out1;

  Logical_Operator_out4640_out1 <= in1072 XOR in1088;

  Logical_Operator_out4641_out1 <= Logical_Operator_out3617_out1 XOR Logical_Operator_out3625_out1;

  Logical_Operator_out4642_out1 <= Logical_Operator_out3618_out1 XOR Logical_Operator_out3626_out1;

  Logical_Operator_out4643_out1 <= Logical_Operator_out3619_out1 XOR Logical_Operator_out3627_out1;

  Logical_Operator_out4644_out1 <= Logical_Operator_out3620_out1 XOR Logical_Operator_out3628_out1;

  Logical_Operator_out4645_out1 <= Logical_Operator_out3621_out1 XOR Logical_Operator_out3629_out1;

  Logical_Operator_out4646_out1 <= Logical_Operator_out3622_out1 XOR Logical_Operator_out3630_out1;

  Logical_Operator_out4647_out1 <= Logical_Operator_out3623_out1 XOR Logical_Operator_out3631_out1;

  Logical_Operator_out4648_out1 <= Logical_Operator_out3624_out1 XOR Logical_Operator_out3632_out1;

  Logical_Operator_out4649_out1 <= Logical_Operator_out2597_out1 XOR Logical_Operator_out2605_out1;

  Logical_Operator_out4650_out1 <= Logical_Operator_out2598_out1 XOR Logical_Operator_out2606_out1;

  Logical_Operator_out4651_out1 <= Logical_Operator_out2599_out1 XOR Logical_Operator_out2607_out1;

  Logical_Operator_out4652_out1 <= Logical_Operator_out2600_out1 XOR Logical_Operator_out2608_out1;

  Logical_Operator_out4653_out1 <= Logical_Operator_out1575_out1 XOR Logical_Operator_out1583_out1;

  Logical_Operator_out4654_out1 <= Logical_Operator_out1576_out1 XOR Logical_Operator_out1584_out1;

  Logical_Operator_out4655_out1 <= Logical_Operator_out552_out1 XOR Logical_Operator_out560_out1;

  Logical_Operator_out4656_out1 <= in1104 XOR in1120;

  Logical_Operator_out4657_out1 <= Logical_Operator_out3633_out1 XOR Logical_Operator_out3641_out1;

  Logical_Operator_out4658_out1 <= Logical_Operator_out3634_out1 XOR Logical_Operator_out3642_out1;

  Logical_Operator_out4659_out1 <= Logical_Operator_out3635_out1 XOR Logical_Operator_out3643_out1;

  Logical_Operator_out4660_out1 <= Logical_Operator_out3636_out1 XOR Logical_Operator_out3644_out1;

  Logical_Operator_out4661_out1 <= Logical_Operator_out3637_out1 XOR Logical_Operator_out3645_out1;

  Logical_Operator_out4662_out1 <= Logical_Operator_out3638_out1 XOR Logical_Operator_out3646_out1;

  Logical_Operator_out4663_out1 <= Logical_Operator_out3639_out1 XOR Logical_Operator_out3647_out1;

  Logical_Operator_out4664_out1 <= Logical_Operator_out3640_out1 XOR Logical_Operator_out3648_out1;

  Logical_Operator_out4665_out1 <= Logical_Operator_out2613_out1 XOR Logical_Operator_out2621_out1;

  Logical_Operator_out4666_out1 <= Logical_Operator_out2614_out1 XOR Logical_Operator_out2622_out1;

  Logical_Operator_out4667_out1 <= Logical_Operator_out2615_out1 XOR Logical_Operator_out2623_out1;

  Logical_Operator_out4668_out1 <= Logical_Operator_out2616_out1 XOR Logical_Operator_out2624_out1;

  Logical_Operator_out4669_out1 <= Logical_Operator_out1591_out1 XOR Logical_Operator_out1599_out1;

  Logical_Operator_out4670_out1 <= Logical_Operator_out1592_out1 XOR Logical_Operator_out1600_out1;

  Logical_Operator_out4671_out1 <= Logical_Operator_out568_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out4672_out1 <= in1136 XOR in1152;

  Logical_Operator_out4673_out1 <= Logical_Operator_out3649_out1 XOR Logical_Operator_out3657_out1;

  Logical_Operator_out4674_out1 <= Logical_Operator_out3650_out1 XOR Logical_Operator_out3658_out1;

  Logical_Operator_out4675_out1 <= Logical_Operator_out3651_out1 XOR Logical_Operator_out3659_out1;

  Logical_Operator_out4676_out1 <= Logical_Operator_out3652_out1 XOR Logical_Operator_out3660_out1;

  Logical_Operator_out4677_out1 <= Logical_Operator_out3653_out1 XOR Logical_Operator_out3661_out1;

  Logical_Operator_out4678_out1 <= Logical_Operator_out3654_out1 XOR Logical_Operator_out3662_out1;

  Logical_Operator_out4679_out1 <= Logical_Operator_out3655_out1 XOR Logical_Operator_out3663_out1;

  Logical_Operator_out4680_out1 <= Logical_Operator_out3656_out1 XOR Logical_Operator_out3664_out1;

  Logical_Operator_out4681_out1 <= Logical_Operator_out2629_out1 XOR Logical_Operator_out2637_out1;

  Logical_Operator_out4682_out1 <= Logical_Operator_out2630_out1 XOR Logical_Operator_out2638_out1;

  Logical_Operator_out4683_out1 <= Logical_Operator_out2631_out1 XOR Logical_Operator_out2639_out1;

  Logical_Operator_out4684_out1 <= Logical_Operator_out2632_out1 XOR Logical_Operator_out2640_out1;

  Logical_Operator_out4685_out1 <= Logical_Operator_out1607_out1 XOR Logical_Operator_out1615_out1;

  Logical_Operator_out4686_out1 <= Logical_Operator_out1608_out1 XOR Logical_Operator_out1616_out1;

  Logical_Operator_out4687_out1 <= Logical_Operator_out584_out1 XOR Logical_Operator_out592_out1;

  Logical_Operator_out4688_out1 <= in1168 XOR in1184;

  Logical_Operator_out4689_out1 <= Logical_Operator_out3665_out1 XOR Logical_Operator_out3673_out1;

  Logical_Operator_out4690_out1 <= Logical_Operator_out3666_out1 XOR Logical_Operator_out3674_out1;

  Logical_Operator_out4691_out1 <= Logical_Operator_out3667_out1 XOR Logical_Operator_out3675_out1;

  Logical_Operator_out4692_out1 <= Logical_Operator_out3668_out1 XOR Logical_Operator_out3676_out1;

  Logical_Operator_out4693_out1 <= Logical_Operator_out3669_out1 XOR Logical_Operator_out3677_out1;

  Logical_Operator_out4694_out1 <= Logical_Operator_out3670_out1 XOR Logical_Operator_out3678_out1;

  Logical_Operator_out4695_out1 <= Logical_Operator_out3671_out1 XOR Logical_Operator_out3679_out1;

  Logical_Operator_out4696_out1 <= Logical_Operator_out3672_out1 XOR Logical_Operator_out3680_out1;

  Logical_Operator_out4697_out1 <= Logical_Operator_out2645_out1 XOR Logical_Operator_out2653_out1;

  Logical_Operator_out4698_out1 <= Logical_Operator_out2646_out1 XOR Logical_Operator_out2654_out1;

  Logical_Operator_out4699_out1 <= Logical_Operator_out2647_out1 XOR Logical_Operator_out2655_out1;

  Logical_Operator_out4700_out1 <= Logical_Operator_out2648_out1 XOR Logical_Operator_out2656_out1;

  Logical_Operator_out4701_out1 <= Logical_Operator_out1623_out1 XOR Logical_Operator_out1631_out1;

  Logical_Operator_out4702_out1 <= Logical_Operator_out1624_out1 XOR Logical_Operator_out1632_out1;

  Logical_Operator_out4703_out1 <= Logical_Operator_out600_out1 XOR Logical_Operator_out608_out1;

  Logical_Operator_out4704_out1 <= in1200 XOR in1216;

  Logical_Operator_out4705_out1 <= Logical_Operator_out3681_out1 XOR Logical_Operator_out3689_out1;

  Logical_Operator_out4706_out1 <= Logical_Operator_out3682_out1 XOR Logical_Operator_out3690_out1;

  Logical_Operator_out4707_out1 <= Logical_Operator_out3683_out1 XOR Logical_Operator_out3691_out1;

  Logical_Operator_out4708_out1 <= Logical_Operator_out3684_out1 XOR Logical_Operator_out3692_out1;

  Logical_Operator_out4709_out1 <= Logical_Operator_out3685_out1 XOR Logical_Operator_out3693_out1;

  Logical_Operator_out4710_out1 <= Logical_Operator_out3686_out1 XOR Logical_Operator_out3694_out1;

  Logical_Operator_out4711_out1 <= Logical_Operator_out3687_out1 XOR Logical_Operator_out3695_out1;

  Logical_Operator_out4712_out1 <= Logical_Operator_out3688_out1 XOR Logical_Operator_out3696_out1;

  Logical_Operator_out4713_out1 <= Logical_Operator_out2661_out1 XOR Logical_Operator_out2669_out1;

  Logical_Operator_out4714_out1 <= Logical_Operator_out2662_out1 XOR Logical_Operator_out2670_out1;

  Logical_Operator_out4715_out1 <= Logical_Operator_out2663_out1 XOR Logical_Operator_out2671_out1;

  Logical_Operator_out4716_out1 <= Logical_Operator_out2664_out1 XOR Logical_Operator_out2672_out1;

  Logical_Operator_out4717_out1 <= Logical_Operator_out1639_out1 XOR Logical_Operator_out1647_out1;

  Logical_Operator_out4718_out1 <= Logical_Operator_out1640_out1 XOR Logical_Operator_out1648_out1;

  Logical_Operator_out4719_out1 <= Logical_Operator_out616_out1 XOR Logical_Operator_out624_out1;

  Logical_Operator_out4720_out1 <= in1232 XOR in1248;

  Logical_Operator_out4721_out1 <= Logical_Operator_out3697_out1 XOR Logical_Operator_out3705_out1;

  Logical_Operator_out4722_out1 <= Logical_Operator_out3698_out1 XOR Logical_Operator_out3706_out1;

  Logical_Operator_out4723_out1 <= Logical_Operator_out3699_out1 XOR Logical_Operator_out3707_out1;

  Logical_Operator_out4724_out1 <= Logical_Operator_out3700_out1 XOR Logical_Operator_out3708_out1;

  Logical_Operator_out4725_out1 <= Logical_Operator_out3701_out1 XOR Logical_Operator_out3709_out1;

  Logical_Operator_out4726_out1 <= Logical_Operator_out3702_out1 XOR Logical_Operator_out3710_out1;

  Logical_Operator_out4727_out1 <= Logical_Operator_out3703_out1 XOR Logical_Operator_out3711_out1;

  Logical_Operator_out4728_out1 <= Logical_Operator_out3704_out1 XOR Logical_Operator_out3712_out1;

  Logical_Operator_out4729_out1 <= Logical_Operator_out2677_out1 XOR Logical_Operator_out2685_out1;

  Logical_Operator_out4730_out1 <= Logical_Operator_out2678_out1 XOR Logical_Operator_out2686_out1;

  Logical_Operator_out4731_out1 <= Logical_Operator_out2679_out1 XOR Logical_Operator_out2687_out1;

  Logical_Operator_out4732_out1 <= Logical_Operator_out2680_out1 XOR Logical_Operator_out2688_out1;

  Logical_Operator_out4733_out1 <= Logical_Operator_out1655_out1 XOR Logical_Operator_out1663_out1;

  Logical_Operator_out4734_out1 <= Logical_Operator_out1656_out1 XOR Logical_Operator_out1664_out1;

  Logical_Operator_out4735_out1 <= Logical_Operator_out632_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out4736_out1 <= in1264 XOR in1280;

  Logical_Operator_out4737_out1 <= Logical_Operator_out3713_out1 XOR Logical_Operator_out3721_out1;

  Logical_Operator_out4738_out1 <= Logical_Operator_out3714_out1 XOR Logical_Operator_out3722_out1;

  Logical_Operator_out4739_out1 <= Logical_Operator_out3715_out1 XOR Logical_Operator_out3723_out1;

  Logical_Operator_out4740_out1 <= Logical_Operator_out3716_out1 XOR Logical_Operator_out3724_out1;

  Logical_Operator_out4741_out1 <= Logical_Operator_out3717_out1 XOR Logical_Operator_out3725_out1;

  Logical_Operator_out4742_out1 <= Logical_Operator_out3718_out1 XOR Logical_Operator_out3726_out1;

  Logical_Operator_out4743_out1 <= Logical_Operator_out3719_out1 XOR Logical_Operator_out3727_out1;

  Logical_Operator_out4744_out1 <= Logical_Operator_out3720_out1 XOR Logical_Operator_out3728_out1;

  Logical_Operator_out4745_out1 <= Logical_Operator_out2693_out1 XOR Logical_Operator_out2701_out1;

  Logical_Operator_out4746_out1 <= Logical_Operator_out2694_out1 XOR Logical_Operator_out2702_out1;

  Logical_Operator_out4747_out1 <= Logical_Operator_out2695_out1 XOR Logical_Operator_out2703_out1;

  Logical_Operator_out4748_out1 <= Logical_Operator_out2696_out1 XOR Logical_Operator_out2704_out1;

  Logical_Operator_out4749_out1 <= Logical_Operator_out1671_out1 XOR Logical_Operator_out1679_out1;

  Logical_Operator_out4750_out1 <= Logical_Operator_out1672_out1 XOR Logical_Operator_out1680_out1;

  Logical_Operator_out4751_out1 <= Logical_Operator_out648_out1 XOR Logical_Operator_out656_out1;

  Logical_Operator_out4752_out1 <= in1296 XOR in1312;

  Logical_Operator_out4753_out1 <= Logical_Operator_out3729_out1 XOR Logical_Operator_out3737_out1;

  Logical_Operator_out4754_out1 <= Logical_Operator_out3730_out1 XOR Logical_Operator_out3738_out1;

  Logical_Operator_out4755_out1 <= Logical_Operator_out3731_out1 XOR Logical_Operator_out3739_out1;

  Logical_Operator_out4756_out1 <= Logical_Operator_out3732_out1 XOR Logical_Operator_out3740_out1;

  Logical_Operator_out4757_out1 <= Logical_Operator_out3733_out1 XOR Logical_Operator_out3741_out1;

  Logical_Operator_out4758_out1 <= Logical_Operator_out3734_out1 XOR Logical_Operator_out3742_out1;

  Logical_Operator_out4759_out1 <= Logical_Operator_out3735_out1 XOR Logical_Operator_out3743_out1;

  Logical_Operator_out4760_out1 <= Logical_Operator_out3736_out1 XOR Logical_Operator_out3744_out1;

  Logical_Operator_out4761_out1 <= Logical_Operator_out2709_out1 XOR Logical_Operator_out2717_out1;

  Logical_Operator_out4762_out1 <= Logical_Operator_out2710_out1 XOR Logical_Operator_out2718_out1;

  Logical_Operator_out4763_out1 <= Logical_Operator_out2711_out1 XOR Logical_Operator_out2719_out1;

  Logical_Operator_out4764_out1 <= Logical_Operator_out2712_out1 XOR Logical_Operator_out2720_out1;

  Logical_Operator_out4765_out1 <= Logical_Operator_out1687_out1 XOR Logical_Operator_out1695_out1;

  Logical_Operator_out4766_out1 <= Logical_Operator_out1688_out1 XOR Logical_Operator_out1696_out1;

  Logical_Operator_out4767_out1 <= Logical_Operator_out664_out1 XOR Logical_Operator_out672_out1;

  Logical_Operator_out4768_out1 <= in1328 XOR in1344;

  Logical_Operator_out4769_out1 <= Logical_Operator_out3745_out1 XOR Logical_Operator_out3753_out1;

  Logical_Operator_out4770_out1 <= Logical_Operator_out3746_out1 XOR Logical_Operator_out3754_out1;

  Logical_Operator_out4771_out1 <= Logical_Operator_out3747_out1 XOR Logical_Operator_out3755_out1;

  Logical_Operator_out4772_out1 <= Logical_Operator_out3748_out1 XOR Logical_Operator_out3756_out1;

  Logical_Operator_out4773_out1 <= Logical_Operator_out3749_out1 XOR Logical_Operator_out3757_out1;

  Logical_Operator_out4774_out1 <= Logical_Operator_out3750_out1 XOR Logical_Operator_out3758_out1;

  Logical_Operator_out4775_out1 <= Logical_Operator_out3751_out1 XOR Logical_Operator_out3759_out1;

  Logical_Operator_out4776_out1 <= Logical_Operator_out3752_out1 XOR Logical_Operator_out3760_out1;

  Logical_Operator_out4777_out1 <= Logical_Operator_out2725_out1 XOR Logical_Operator_out2733_out1;

  Logical_Operator_out4778_out1 <= Logical_Operator_out2726_out1 XOR Logical_Operator_out2734_out1;

  Logical_Operator_out4779_out1 <= Logical_Operator_out2727_out1 XOR Logical_Operator_out2735_out1;

  Logical_Operator_out4780_out1 <= Logical_Operator_out2728_out1 XOR Logical_Operator_out2736_out1;

  Logical_Operator_out4781_out1 <= Logical_Operator_out1703_out1 XOR Logical_Operator_out1711_out1;

  Logical_Operator_out4782_out1 <= Logical_Operator_out1704_out1 XOR Logical_Operator_out1712_out1;

  Logical_Operator_out4783_out1 <= Logical_Operator_out680_out1 XOR Logical_Operator_out688_out1;

  Logical_Operator_out4784_out1 <= in1360 XOR in1376;

  Logical_Operator_out4785_out1 <= Logical_Operator_out3761_out1 XOR Logical_Operator_out3769_out1;

  Logical_Operator_out4786_out1 <= Logical_Operator_out3762_out1 XOR Logical_Operator_out3770_out1;

  Logical_Operator_out4787_out1 <= Logical_Operator_out3763_out1 XOR Logical_Operator_out3771_out1;

  Logical_Operator_out4788_out1 <= Logical_Operator_out3764_out1 XOR Logical_Operator_out3772_out1;

  Logical_Operator_out4789_out1 <= Logical_Operator_out3765_out1 XOR Logical_Operator_out3773_out1;

  Logical_Operator_out4790_out1 <= Logical_Operator_out3766_out1 XOR Logical_Operator_out3774_out1;

  Logical_Operator_out4791_out1 <= Logical_Operator_out3767_out1 XOR Logical_Operator_out3775_out1;

  Logical_Operator_out4792_out1 <= Logical_Operator_out3768_out1 XOR Logical_Operator_out3776_out1;

  Logical_Operator_out4793_out1 <= Logical_Operator_out2741_out1 XOR Logical_Operator_out2749_out1;

  Logical_Operator_out4794_out1 <= Logical_Operator_out2742_out1 XOR Logical_Operator_out2750_out1;

  Logical_Operator_out4795_out1 <= Logical_Operator_out2743_out1 XOR Logical_Operator_out2751_out1;

  Logical_Operator_out4796_out1 <= Logical_Operator_out2744_out1 XOR Logical_Operator_out2752_out1;

  Logical_Operator_out4797_out1 <= Logical_Operator_out1719_out1 XOR Logical_Operator_out1727_out1;

  Logical_Operator_out4798_out1 <= Logical_Operator_out1720_out1 XOR Logical_Operator_out1728_out1;

  Logical_Operator_out4799_out1 <= Logical_Operator_out696_out1 XOR Logical_Operator_out704_out1;

  Logical_Operator_out4800_out1 <= in1392 XOR in1408;

  Logical_Operator_out4801_out1 <= Logical_Operator_out3777_out1 XOR Logical_Operator_out3785_out1;

  Logical_Operator_out4802_out1 <= Logical_Operator_out3778_out1 XOR Logical_Operator_out3786_out1;

  Logical_Operator_out4803_out1 <= Logical_Operator_out3779_out1 XOR Logical_Operator_out3787_out1;

  Logical_Operator_out4804_out1 <= Logical_Operator_out3780_out1 XOR Logical_Operator_out3788_out1;

  Logical_Operator_out4805_out1 <= Logical_Operator_out3781_out1 XOR Logical_Operator_out3789_out1;

  Logical_Operator_out4806_out1 <= Logical_Operator_out3782_out1 XOR Logical_Operator_out3790_out1;

  Logical_Operator_out4807_out1 <= Logical_Operator_out3783_out1 XOR Logical_Operator_out3791_out1;

  Logical_Operator_out4808_out1 <= Logical_Operator_out3784_out1 XOR Logical_Operator_out3792_out1;

  Logical_Operator_out4809_out1 <= Logical_Operator_out2757_out1 XOR Logical_Operator_out2765_out1;

  Logical_Operator_out4810_out1 <= Logical_Operator_out2758_out1 XOR Logical_Operator_out2766_out1;

  Logical_Operator_out4811_out1 <= Logical_Operator_out2759_out1 XOR Logical_Operator_out2767_out1;

  Logical_Operator_out4812_out1 <= Logical_Operator_out2760_out1 XOR Logical_Operator_out2768_out1;

  Logical_Operator_out4813_out1 <= Logical_Operator_out1735_out1 XOR Logical_Operator_out1743_out1;

  Logical_Operator_out4814_out1 <= Logical_Operator_out1736_out1 XOR Logical_Operator_out1744_out1;

  Logical_Operator_out4815_out1 <= Logical_Operator_out712_out1 XOR Logical_Operator_out720_out1;

  Logical_Operator_out4816_out1 <= in1424 XOR in1440;

  Logical_Operator_out4817_out1 <= Logical_Operator_out3793_out1 XOR Logical_Operator_out3801_out1;

  Logical_Operator_out4818_out1 <= Logical_Operator_out3794_out1 XOR Logical_Operator_out3802_out1;

  Logical_Operator_out4819_out1 <= Logical_Operator_out3795_out1 XOR Logical_Operator_out3803_out1;

  Logical_Operator_out4820_out1 <= Logical_Operator_out3796_out1 XOR Logical_Operator_out3804_out1;

  Logical_Operator_out4821_out1 <= Logical_Operator_out3797_out1 XOR Logical_Operator_out3805_out1;

  Logical_Operator_out4822_out1 <= Logical_Operator_out3798_out1 XOR Logical_Operator_out3806_out1;

  Logical_Operator_out4823_out1 <= Logical_Operator_out3799_out1 XOR Logical_Operator_out3807_out1;

  Logical_Operator_out4824_out1 <= Logical_Operator_out3800_out1 XOR Logical_Operator_out3808_out1;

  Logical_Operator_out4825_out1 <= Logical_Operator_out2773_out1 XOR Logical_Operator_out2781_out1;

  Logical_Operator_out4826_out1 <= Logical_Operator_out2774_out1 XOR Logical_Operator_out2782_out1;

  Logical_Operator_out4827_out1 <= Logical_Operator_out2775_out1 XOR Logical_Operator_out2783_out1;

  Logical_Operator_out4828_out1 <= Logical_Operator_out2776_out1 XOR Logical_Operator_out2784_out1;

  Logical_Operator_out4829_out1 <= Logical_Operator_out1751_out1 XOR Logical_Operator_out1759_out1;

  Logical_Operator_out4830_out1 <= Logical_Operator_out1752_out1 XOR Logical_Operator_out1760_out1;

  Logical_Operator_out4831_out1 <= Logical_Operator_out728_out1 XOR Logical_Operator_out736_out1;

  Logical_Operator_out4832_out1 <= in1456 XOR in1472;

  Logical_Operator_out4833_out1 <= Logical_Operator_out3809_out1 XOR Logical_Operator_out3817_out1;

  Logical_Operator_out4834_out1 <= Logical_Operator_out3810_out1 XOR Logical_Operator_out3818_out1;

  Logical_Operator_out4835_out1 <= Logical_Operator_out3811_out1 XOR Logical_Operator_out3819_out1;

  Logical_Operator_out4836_out1 <= Logical_Operator_out3812_out1 XOR Logical_Operator_out3820_out1;

  Logical_Operator_out4837_out1 <= Logical_Operator_out3813_out1 XOR Logical_Operator_out3821_out1;

  Logical_Operator_out4838_out1 <= Logical_Operator_out3814_out1 XOR Logical_Operator_out3822_out1;

  Logical_Operator_out4839_out1 <= Logical_Operator_out3815_out1 XOR Logical_Operator_out3823_out1;

  Logical_Operator_out4840_out1 <= Logical_Operator_out3816_out1 XOR Logical_Operator_out3824_out1;

  Logical_Operator_out4841_out1 <= Logical_Operator_out2789_out1 XOR Logical_Operator_out2797_out1;

  Logical_Operator_out4842_out1 <= Logical_Operator_out2790_out1 XOR Logical_Operator_out2798_out1;

  Logical_Operator_out4843_out1 <= Logical_Operator_out2791_out1 XOR Logical_Operator_out2799_out1;

  Logical_Operator_out4844_out1 <= Logical_Operator_out2792_out1 XOR Logical_Operator_out2800_out1;

  Logical_Operator_out4845_out1 <= Logical_Operator_out1767_out1 XOR Logical_Operator_out1775_out1;

  Logical_Operator_out4846_out1 <= Logical_Operator_out1768_out1 XOR Logical_Operator_out1776_out1;

  Logical_Operator_out4847_out1 <= Logical_Operator_out744_out1 XOR Logical_Operator_out752_out1;

  Logical_Operator_out4848_out1 <= in1488 XOR in1504;

  Logical_Operator_out4849_out1 <= Logical_Operator_out3825_out1 XOR Logical_Operator_out3833_out1;

  Logical_Operator_out4850_out1 <= Logical_Operator_out3826_out1 XOR Logical_Operator_out3834_out1;

  Logical_Operator_out4851_out1 <= Logical_Operator_out3827_out1 XOR Logical_Operator_out3835_out1;

  Logical_Operator_out4852_out1 <= Logical_Operator_out3828_out1 XOR Logical_Operator_out3836_out1;

  Logical_Operator_out4853_out1 <= Logical_Operator_out3829_out1 XOR Logical_Operator_out3837_out1;

  Logical_Operator_out4854_out1 <= Logical_Operator_out3830_out1 XOR Logical_Operator_out3838_out1;

  Logical_Operator_out4855_out1 <= Logical_Operator_out3831_out1 XOR Logical_Operator_out3839_out1;

  Logical_Operator_out4856_out1 <= Logical_Operator_out3832_out1 XOR Logical_Operator_out3840_out1;

  Logical_Operator_out4857_out1 <= Logical_Operator_out2805_out1 XOR Logical_Operator_out2813_out1;

  Logical_Operator_out4858_out1 <= Logical_Operator_out2806_out1 XOR Logical_Operator_out2814_out1;

  Logical_Operator_out4859_out1 <= Logical_Operator_out2807_out1 XOR Logical_Operator_out2815_out1;

  Logical_Operator_out4860_out1 <= Logical_Operator_out2808_out1 XOR Logical_Operator_out2816_out1;

  Logical_Operator_out4861_out1 <= Logical_Operator_out1783_out1 XOR Logical_Operator_out1791_out1;

  Logical_Operator_out4862_out1 <= Logical_Operator_out1784_out1 XOR Logical_Operator_out1792_out1;

  Logical_Operator_out4863_out1 <= Logical_Operator_out760_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out4864_out1 <= in1520 XOR in1536;

  Logical_Operator_out4865_out1 <= Logical_Operator_out3841_out1 XOR Logical_Operator_out3849_out1;

  Logical_Operator_out4866_out1 <= Logical_Operator_out3842_out1 XOR Logical_Operator_out3850_out1;

  Logical_Operator_out4867_out1 <= Logical_Operator_out3843_out1 XOR Logical_Operator_out3851_out1;

  Logical_Operator_out4868_out1 <= Logical_Operator_out3844_out1 XOR Logical_Operator_out3852_out1;

  Logical_Operator_out4869_out1 <= Logical_Operator_out3845_out1 XOR Logical_Operator_out3853_out1;

  Logical_Operator_out4870_out1 <= Logical_Operator_out3846_out1 XOR Logical_Operator_out3854_out1;

  Logical_Operator_out4871_out1 <= Logical_Operator_out3847_out1 XOR Logical_Operator_out3855_out1;

  Logical_Operator_out4872_out1 <= Logical_Operator_out3848_out1 XOR Logical_Operator_out3856_out1;

  Logical_Operator_out4873_out1 <= Logical_Operator_out2821_out1 XOR Logical_Operator_out2829_out1;

  Logical_Operator_out4874_out1 <= Logical_Operator_out2822_out1 XOR Logical_Operator_out2830_out1;

  Logical_Operator_out4875_out1 <= Logical_Operator_out2823_out1 XOR Logical_Operator_out2831_out1;

  Logical_Operator_out4876_out1 <= Logical_Operator_out2824_out1 XOR Logical_Operator_out2832_out1;

  Logical_Operator_out4877_out1 <= Logical_Operator_out1799_out1 XOR Logical_Operator_out1807_out1;

  Logical_Operator_out4878_out1 <= Logical_Operator_out1800_out1 XOR Logical_Operator_out1808_out1;

  Logical_Operator_out4879_out1 <= Logical_Operator_out776_out1 XOR Logical_Operator_out784_out1;

  Logical_Operator_out4880_out1 <= in1552 XOR in1568;

  Logical_Operator_out4881_out1 <= Logical_Operator_out3857_out1 XOR Logical_Operator_out3865_out1;

  Logical_Operator_out4882_out1 <= Logical_Operator_out3858_out1 XOR Logical_Operator_out3866_out1;

  Logical_Operator_out4883_out1 <= Logical_Operator_out3859_out1 XOR Logical_Operator_out3867_out1;

  Logical_Operator_out4884_out1 <= Logical_Operator_out3860_out1 XOR Logical_Operator_out3868_out1;

  Logical_Operator_out4885_out1 <= Logical_Operator_out3861_out1 XOR Logical_Operator_out3869_out1;

  Logical_Operator_out4886_out1 <= Logical_Operator_out3862_out1 XOR Logical_Operator_out3870_out1;

  Logical_Operator_out4887_out1 <= Logical_Operator_out3863_out1 XOR Logical_Operator_out3871_out1;

  Logical_Operator_out4888_out1 <= Logical_Operator_out3864_out1 XOR Logical_Operator_out3872_out1;

  Logical_Operator_out4889_out1 <= Logical_Operator_out2837_out1 XOR Logical_Operator_out2845_out1;

  Logical_Operator_out4890_out1 <= Logical_Operator_out2838_out1 XOR Logical_Operator_out2846_out1;

  Logical_Operator_out4891_out1 <= Logical_Operator_out2839_out1 XOR Logical_Operator_out2847_out1;

  Logical_Operator_out4892_out1 <= Logical_Operator_out2840_out1 XOR Logical_Operator_out2848_out1;

  Logical_Operator_out4893_out1 <= Logical_Operator_out1815_out1 XOR Logical_Operator_out1823_out1;

  Logical_Operator_out4894_out1 <= Logical_Operator_out1816_out1 XOR Logical_Operator_out1824_out1;

  Logical_Operator_out4895_out1 <= Logical_Operator_out792_out1 XOR Logical_Operator_out800_out1;

  Logical_Operator_out4896_out1 <= in1584 XOR in1600;

  Logical_Operator_out4897_out1 <= Logical_Operator_out3873_out1 XOR Logical_Operator_out3881_out1;

  Logical_Operator_out4898_out1 <= Logical_Operator_out3874_out1 XOR Logical_Operator_out3882_out1;

  Logical_Operator_out4899_out1 <= Logical_Operator_out3875_out1 XOR Logical_Operator_out3883_out1;

  Logical_Operator_out4900_out1 <= Logical_Operator_out3876_out1 XOR Logical_Operator_out3884_out1;

  Logical_Operator_out4901_out1 <= Logical_Operator_out3877_out1 XOR Logical_Operator_out3885_out1;

  Logical_Operator_out4902_out1 <= Logical_Operator_out3878_out1 XOR Logical_Operator_out3886_out1;

  Logical_Operator_out4903_out1 <= Logical_Operator_out3879_out1 XOR Logical_Operator_out3887_out1;

  Logical_Operator_out4904_out1 <= Logical_Operator_out3880_out1 XOR Logical_Operator_out3888_out1;

  Logical_Operator_out4905_out1 <= Logical_Operator_out2853_out1 XOR Logical_Operator_out2861_out1;

  Logical_Operator_out4906_out1 <= Logical_Operator_out2854_out1 XOR Logical_Operator_out2862_out1;

  Logical_Operator_out4907_out1 <= Logical_Operator_out2855_out1 XOR Logical_Operator_out2863_out1;

  Logical_Operator_out4908_out1 <= Logical_Operator_out2856_out1 XOR Logical_Operator_out2864_out1;

  Logical_Operator_out4909_out1 <= Logical_Operator_out1831_out1 XOR Logical_Operator_out1839_out1;

  Logical_Operator_out4910_out1 <= Logical_Operator_out1832_out1 XOR Logical_Operator_out1840_out1;

  Logical_Operator_out4911_out1 <= Logical_Operator_out808_out1 XOR Logical_Operator_out816_out1;

  Logical_Operator_out4912_out1 <= in1616 XOR in1632;

  Logical_Operator_out4913_out1 <= Logical_Operator_out3889_out1 XOR Logical_Operator_out3897_out1;

  Logical_Operator_out4914_out1 <= Logical_Operator_out3890_out1 XOR Logical_Operator_out3898_out1;

  Logical_Operator_out4915_out1 <= Logical_Operator_out3891_out1 XOR Logical_Operator_out3899_out1;

  Logical_Operator_out4916_out1 <= Logical_Operator_out3892_out1 XOR Logical_Operator_out3900_out1;

  Logical_Operator_out4917_out1 <= Logical_Operator_out3893_out1 XOR Logical_Operator_out3901_out1;

  Logical_Operator_out4918_out1 <= Logical_Operator_out3894_out1 XOR Logical_Operator_out3902_out1;

  Logical_Operator_out4919_out1 <= Logical_Operator_out3895_out1 XOR Logical_Operator_out3903_out1;

  Logical_Operator_out4920_out1 <= Logical_Operator_out3896_out1 XOR Logical_Operator_out3904_out1;

  Logical_Operator_out4921_out1 <= Logical_Operator_out2869_out1 XOR Logical_Operator_out2877_out1;

  Logical_Operator_out4922_out1 <= Logical_Operator_out2870_out1 XOR Logical_Operator_out2878_out1;

  Logical_Operator_out4923_out1 <= Logical_Operator_out2871_out1 XOR Logical_Operator_out2879_out1;

  Logical_Operator_out4924_out1 <= Logical_Operator_out2872_out1 XOR Logical_Operator_out2880_out1;

  Logical_Operator_out4925_out1 <= Logical_Operator_out1847_out1 XOR Logical_Operator_out1855_out1;

  Logical_Operator_out4926_out1 <= Logical_Operator_out1848_out1 XOR Logical_Operator_out1856_out1;

  Logical_Operator_out4927_out1 <= Logical_Operator_out824_out1 XOR Logical_Operator_out832_out1;

  Logical_Operator_out4928_out1 <= in1648 XOR in1664;

  Logical_Operator_out4929_out1 <= Logical_Operator_out3905_out1 XOR Logical_Operator_out3913_out1;

  Logical_Operator_out4930_out1 <= Logical_Operator_out3906_out1 XOR Logical_Operator_out3914_out1;

  Logical_Operator_out4931_out1 <= Logical_Operator_out3907_out1 XOR Logical_Operator_out3915_out1;

  Logical_Operator_out4932_out1 <= Logical_Operator_out3908_out1 XOR Logical_Operator_out3916_out1;

  Logical_Operator_out4933_out1 <= Logical_Operator_out3909_out1 XOR Logical_Operator_out3917_out1;

  Logical_Operator_out4934_out1 <= Logical_Operator_out3910_out1 XOR Logical_Operator_out3918_out1;

  Logical_Operator_out4935_out1 <= Logical_Operator_out3911_out1 XOR Logical_Operator_out3919_out1;

  Logical_Operator_out4936_out1 <= Logical_Operator_out3912_out1 XOR Logical_Operator_out3920_out1;

  Logical_Operator_out4937_out1 <= Logical_Operator_out2885_out1 XOR Logical_Operator_out2893_out1;

  Logical_Operator_out4938_out1 <= Logical_Operator_out2886_out1 XOR Logical_Operator_out2894_out1;

  Logical_Operator_out4939_out1 <= Logical_Operator_out2887_out1 XOR Logical_Operator_out2895_out1;

  Logical_Operator_out4940_out1 <= Logical_Operator_out2888_out1 XOR Logical_Operator_out2896_out1;

  Logical_Operator_out4941_out1 <= Logical_Operator_out1863_out1 XOR Logical_Operator_out1871_out1;

  Logical_Operator_out4942_out1 <= Logical_Operator_out1864_out1 XOR Logical_Operator_out1872_out1;

  Logical_Operator_out4943_out1 <= Logical_Operator_out840_out1 XOR Logical_Operator_out848_out1;

  Logical_Operator_out4944_out1 <= in1680 XOR in1696;

  Logical_Operator_out4945_out1 <= Logical_Operator_out3921_out1 XOR Logical_Operator_out3929_out1;

  Logical_Operator_out4946_out1 <= Logical_Operator_out3922_out1 XOR Logical_Operator_out3930_out1;

  Logical_Operator_out4947_out1 <= Logical_Operator_out3923_out1 XOR Logical_Operator_out3931_out1;

  Logical_Operator_out4948_out1 <= Logical_Operator_out3924_out1 XOR Logical_Operator_out3932_out1;

  Logical_Operator_out4949_out1 <= Logical_Operator_out3925_out1 XOR Logical_Operator_out3933_out1;

  Logical_Operator_out4950_out1 <= Logical_Operator_out3926_out1 XOR Logical_Operator_out3934_out1;

  Logical_Operator_out4951_out1 <= Logical_Operator_out3927_out1 XOR Logical_Operator_out3935_out1;

  Logical_Operator_out4952_out1 <= Logical_Operator_out3928_out1 XOR Logical_Operator_out3936_out1;

  Logical_Operator_out4953_out1 <= Logical_Operator_out2901_out1 XOR Logical_Operator_out2909_out1;

  Logical_Operator_out4954_out1 <= Logical_Operator_out2902_out1 XOR Logical_Operator_out2910_out1;

  Logical_Operator_out4955_out1 <= Logical_Operator_out2903_out1 XOR Logical_Operator_out2911_out1;

  Logical_Operator_out4956_out1 <= Logical_Operator_out2904_out1 XOR Logical_Operator_out2912_out1;

  Logical_Operator_out4957_out1 <= Logical_Operator_out1879_out1 XOR Logical_Operator_out1887_out1;

  Logical_Operator_out4958_out1 <= Logical_Operator_out1880_out1 XOR Logical_Operator_out1888_out1;

  Logical_Operator_out4959_out1 <= Logical_Operator_out856_out1 XOR Logical_Operator_out864_out1;

  Logical_Operator_out4960_out1 <= in1712 XOR in1728;

  Logical_Operator_out4961_out1 <= Logical_Operator_out3937_out1 XOR Logical_Operator_out3945_out1;

  Logical_Operator_out4962_out1 <= Logical_Operator_out3938_out1 XOR Logical_Operator_out3946_out1;

  Logical_Operator_out4963_out1 <= Logical_Operator_out3939_out1 XOR Logical_Operator_out3947_out1;

  Logical_Operator_out4964_out1 <= Logical_Operator_out3940_out1 XOR Logical_Operator_out3948_out1;

  Logical_Operator_out4965_out1 <= Logical_Operator_out3941_out1 XOR Logical_Operator_out3949_out1;

  Logical_Operator_out4966_out1 <= Logical_Operator_out3942_out1 XOR Logical_Operator_out3950_out1;

  Logical_Operator_out4967_out1 <= Logical_Operator_out3943_out1 XOR Logical_Operator_out3951_out1;

  Logical_Operator_out4968_out1 <= Logical_Operator_out3944_out1 XOR Logical_Operator_out3952_out1;

  Logical_Operator_out4969_out1 <= Logical_Operator_out2917_out1 XOR Logical_Operator_out2925_out1;

  Logical_Operator_out4970_out1 <= Logical_Operator_out2918_out1 XOR Logical_Operator_out2926_out1;

  Logical_Operator_out4971_out1 <= Logical_Operator_out2919_out1 XOR Logical_Operator_out2927_out1;

  Logical_Operator_out4972_out1 <= Logical_Operator_out2920_out1 XOR Logical_Operator_out2928_out1;

  Logical_Operator_out4973_out1 <= Logical_Operator_out1895_out1 XOR Logical_Operator_out1903_out1;

  Logical_Operator_out4974_out1 <= Logical_Operator_out1896_out1 XOR Logical_Operator_out1904_out1;

  Logical_Operator_out4975_out1 <= Logical_Operator_out872_out1 XOR Logical_Operator_out880_out1;

  Logical_Operator_out4976_out1 <= in1744 XOR in1760;

  Logical_Operator_out4977_out1 <= Logical_Operator_out3953_out1 XOR Logical_Operator_out3961_out1;

  Logical_Operator_out4978_out1 <= Logical_Operator_out3954_out1 XOR Logical_Operator_out3962_out1;

  Logical_Operator_out4979_out1 <= Logical_Operator_out3955_out1 XOR Logical_Operator_out3963_out1;

  Logical_Operator_out4980_out1 <= Logical_Operator_out3956_out1 XOR Logical_Operator_out3964_out1;

  Logical_Operator_out4981_out1 <= Logical_Operator_out3957_out1 XOR Logical_Operator_out3965_out1;

  Logical_Operator_out4982_out1 <= Logical_Operator_out3958_out1 XOR Logical_Operator_out3966_out1;

  Logical_Operator_out4983_out1 <= Logical_Operator_out3959_out1 XOR Logical_Operator_out3967_out1;

  Logical_Operator_out4984_out1 <= Logical_Operator_out3960_out1 XOR Logical_Operator_out3968_out1;

  Logical_Operator_out4985_out1 <= Logical_Operator_out2933_out1 XOR Logical_Operator_out2941_out1;

  Logical_Operator_out4986_out1 <= Logical_Operator_out2934_out1 XOR Logical_Operator_out2942_out1;

  Logical_Operator_out4987_out1 <= Logical_Operator_out2935_out1 XOR Logical_Operator_out2943_out1;

  Logical_Operator_out4988_out1 <= Logical_Operator_out2936_out1 XOR Logical_Operator_out2944_out1;

  Logical_Operator_out4989_out1 <= Logical_Operator_out1911_out1 XOR Logical_Operator_out1919_out1;

  Logical_Operator_out4990_out1 <= Logical_Operator_out1912_out1 XOR Logical_Operator_out1920_out1;

  Logical_Operator_out4991_out1 <= Logical_Operator_out888_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out4992_out1 <= in1776 XOR in1792;

  Logical_Operator_out4993_out1 <= Logical_Operator_out3969_out1 XOR Logical_Operator_out3977_out1;

  Logical_Operator_out4994_out1 <= Logical_Operator_out3970_out1 XOR Logical_Operator_out3978_out1;

  Logical_Operator_out4995_out1 <= Logical_Operator_out3971_out1 XOR Logical_Operator_out3979_out1;

  Logical_Operator_out4996_out1 <= Logical_Operator_out3972_out1 XOR Logical_Operator_out3980_out1;

  Logical_Operator_out4997_out1 <= Logical_Operator_out3973_out1 XOR Logical_Operator_out3981_out1;

  Logical_Operator_out4998_out1 <= Logical_Operator_out3974_out1 XOR Logical_Operator_out3982_out1;

  Logical_Operator_out4999_out1 <= Logical_Operator_out3975_out1 XOR Logical_Operator_out3983_out1;

  Logical_Operator_out5000_out1 <= Logical_Operator_out3976_out1 XOR Logical_Operator_out3984_out1;

  Logical_Operator_out5001_out1 <= Logical_Operator_out2949_out1 XOR Logical_Operator_out2957_out1;

  Logical_Operator_out5002_out1 <= Logical_Operator_out2950_out1 XOR Logical_Operator_out2958_out1;

  Logical_Operator_out5003_out1 <= Logical_Operator_out2951_out1 XOR Logical_Operator_out2959_out1;

  Logical_Operator_out5004_out1 <= Logical_Operator_out2952_out1 XOR Logical_Operator_out2960_out1;

  Logical_Operator_out5005_out1 <= Logical_Operator_out1927_out1 XOR Logical_Operator_out1935_out1;

  Logical_Operator_out5006_out1 <= Logical_Operator_out1928_out1 XOR Logical_Operator_out1936_out1;

  Logical_Operator_out5007_out1 <= Logical_Operator_out904_out1 XOR Logical_Operator_out912_out1;

  Logical_Operator_out5008_out1 <= in1808 XOR in1824;

  Logical_Operator_out5009_out1 <= Logical_Operator_out3985_out1 XOR Logical_Operator_out3993_out1;

  Logical_Operator_out5010_out1 <= Logical_Operator_out3986_out1 XOR Logical_Operator_out3994_out1;

  Logical_Operator_out5011_out1 <= Logical_Operator_out3987_out1 XOR Logical_Operator_out3995_out1;

  Logical_Operator_out5012_out1 <= Logical_Operator_out3988_out1 XOR Logical_Operator_out3996_out1;

  Logical_Operator_out5013_out1 <= Logical_Operator_out3989_out1 XOR Logical_Operator_out3997_out1;

  Logical_Operator_out5014_out1 <= Logical_Operator_out3990_out1 XOR Logical_Operator_out3998_out1;

  Logical_Operator_out5015_out1 <= Logical_Operator_out3991_out1 XOR Logical_Operator_out3999_out1;

  Logical_Operator_out5016_out1 <= Logical_Operator_out3992_out1 XOR Logical_Operator_out4000_out1;

  Logical_Operator_out5017_out1 <= Logical_Operator_out2965_out1 XOR Logical_Operator_out2973_out1;

  Logical_Operator_out5018_out1 <= Logical_Operator_out2966_out1 XOR Logical_Operator_out2974_out1;

  Logical_Operator_out5019_out1 <= Logical_Operator_out2967_out1 XOR Logical_Operator_out2975_out1;

  Logical_Operator_out5020_out1 <= Logical_Operator_out2968_out1 XOR Logical_Operator_out2976_out1;

  Logical_Operator_out5021_out1 <= Logical_Operator_out1943_out1 XOR Logical_Operator_out1951_out1;

  Logical_Operator_out5022_out1 <= Logical_Operator_out1944_out1 XOR Logical_Operator_out1952_out1;

  Logical_Operator_out5023_out1 <= Logical_Operator_out920_out1 XOR Logical_Operator_out928_out1;

  Logical_Operator_out5024_out1 <= in1840 XOR in1856;

  Logical_Operator_out5025_out1 <= Logical_Operator_out4001_out1 XOR Logical_Operator_out4009_out1;

  Logical_Operator_out5026_out1 <= Logical_Operator_out4002_out1 XOR Logical_Operator_out4010_out1;

  Logical_Operator_out5027_out1 <= Logical_Operator_out4003_out1 XOR Logical_Operator_out4011_out1;

  Logical_Operator_out5028_out1 <= Logical_Operator_out4004_out1 XOR Logical_Operator_out4012_out1;

  Logical_Operator_out5029_out1 <= Logical_Operator_out4005_out1 XOR Logical_Operator_out4013_out1;

  Logical_Operator_out5030_out1 <= Logical_Operator_out4006_out1 XOR Logical_Operator_out4014_out1;

  Logical_Operator_out5031_out1 <= Logical_Operator_out4007_out1 XOR Logical_Operator_out4015_out1;

  Logical_Operator_out5032_out1 <= Logical_Operator_out4008_out1 XOR Logical_Operator_out4016_out1;

  Logical_Operator_out5033_out1 <= Logical_Operator_out2981_out1 XOR Logical_Operator_out2989_out1;

  Logical_Operator_out5034_out1 <= Logical_Operator_out2982_out1 XOR Logical_Operator_out2990_out1;

  Logical_Operator_out5035_out1 <= Logical_Operator_out2983_out1 XOR Logical_Operator_out2991_out1;

  Logical_Operator_out5036_out1 <= Logical_Operator_out2984_out1 XOR Logical_Operator_out2992_out1;

  Logical_Operator_out5037_out1 <= Logical_Operator_out1959_out1 XOR Logical_Operator_out1967_out1;

  Logical_Operator_out5038_out1 <= Logical_Operator_out1960_out1 XOR Logical_Operator_out1968_out1;

  Logical_Operator_out5039_out1 <= Logical_Operator_out936_out1 XOR Logical_Operator_out944_out1;

  Logical_Operator_out5040_out1 <= in1872 XOR in1888;

  Logical_Operator_out5041_out1 <= Logical_Operator_out4017_out1 XOR Logical_Operator_out4025_out1;

  Logical_Operator_out5042_out1 <= Logical_Operator_out4018_out1 XOR Logical_Operator_out4026_out1;

  Logical_Operator_out5043_out1 <= Logical_Operator_out4019_out1 XOR Logical_Operator_out4027_out1;

  Logical_Operator_out5044_out1 <= Logical_Operator_out4020_out1 XOR Logical_Operator_out4028_out1;

  Logical_Operator_out5045_out1 <= Logical_Operator_out4021_out1 XOR Logical_Operator_out4029_out1;

  Logical_Operator_out5046_out1 <= Logical_Operator_out4022_out1 XOR Logical_Operator_out4030_out1;

  Logical_Operator_out5047_out1 <= Logical_Operator_out4023_out1 XOR Logical_Operator_out4031_out1;

  Logical_Operator_out5048_out1 <= Logical_Operator_out4024_out1 XOR Logical_Operator_out4032_out1;

  Logical_Operator_out5049_out1 <= Logical_Operator_out2997_out1 XOR Logical_Operator_out3005_out1;

  Logical_Operator_out5050_out1 <= Logical_Operator_out2998_out1 XOR Logical_Operator_out3006_out1;

  Logical_Operator_out5051_out1 <= Logical_Operator_out2999_out1 XOR Logical_Operator_out3007_out1;

  Logical_Operator_out5052_out1 <= Logical_Operator_out3000_out1 XOR Logical_Operator_out3008_out1;

  Logical_Operator_out5053_out1 <= Logical_Operator_out1975_out1 XOR Logical_Operator_out1983_out1;

  Logical_Operator_out5054_out1 <= Logical_Operator_out1976_out1 XOR Logical_Operator_out1984_out1;

  Logical_Operator_out5055_out1 <= Logical_Operator_out952_out1 XOR Logical_Operator_out960_out1;

  Logical_Operator_out5056_out1 <= in1904 XOR in1920;

  Logical_Operator_out5057_out1 <= Logical_Operator_out4033_out1 XOR Logical_Operator_out4041_out1;

  Logical_Operator_out5058_out1 <= Logical_Operator_out4034_out1 XOR Logical_Operator_out4042_out1;

  Logical_Operator_out5059_out1 <= Logical_Operator_out4035_out1 XOR Logical_Operator_out4043_out1;

  Logical_Operator_out5060_out1 <= Logical_Operator_out4036_out1 XOR Logical_Operator_out4044_out1;

  Logical_Operator_out5061_out1 <= Logical_Operator_out4037_out1 XOR Logical_Operator_out4045_out1;

  Logical_Operator_out5062_out1 <= Logical_Operator_out4038_out1 XOR Logical_Operator_out4046_out1;

  Logical_Operator_out5063_out1 <= Logical_Operator_out4039_out1 XOR Logical_Operator_out4047_out1;

  Logical_Operator_out5064_out1 <= Logical_Operator_out4040_out1 XOR Logical_Operator_out4048_out1;

  Logical_Operator_out5065_out1 <= Logical_Operator_out3013_out1 XOR Logical_Operator_out3021_out1;

  Logical_Operator_out5066_out1 <= Logical_Operator_out3014_out1 XOR Logical_Operator_out3022_out1;

  Logical_Operator_out5067_out1 <= Logical_Operator_out3015_out1 XOR Logical_Operator_out3023_out1;

  Logical_Operator_out5068_out1 <= Logical_Operator_out3016_out1 XOR Logical_Operator_out3024_out1;

  Logical_Operator_out5069_out1 <= Logical_Operator_out1991_out1 XOR Logical_Operator_out1999_out1;

  Logical_Operator_out5070_out1 <= Logical_Operator_out1992_out1 XOR Logical_Operator_out2000_out1;

  Logical_Operator_out5071_out1 <= Logical_Operator_out968_out1 XOR Logical_Operator_out976_out1;

  Logical_Operator_out5072_out1 <= in1936 XOR in1952;

  Logical_Operator_out5073_out1 <= Logical_Operator_out4049_out1 XOR Logical_Operator_out4057_out1;

  Logical_Operator_out5074_out1 <= Logical_Operator_out4050_out1 XOR Logical_Operator_out4058_out1;

  Logical_Operator_out5075_out1 <= Logical_Operator_out4051_out1 XOR Logical_Operator_out4059_out1;

  Logical_Operator_out5076_out1 <= Logical_Operator_out4052_out1 XOR Logical_Operator_out4060_out1;

  Logical_Operator_out5077_out1 <= Logical_Operator_out4053_out1 XOR Logical_Operator_out4061_out1;

  Logical_Operator_out5078_out1 <= Logical_Operator_out4054_out1 XOR Logical_Operator_out4062_out1;

  Logical_Operator_out5079_out1 <= Logical_Operator_out4055_out1 XOR Logical_Operator_out4063_out1;

  Logical_Operator_out5080_out1 <= Logical_Operator_out4056_out1 XOR Logical_Operator_out4064_out1;

  Logical_Operator_out5081_out1 <= Logical_Operator_out3029_out1 XOR Logical_Operator_out3037_out1;

  Logical_Operator_out5082_out1 <= Logical_Operator_out3030_out1 XOR Logical_Operator_out3038_out1;

  Logical_Operator_out5083_out1 <= Logical_Operator_out3031_out1 XOR Logical_Operator_out3039_out1;

  Logical_Operator_out5084_out1 <= Logical_Operator_out3032_out1 XOR Logical_Operator_out3040_out1;

  Logical_Operator_out5085_out1 <= Logical_Operator_out2007_out1 XOR Logical_Operator_out2015_out1;

  Logical_Operator_out5086_out1 <= Logical_Operator_out2008_out1 XOR Logical_Operator_out2016_out1;

  Logical_Operator_out5087_out1 <= Logical_Operator_out984_out1 XOR Logical_Operator_out992_out1;

  Logical_Operator_out5088_out1 <= in1968 XOR in1984;

  Logical_Operator_out5089_out1 <= Logical_Operator_out4065_out1 XOR Logical_Operator_out4073_out1;

  Logical_Operator_out5090_out1 <= Logical_Operator_out4066_out1 XOR Logical_Operator_out4074_out1;

  Logical_Operator_out5091_out1 <= Logical_Operator_out4067_out1 XOR Logical_Operator_out4075_out1;

  Logical_Operator_out5092_out1 <= Logical_Operator_out4068_out1 XOR Logical_Operator_out4076_out1;

  Logical_Operator_out5093_out1 <= Logical_Operator_out4069_out1 XOR Logical_Operator_out4077_out1;

  Logical_Operator_out5094_out1 <= Logical_Operator_out4070_out1 XOR Logical_Operator_out4078_out1;

  Logical_Operator_out5095_out1 <= Logical_Operator_out4071_out1 XOR Logical_Operator_out4079_out1;

  Logical_Operator_out5096_out1 <= Logical_Operator_out4072_out1 XOR Logical_Operator_out4080_out1;

  Logical_Operator_out5097_out1 <= Logical_Operator_out3045_out1 XOR Logical_Operator_out3053_out1;

  Logical_Operator_out5098_out1 <= Logical_Operator_out3046_out1 XOR Logical_Operator_out3054_out1;

  Logical_Operator_out5099_out1 <= Logical_Operator_out3047_out1 XOR Logical_Operator_out3055_out1;

  Logical_Operator_out5100_out1 <= Logical_Operator_out3048_out1 XOR Logical_Operator_out3056_out1;

  Logical_Operator_out5101_out1 <= Logical_Operator_out2023_out1 XOR Logical_Operator_out2031_out1;

  Logical_Operator_out5102_out1 <= Logical_Operator_out2024_out1 XOR Logical_Operator_out2032_out1;

  Logical_Operator_out5103_out1 <= Logical_Operator_out1000_out1 XOR Logical_Operator_out1008_out1;

  Logical_Operator_out5104_out1 <= in2000 XOR in2016;

  Logical_Operator_out5105_out1 <= Logical_Operator_out4081_out1 XOR Logical_Operator_out4089_out1;

  Logical_Operator_out5106_out1 <= Logical_Operator_out4082_out1 XOR Logical_Operator_out4090_out1;

  Logical_Operator_out5107_out1 <= Logical_Operator_out4083_out1 XOR Logical_Operator_out4091_out1;

  Logical_Operator_out5108_out1 <= Logical_Operator_out4084_out1 XOR Logical_Operator_out4092_out1;

  Logical_Operator_out5109_out1 <= Logical_Operator_out4085_out1 XOR Logical_Operator_out4093_out1;

  Logical_Operator_out5110_out1 <= Logical_Operator_out4086_out1 XOR Logical_Operator_out4094_out1;

  Logical_Operator_out5111_out1 <= Logical_Operator_out4087_out1 XOR Logical_Operator_out4095_out1;

  Logical_Operator_out5112_out1 <= Logical_Operator_out4088_out1 XOR Logical_Operator_out4096_out1;

  Logical_Operator_out5113_out1 <= Logical_Operator_out3061_out1 XOR Logical_Operator_out3069_out1;

  Logical_Operator_out5114_out1 <= Logical_Operator_out3062_out1 XOR Logical_Operator_out3070_out1;

  Logical_Operator_out5115_out1 <= Logical_Operator_out3063_out1 XOR Logical_Operator_out3071_out1;

  Logical_Operator_out5116_out1 <= Logical_Operator_out3064_out1 XOR Logical_Operator_out3072_out1;

  Logical_Operator_out5117_out1 <= Logical_Operator_out2039_out1 XOR Logical_Operator_out2047_out1;

  Logical_Operator_out5118_out1 <= Logical_Operator_out2040_out1 XOR Logical_Operator_out2048_out1;

  Logical_Operator_out5119_out1 <= Logical_Operator_out1016_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out5120_out1 <= in2032 XOR in2048;

  Logical_Operator_out5121_out1 <= Logical_Operator_out4097_out1 XOR Logical_Operator_out4113_out1;

  Logical_Operator_out5122_out1 <= Logical_Operator_out4098_out1 XOR Logical_Operator_out4114_out1;

  Logical_Operator_out5123_out1 <= Logical_Operator_out4099_out1 XOR Logical_Operator_out4115_out1;

  Logical_Operator_out5124_out1 <= Logical_Operator_out4100_out1 XOR Logical_Operator_out4116_out1;

  Logical_Operator_out5125_out1 <= Logical_Operator_out4101_out1 XOR Logical_Operator_out4117_out1;

  Logical_Operator_out5126_out1 <= Logical_Operator_out4102_out1 XOR Logical_Operator_out4118_out1;

  Logical_Operator_out5127_out1 <= Logical_Operator_out4103_out1 XOR Logical_Operator_out4119_out1;

  Logical_Operator_out5128_out1 <= Logical_Operator_out4104_out1 XOR Logical_Operator_out4120_out1;

  Logical_Operator_out5129_out1 <= Logical_Operator_out4105_out1 XOR Logical_Operator_out4121_out1;

  Logical_Operator_out5130_out1 <= Logical_Operator_out4106_out1 XOR Logical_Operator_out4122_out1;

  Logical_Operator_out5131_out1 <= Logical_Operator_out4107_out1 XOR Logical_Operator_out4123_out1;

  Logical_Operator_out5132_out1 <= Logical_Operator_out4108_out1 XOR Logical_Operator_out4124_out1;

  Logical_Operator_out5133_out1 <= Logical_Operator_out4109_out1 XOR Logical_Operator_out4125_out1;

  Logical_Operator_out5134_out1 <= Logical_Operator_out4110_out1 XOR Logical_Operator_out4126_out1;

  Logical_Operator_out5135_out1 <= Logical_Operator_out4111_out1 XOR Logical_Operator_out4127_out1;

  Logical_Operator_out5136_out1 <= Logical_Operator_out4112_out1 XOR Logical_Operator_out4128_out1;

  Logical_Operator_out5137_out1 <= Logical_Operator_out3081_out1 XOR Logical_Operator_out3097_out1;

  Logical_Operator_out5138_out1 <= Logical_Operator_out3082_out1 XOR Logical_Operator_out3098_out1;

  Logical_Operator_out5139_out1 <= Logical_Operator_out3083_out1 XOR Logical_Operator_out3099_out1;

  Logical_Operator_out5140_out1 <= Logical_Operator_out3084_out1 XOR Logical_Operator_out3100_out1;

  Logical_Operator_out5141_out1 <= Logical_Operator_out3085_out1 XOR Logical_Operator_out3101_out1;

  Logical_Operator_out5142_out1 <= Logical_Operator_out3086_out1 XOR Logical_Operator_out3102_out1;

  Logical_Operator_out5143_out1 <= Logical_Operator_out3087_out1 XOR Logical_Operator_out3103_out1;

  Logical_Operator_out5144_out1 <= Logical_Operator_out3088_out1 XOR Logical_Operator_out3104_out1;

  Logical_Operator_out5145_out1 <= Logical_Operator_out2061_out1 XOR Logical_Operator_out2077_out1;

  Logical_Operator_out5146_out1 <= Logical_Operator_out2062_out1 XOR Logical_Operator_out2078_out1;

  Logical_Operator_out5147_out1 <= Logical_Operator_out2063_out1 XOR Logical_Operator_out2079_out1;

  Logical_Operator_out5148_out1 <= Logical_Operator_out2064_out1 XOR Logical_Operator_out2080_out1;

  Logical_Operator_out5149_out1 <= Logical_Operator_out1039_out1 XOR Logical_Operator_out1055_out1;

  Logical_Operator_out5150_out1 <= Logical_Operator_out1040_out1 XOR Logical_Operator_out1056_out1;

  Logical_Operator_out5151_out1 <= Logical_Operator_out16_out1 XOR Logical_Operator_out32_out1;

  Logical_Operator_out5152_out1 <= in32 XOR in64;

  Logical_Operator_out5153_out1 <= Logical_Operator_out4129_out1 XOR Logical_Operator_out4145_out1;

  Logical_Operator_out5154_out1 <= Logical_Operator_out4130_out1 XOR Logical_Operator_out4146_out1;

  Logical_Operator_out5155_out1 <= Logical_Operator_out4131_out1 XOR Logical_Operator_out4147_out1;

  Logical_Operator_out5156_out1 <= Logical_Operator_out4132_out1 XOR Logical_Operator_out4148_out1;

  Logical_Operator_out5157_out1 <= Logical_Operator_out4133_out1 XOR Logical_Operator_out4149_out1;

  Logical_Operator_out5158_out1 <= Logical_Operator_out4134_out1 XOR Logical_Operator_out4150_out1;

  Logical_Operator_out5159_out1 <= Logical_Operator_out4135_out1 XOR Logical_Operator_out4151_out1;

  Logical_Operator_out5160_out1 <= Logical_Operator_out4136_out1 XOR Logical_Operator_out4152_out1;

  Logical_Operator_out5161_out1 <= Logical_Operator_out4137_out1 XOR Logical_Operator_out4153_out1;

  Logical_Operator_out5162_out1 <= Logical_Operator_out4138_out1 XOR Logical_Operator_out4154_out1;

  Logical_Operator_out5163_out1 <= Logical_Operator_out4139_out1 XOR Logical_Operator_out4155_out1;

  Logical_Operator_out5164_out1 <= Logical_Operator_out4140_out1 XOR Logical_Operator_out4156_out1;

  Logical_Operator_out5165_out1 <= Logical_Operator_out4141_out1 XOR Logical_Operator_out4157_out1;

  Logical_Operator_out5166_out1 <= Logical_Operator_out4142_out1 XOR Logical_Operator_out4158_out1;

  Logical_Operator_out5167_out1 <= Logical_Operator_out4143_out1 XOR Logical_Operator_out4159_out1;

  Logical_Operator_out5168_out1 <= Logical_Operator_out4144_out1 XOR Logical_Operator_out4160_out1;

  Logical_Operator_out5169_out1 <= Logical_Operator_out3113_out1 XOR Logical_Operator_out3129_out1;

  Logical_Operator_out5170_out1 <= Logical_Operator_out3114_out1 XOR Logical_Operator_out3130_out1;

  Logical_Operator_out5171_out1 <= Logical_Operator_out3115_out1 XOR Logical_Operator_out3131_out1;

  Logical_Operator_out5172_out1 <= Logical_Operator_out3116_out1 XOR Logical_Operator_out3132_out1;

  Logical_Operator_out5173_out1 <= Logical_Operator_out3117_out1 XOR Logical_Operator_out3133_out1;

  Logical_Operator_out5174_out1 <= Logical_Operator_out3118_out1 XOR Logical_Operator_out3134_out1;

  Logical_Operator_out5175_out1 <= Logical_Operator_out3119_out1 XOR Logical_Operator_out3135_out1;

  Logical_Operator_out5176_out1 <= Logical_Operator_out3120_out1 XOR Logical_Operator_out3136_out1;

  Logical_Operator_out5177_out1 <= Logical_Operator_out2093_out1 XOR Logical_Operator_out2109_out1;

  Logical_Operator_out5178_out1 <= Logical_Operator_out2094_out1 XOR Logical_Operator_out2110_out1;

  Logical_Operator_out5179_out1 <= Logical_Operator_out2095_out1 XOR Logical_Operator_out2111_out1;

  Logical_Operator_out5180_out1 <= Logical_Operator_out2096_out1 XOR Logical_Operator_out2112_out1;

  Logical_Operator_out5181_out1 <= Logical_Operator_out1071_out1 XOR Logical_Operator_out1087_out1;

  Logical_Operator_out5182_out1 <= Logical_Operator_out1072_out1 XOR Logical_Operator_out1088_out1;

  Logical_Operator_out5183_out1 <= Logical_Operator_out48_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out5184_out1 <= in96 XOR in128;

  Logical_Operator_out5185_out1 <= Logical_Operator_out4161_out1 XOR Logical_Operator_out4177_out1;

  Logical_Operator_out5186_out1 <= Logical_Operator_out4162_out1 XOR Logical_Operator_out4178_out1;

  Logical_Operator_out5187_out1 <= Logical_Operator_out4163_out1 XOR Logical_Operator_out4179_out1;

  Logical_Operator_out5188_out1 <= Logical_Operator_out4164_out1 XOR Logical_Operator_out4180_out1;

  Logical_Operator_out5189_out1 <= Logical_Operator_out4165_out1 XOR Logical_Operator_out4181_out1;

  Logical_Operator_out5190_out1 <= Logical_Operator_out4166_out1 XOR Logical_Operator_out4182_out1;

  Logical_Operator_out5191_out1 <= Logical_Operator_out4167_out1 XOR Logical_Operator_out4183_out1;

  Logical_Operator_out5192_out1 <= Logical_Operator_out4168_out1 XOR Logical_Operator_out4184_out1;

  Logical_Operator_out5193_out1 <= Logical_Operator_out4169_out1 XOR Logical_Operator_out4185_out1;

  Logical_Operator_out5194_out1 <= Logical_Operator_out4170_out1 XOR Logical_Operator_out4186_out1;

  Logical_Operator_out5195_out1 <= Logical_Operator_out4171_out1 XOR Logical_Operator_out4187_out1;

  Logical_Operator_out5196_out1 <= Logical_Operator_out4172_out1 XOR Logical_Operator_out4188_out1;

  Logical_Operator_out5197_out1 <= Logical_Operator_out4173_out1 XOR Logical_Operator_out4189_out1;

  Logical_Operator_out5198_out1 <= Logical_Operator_out4174_out1 XOR Logical_Operator_out4190_out1;

  Logical_Operator_out5199_out1 <= Logical_Operator_out4175_out1 XOR Logical_Operator_out4191_out1;

  Logical_Operator_out5200_out1 <= Logical_Operator_out4176_out1 XOR Logical_Operator_out4192_out1;

  Logical_Operator_out5201_out1 <= Logical_Operator_out3145_out1 XOR Logical_Operator_out3161_out1;

  Logical_Operator_out5202_out1 <= Logical_Operator_out3146_out1 XOR Logical_Operator_out3162_out1;

  Logical_Operator_out5203_out1 <= Logical_Operator_out3147_out1 XOR Logical_Operator_out3163_out1;

  Logical_Operator_out5204_out1 <= Logical_Operator_out3148_out1 XOR Logical_Operator_out3164_out1;

  Logical_Operator_out5205_out1 <= Logical_Operator_out3149_out1 XOR Logical_Operator_out3165_out1;

  Logical_Operator_out5206_out1 <= Logical_Operator_out3150_out1 XOR Logical_Operator_out3166_out1;

  Logical_Operator_out5207_out1 <= Logical_Operator_out3151_out1 XOR Logical_Operator_out3167_out1;

  Logical_Operator_out5208_out1 <= Logical_Operator_out3152_out1 XOR Logical_Operator_out3168_out1;

  Logical_Operator_out5209_out1 <= Logical_Operator_out2125_out1 XOR Logical_Operator_out2141_out1;

  Logical_Operator_out5210_out1 <= Logical_Operator_out2126_out1 XOR Logical_Operator_out2142_out1;

  Logical_Operator_out5211_out1 <= Logical_Operator_out2127_out1 XOR Logical_Operator_out2143_out1;

  Logical_Operator_out5212_out1 <= Logical_Operator_out2128_out1 XOR Logical_Operator_out2144_out1;

  Logical_Operator_out5213_out1 <= Logical_Operator_out1103_out1 XOR Logical_Operator_out1119_out1;

  Logical_Operator_out5214_out1 <= Logical_Operator_out1104_out1 XOR Logical_Operator_out1120_out1;

  Logical_Operator_out5215_out1 <= Logical_Operator_out80_out1 XOR Logical_Operator_out96_out1;

  Logical_Operator_out5216_out1 <= in160 XOR in192;

  Logical_Operator_out5217_out1 <= Logical_Operator_out4193_out1 XOR Logical_Operator_out4209_out1;

  Logical_Operator_out5218_out1 <= Logical_Operator_out4194_out1 XOR Logical_Operator_out4210_out1;

  Logical_Operator_out5219_out1 <= Logical_Operator_out4195_out1 XOR Logical_Operator_out4211_out1;

  Logical_Operator_out5220_out1 <= Logical_Operator_out4196_out1 XOR Logical_Operator_out4212_out1;

  Logical_Operator_out5221_out1 <= Logical_Operator_out4197_out1 XOR Logical_Operator_out4213_out1;

  Logical_Operator_out5222_out1 <= Logical_Operator_out4198_out1 XOR Logical_Operator_out4214_out1;

  Logical_Operator_out5223_out1 <= Logical_Operator_out4199_out1 XOR Logical_Operator_out4215_out1;

  Logical_Operator_out5224_out1 <= Logical_Operator_out4200_out1 XOR Logical_Operator_out4216_out1;

  Logical_Operator_out5225_out1 <= Logical_Operator_out4201_out1 XOR Logical_Operator_out4217_out1;

  Logical_Operator_out5226_out1 <= Logical_Operator_out4202_out1 XOR Logical_Operator_out4218_out1;

  Logical_Operator_out5227_out1 <= Logical_Operator_out4203_out1 XOR Logical_Operator_out4219_out1;

  Logical_Operator_out5228_out1 <= Logical_Operator_out4204_out1 XOR Logical_Operator_out4220_out1;

  Logical_Operator_out5229_out1 <= Logical_Operator_out4205_out1 XOR Logical_Operator_out4221_out1;

  Logical_Operator_out5230_out1 <= Logical_Operator_out4206_out1 XOR Logical_Operator_out4222_out1;

  Logical_Operator_out5231_out1 <= Logical_Operator_out4207_out1 XOR Logical_Operator_out4223_out1;

  Logical_Operator_out5232_out1 <= Logical_Operator_out4208_out1 XOR Logical_Operator_out4224_out1;

  Logical_Operator_out5233_out1 <= Logical_Operator_out3177_out1 XOR Logical_Operator_out3193_out1;

  Logical_Operator_out5234_out1 <= Logical_Operator_out3178_out1 XOR Logical_Operator_out3194_out1;

  Logical_Operator_out5235_out1 <= Logical_Operator_out3179_out1 XOR Logical_Operator_out3195_out1;

  Logical_Operator_out5236_out1 <= Logical_Operator_out3180_out1 XOR Logical_Operator_out3196_out1;

  Logical_Operator_out5237_out1 <= Logical_Operator_out3181_out1 XOR Logical_Operator_out3197_out1;

  Logical_Operator_out5238_out1 <= Logical_Operator_out3182_out1 XOR Logical_Operator_out3198_out1;

  Logical_Operator_out5239_out1 <= Logical_Operator_out3183_out1 XOR Logical_Operator_out3199_out1;

  Logical_Operator_out5240_out1 <= Logical_Operator_out3184_out1 XOR Logical_Operator_out3200_out1;

  Logical_Operator_out5241_out1 <= Logical_Operator_out2157_out1 XOR Logical_Operator_out2173_out1;

  Logical_Operator_out5242_out1 <= Logical_Operator_out2158_out1 XOR Logical_Operator_out2174_out1;

  Logical_Operator_out5243_out1 <= Logical_Operator_out2159_out1 XOR Logical_Operator_out2175_out1;

  Logical_Operator_out5244_out1 <= Logical_Operator_out2160_out1 XOR Logical_Operator_out2176_out1;

  Logical_Operator_out5245_out1 <= Logical_Operator_out1135_out1 XOR Logical_Operator_out1151_out1;

  Logical_Operator_out5246_out1 <= Logical_Operator_out1136_out1 XOR Logical_Operator_out1152_out1;

  Logical_Operator_out5247_out1 <= Logical_Operator_out112_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out5248_out1 <= in224 XOR in256;

  Logical_Operator_out5249_out1 <= Logical_Operator_out4225_out1 XOR Logical_Operator_out4241_out1;

  Logical_Operator_out5250_out1 <= Logical_Operator_out4226_out1 XOR Logical_Operator_out4242_out1;

  Logical_Operator_out5251_out1 <= Logical_Operator_out4227_out1 XOR Logical_Operator_out4243_out1;

  Logical_Operator_out5252_out1 <= Logical_Operator_out4228_out1 XOR Logical_Operator_out4244_out1;

  Logical_Operator_out5253_out1 <= Logical_Operator_out4229_out1 XOR Logical_Operator_out4245_out1;

  Logical_Operator_out5254_out1 <= Logical_Operator_out4230_out1 XOR Logical_Operator_out4246_out1;

  Logical_Operator_out5255_out1 <= Logical_Operator_out4231_out1 XOR Logical_Operator_out4247_out1;

  Logical_Operator_out5256_out1 <= Logical_Operator_out4232_out1 XOR Logical_Operator_out4248_out1;

  Logical_Operator_out5257_out1 <= Logical_Operator_out4233_out1 XOR Logical_Operator_out4249_out1;

  Logical_Operator_out5258_out1 <= Logical_Operator_out4234_out1 XOR Logical_Operator_out4250_out1;

  Logical_Operator_out5259_out1 <= Logical_Operator_out4235_out1 XOR Logical_Operator_out4251_out1;

  Logical_Operator_out5260_out1 <= Logical_Operator_out4236_out1 XOR Logical_Operator_out4252_out1;

  Logical_Operator_out5261_out1 <= Logical_Operator_out4237_out1 XOR Logical_Operator_out4253_out1;

  Logical_Operator_out5262_out1 <= Logical_Operator_out4238_out1 XOR Logical_Operator_out4254_out1;

  Logical_Operator_out5263_out1 <= Logical_Operator_out4239_out1 XOR Logical_Operator_out4255_out1;

  Logical_Operator_out5264_out1 <= Logical_Operator_out4240_out1 XOR Logical_Operator_out4256_out1;

  Logical_Operator_out5265_out1 <= Logical_Operator_out3209_out1 XOR Logical_Operator_out3225_out1;

  Logical_Operator_out5266_out1 <= Logical_Operator_out3210_out1 XOR Logical_Operator_out3226_out1;

  Logical_Operator_out5267_out1 <= Logical_Operator_out3211_out1 XOR Logical_Operator_out3227_out1;

  Logical_Operator_out5268_out1 <= Logical_Operator_out3212_out1 XOR Logical_Operator_out3228_out1;

  Logical_Operator_out5269_out1 <= Logical_Operator_out3213_out1 XOR Logical_Operator_out3229_out1;

  Logical_Operator_out5270_out1 <= Logical_Operator_out3214_out1 XOR Logical_Operator_out3230_out1;

  Logical_Operator_out5271_out1 <= Logical_Operator_out3215_out1 XOR Logical_Operator_out3231_out1;

  Logical_Operator_out5272_out1 <= Logical_Operator_out3216_out1 XOR Logical_Operator_out3232_out1;

  Logical_Operator_out5273_out1 <= Logical_Operator_out2189_out1 XOR Logical_Operator_out2205_out1;

  Logical_Operator_out5274_out1 <= Logical_Operator_out2190_out1 XOR Logical_Operator_out2206_out1;

  Logical_Operator_out5275_out1 <= Logical_Operator_out2191_out1 XOR Logical_Operator_out2207_out1;

  Logical_Operator_out5276_out1 <= Logical_Operator_out2192_out1 XOR Logical_Operator_out2208_out1;

  Logical_Operator_out5277_out1 <= Logical_Operator_out1167_out1 XOR Logical_Operator_out1183_out1;

  Logical_Operator_out5278_out1 <= Logical_Operator_out1168_out1 XOR Logical_Operator_out1184_out1;

  Logical_Operator_out5279_out1 <= Logical_Operator_out144_out1 XOR Logical_Operator_out160_out1;

  Logical_Operator_out5280_out1 <= in288 XOR in320;

  Logical_Operator_out5281_out1 <= Logical_Operator_out4257_out1 XOR Logical_Operator_out4273_out1;

  Logical_Operator_out5282_out1 <= Logical_Operator_out4258_out1 XOR Logical_Operator_out4274_out1;

  Logical_Operator_out5283_out1 <= Logical_Operator_out4259_out1 XOR Logical_Operator_out4275_out1;

  Logical_Operator_out5284_out1 <= Logical_Operator_out4260_out1 XOR Logical_Operator_out4276_out1;

  Logical_Operator_out5285_out1 <= Logical_Operator_out4261_out1 XOR Logical_Operator_out4277_out1;

  Logical_Operator_out5286_out1 <= Logical_Operator_out4262_out1 XOR Logical_Operator_out4278_out1;

  Logical_Operator_out5287_out1 <= Logical_Operator_out4263_out1 XOR Logical_Operator_out4279_out1;

  Logical_Operator_out5288_out1 <= Logical_Operator_out4264_out1 XOR Logical_Operator_out4280_out1;

  Logical_Operator_out5289_out1 <= Logical_Operator_out4265_out1 XOR Logical_Operator_out4281_out1;

  Logical_Operator_out5290_out1 <= Logical_Operator_out4266_out1 XOR Logical_Operator_out4282_out1;

  Logical_Operator_out5291_out1 <= Logical_Operator_out4267_out1 XOR Logical_Operator_out4283_out1;

  Logical_Operator_out5292_out1 <= Logical_Operator_out4268_out1 XOR Logical_Operator_out4284_out1;

  Logical_Operator_out5293_out1 <= Logical_Operator_out4269_out1 XOR Logical_Operator_out4285_out1;

  Logical_Operator_out5294_out1 <= Logical_Operator_out4270_out1 XOR Logical_Operator_out4286_out1;

  Logical_Operator_out5295_out1 <= Logical_Operator_out4271_out1 XOR Logical_Operator_out4287_out1;

  Logical_Operator_out5296_out1 <= Logical_Operator_out4272_out1 XOR Logical_Operator_out4288_out1;

  Logical_Operator_out5297_out1 <= Logical_Operator_out3241_out1 XOR Logical_Operator_out3257_out1;

  Logical_Operator_out5298_out1 <= Logical_Operator_out3242_out1 XOR Logical_Operator_out3258_out1;

  Logical_Operator_out5299_out1 <= Logical_Operator_out3243_out1 XOR Logical_Operator_out3259_out1;

  Logical_Operator_out5300_out1 <= Logical_Operator_out3244_out1 XOR Logical_Operator_out3260_out1;

  Logical_Operator_out5301_out1 <= Logical_Operator_out3245_out1 XOR Logical_Operator_out3261_out1;

  Logical_Operator_out5302_out1 <= Logical_Operator_out3246_out1 XOR Logical_Operator_out3262_out1;

  Logical_Operator_out5303_out1 <= Logical_Operator_out3247_out1 XOR Logical_Operator_out3263_out1;

  Logical_Operator_out5304_out1 <= Logical_Operator_out3248_out1 XOR Logical_Operator_out3264_out1;

  Logical_Operator_out5305_out1 <= Logical_Operator_out2221_out1 XOR Logical_Operator_out2237_out1;

  Logical_Operator_out5306_out1 <= Logical_Operator_out2222_out1 XOR Logical_Operator_out2238_out1;

  Logical_Operator_out5307_out1 <= Logical_Operator_out2223_out1 XOR Logical_Operator_out2239_out1;

  Logical_Operator_out5308_out1 <= Logical_Operator_out2224_out1 XOR Logical_Operator_out2240_out1;

  Logical_Operator_out5309_out1 <= Logical_Operator_out1199_out1 XOR Logical_Operator_out1215_out1;

  Logical_Operator_out5310_out1 <= Logical_Operator_out1200_out1 XOR Logical_Operator_out1216_out1;

  Logical_Operator_out5311_out1 <= Logical_Operator_out176_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out5312_out1 <= in352 XOR in384;

  Logical_Operator_out5313_out1 <= Logical_Operator_out4289_out1 XOR Logical_Operator_out4305_out1;

  Logical_Operator_out5314_out1 <= Logical_Operator_out4290_out1 XOR Logical_Operator_out4306_out1;

  Logical_Operator_out5315_out1 <= Logical_Operator_out4291_out1 XOR Logical_Operator_out4307_out1;

  Logical_Operator_out5316_out1 <= Logical_Operator_out4292_out1 XOR Logical_Operator_out4308_out1;

  Logical_Operator_out5317_out1 <= Logical_Operator_out4293_out1 XOR Logical_Operator_out4309_out1;

  Logical_Operator_out5318_out1 <= Logical_Operator_out4294_out1 XOR Logical_Operator_out4310_out1;

  Logical_Operator_out5319_out1 <= Logical_Operator_out4295_out1 XOR Logical_Operator_out4311_out1;

  Logical_Operator_out5320_out1 <= Logical_Operator_out4296_out1 XOR Logical_Operator_out4312_out1;

  Logical_Operator_out5321_out1 <= Logical_Operator_out4297_out1 XOR Logical_Operator_out4313_out1;

  Logical_Operator_out5322_out1 <= Logical_Operator_out4298_out1 XOR Logical_Operator_out4314_out1;

  Logical_Operator_out5323_out1 <= Logical_Operator_out4299_out1 XOR Logical_Operator_out4315_out1;

  Logical_Operator_out5324_out1 <= Logical_Operator_out4300_out1 XOR Logical_Operator_out4316_out1;

  Logical_Operator_out5325_out1 <= Logical_Operator_out4301_out1 XOR Logical_Operator_out4317_out1;

  Logical_Operator_out5326_out1 <= Logical_Operator_out4302_out1 XOR Logical_Operator_out4318_out1;

  Logical_Operator_out5327_out1 <= Logical_Operator_out4303_out1 XOR Logical_Operator_out4319_out1;

  Logical_Operator_out5328_out1 <= Logical_Operator_out4304_out1 XOR Logical_Operator_out4320_out1;

  Logical_Operator_out5329_out1 <= Logical_Operator_out3273_out1 XOR Logical_Operator_out3289_out1;

  Logical_Operator_out5330_out1 <= Logical_Operator_out3274_out1 XOR Logical_Operator_out3290_out1;

  Logical_Operator_out5331_out1 <= Logical_Operator_out3275_out1 XOR Logical_Operator_out3291_out1;

  Logical_Operator_out5332_out1 <= Logical_Operator_out3276_out1 XOR Logical_Operator_out3292_out1;

  Logical_Operator_out5333_out1 <= Logical_Operator_out3277_out1 XOR Logical_Operator_out3293_out1;

  Logical_Operator_out5334_out1 <= Logical_Operator_out3278_out1 XOR Logical_Operator_out3294_out1;

  Logical_Operator_out5335_out1 <= Logical_Operator_out3279_out1 XOR Logical_Operator_out3295_out1;

  Logical_Operator_out5336_out1 <= Logical_Operator_out3280_out1 XOR Logical_Operator_out3296_out1;

  Logical_Operator_out5337_out1 <= Logical_Operator_out2253_out1 XOR Logical_Operator_out2269_out1;

  Logical_Operator_out5338_out1 <= Logical_Operator_out2254_out1 XOR Logical_Operator_out2270_out1;

  Logical_Operator_out5339_out1 <= Logical_Operator_out2255_out1 XOR Logical_Operator_out2271_out1;

  Logical_Operator_out5340_out1 <= Logical_Operator_out2256_out1 XOR Logical_Operator_out2272_out1;

  Logical_Operator_out5341_out1 <= Logical_Operator_out1231_out1 XOR Logical_Operator_out1247_out1;

  Logical_Operator_out5342_out1 <= Logical_Operator_out1232_out1 XOR Logical_Operator_out1248_out1;

  Logical_Operator_out5343_out1 <= Logical_Operator_out208_out1 XOR Logical_Operator_out224_out1;

  Logical_Operator_out5344_out1 <= in416 XOR in448;

  Logical_Operator_out5345_out1 <= Logical_Operator_out4321_out1 XOR Logical_Operator_out4337_out1;

  Logical_Operator_out5346_out1 <= Logical_Operator_out4322_out1 XOR Logical_Operator_out4338_out1;

  Logical_Operator_out5347_out1 <= Logical_Operator_out4323_out1 XOR Logical_Operator_out4339_out1;

  Logical_Operator_out5348_out1 <= Logical_Operator_out4324_out1 XOR Logical_Operator_out4340_out1;

  Logical_Operator_out5349_out1 <= Logical_Operator_out4325_out1 XOR Logical_Operator_out4341_out1;

  Logical_Operator_out5350_out1 <= Logical_Operator_out4326_out1 XOR Logical_Operator_out4342_out1;

  Logical_Operator_out5351_out1 <= Logical_Operator_out4327_out1 XOR Logical_Operator_out4343_out1;

  Logical_Operator_out5352_out1 <= Logical_Operator_out4328_out1 XOR Logical_Operator_out4344_out1;

  Logical_Operator_out5353_out1 <= Logical_Operator_out4329_out1 XOR Logical_Operator_out4345_out1;

  Logical_Operator_out5354_out1 <= Logical_Operator_out4330_out1 XOR Logical_Operator_out4346_out1;

  Logical_Operator_out5355_out1 <= Logical_Operator_out4331_out1 XOR Logical_Operator_out4347_out1;

  Logical_Operator_out5356_out1 <= Logical_Operator_out4332_out1 XOR Logical_Operator_out4348_out1;

  Logical_Operator_out5357_out1 <= Logical_Operator_out4333_out1 XOR Logical_Operator_out4349_out1;

  Logical_Operator_out5358_out1 <= Logical_Operator_out4334_out1 XOR Logical_Operator_out4350_out1;

  Logical_Operator_out5359_out1 <= Logical_Operator_out4335_out1 XOR Logical_Operator_out4351_out1;

  Logical_Operator_out5360_out1 <= Logical_Operator_out4336_out1 XOR Logical_Operator_out4352_out1;

  Logical_Operator_out5361_out1 <= Logical_Operator_out3305_out1 XOR Logical_Operator_out3321_out1;

  Logical_Operator_out5362_out1 <= Logical_Operator_out3306_out1 XOR Logical_Operator_out3322_out1;

  Logical_Operator_out5363_out1 <= Logical_Operator_out3307_out1 XOR Logical_Operator_out3323_out1;

  Logical_Operator_out5364_out1 <= Logical_Operator_out3308_out1 XOR Logical_Operator_out3324_out1;

  Logical_Operator_out5365_out1 <= Logical_Operator_out3309_out1 XOR Logical_Operator_out3325_out1;

  Logical_Operator_out5366_out1 <= Logical_Operator_out3310_out1 XOR Logical_Operator_out3326_out1;

  Logical_Operator_out5367_out1 <= Logical_Operator_out3311_out1 XOR Logical_Operator_out3327_out1;

  Logical_Operator_out5368_out1 <= Logical_Operator_out3312_out1 XOR Logical_Operator_out3328_out1;

  Logical_Operator_out5369_out1 <= Logical_Operator_out2285_out1 XOR Logical_Operator_out2301_out1;

  Logical_Operator_out5370_out1 <= Logical_Operator_out2286_out1 XOR Logical_Operator_out2302_out1;

  Logical_Operator_out5371_out1 <= Logical_Operator_out2287_out1 XOR Logical_Operator_out2303_out1;

  Logical_Operator_out5372_out1 <= Logical_Operator_out2288_out1 XOR Logical_Operator_out2304_out1;

  Logical_Operator_out5373_out1 <= Logical_Operator_out1263_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out5374_out1 <= Logical_Operator_out1264_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out5375_out1 <= Logical_Operator_out240_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out5376_out1 <= in480 XOR in512;

  Logical_Operator_out5377_out1 <= Logical_Operator_out4353_out1 XOR Logical_Operator_out4369_out1;

  Logical_Operator_out5378_out1 <= Logical_Operator_out4354_out1 XOR Logical_Operator_out4370_out1;

  Logical_Operator_out5379_out1 <= Logical_Operator_out4355_out1 XOR Logical_Operator_out4371_out1;

  Logical_Operator_out5380_out1 <= Logical_Operator_out4356_out1 XOR Logical_Operator_out4372_out1;

  Logical_Operator_out5381_out1 <= Logical_Operator_out4357_out1 XOR Logical_Operator_out4373_out1;

  Logical_Operator_out5382_out1 <= Logical_Operator_out4358_out1 XOR Logical_Operator_out4374_out1;

  Logical_Operator_out5383_out1 <= Logical_Operator_out4359_out1 XOR Logical_Operator_out4375_out1;

  Logical_Operator_out5384_out1 <= Logical_Operator_out4360_out1 XOR Logical_Operator_out4376_out1;

  Logical_Operator_out5385_out1 <= Logical_Operator_out4361_out1 XOR Logical_Operator_out4377_out1;

  Logical_Operator_out5386_out1 <= Logical_Operator_out4362_out1 XOR Logical_Operator_out4378_out1;

  Logical_Operator_out5387_out1 <= Logical_Operator_out4363_out1 XOR Logical_Operator_out4379_out1;

  Logical_Operator_out5388_out1 <= Logical_Operator_out4364_out1 XOR Logical_Operator_out4380_out1;

  Logical_Operator_out5389_out1 <= Logical_Operator_out4365_out1 XOR Logical_Operator_out4381_out1;

  Logical_Operator_out5390_out1 <= Logical_Operator_out4366_out1 XOR Logical_Operator_out4382_out1;

  Logical_Operator_out5391_out1 <= Logical_Operator_out4367_out1 XOR Logical_Operator_out4383_out1;

  Logical_Operator_out5392_out1 <= Logical_Operator_out4368_out1 XOR Logical_Operator_out4384_out1;

  Logical_Operator_out5393_out1 <= Logical_Operator_out3337_out1 XOR Logical_Operator_out3353_out1;

  Logical_Operator_out5394_out1 <= Logical_Operator_out3338_out1 XOR Logical_Operator_out3354_out1;

  Logical_Operator_out5395_out1 <= Logical_Operator_out3339_out1 XOR Logical_Operator_out3355_out1;

  Logical_Operator_out5396_out1 <= Logical_Operator_out3340_out1 XOR Logical_Operator_out3356_out1;

  Logical_Operator_out5397_out1 <= Logical_Operator_out3341_out1 XOR Logical_Operator_out3357_out1;

  Logical_Operator_out5398_out1 <= Logical_Operator_out3342_out1 XOR Logical_Operator_out3358_out1;

  Logical_Operator_out5399_out1 <= Logical_Operator_out3343_out1 XOR Logical_Operator_out3359_out1;

  Logical_Operator_out5400_out1 <= Logical_Operator_out3344_out1 XOR Logical_Operator_out3360_out1;

  Logical_Operator_out5401_out1 <= Logical_Operator_out2317_out1 XOR Logical_Operator_out2333_out1;

  Logical_Operator_out5402_out1 <= Logical_Operator_out2318_out1 XOR Logical_Operator_out2334_out1;

  Logical_Operator_out5403_out1 <= Logical_Operator_out2319_out1 XOR Logical_Operator_out2335_out1;

  Logical_Operator_out5404_out1 <= Logical_Operator_out2320_out1 XOR Logical_Operator_out2336_out1;

  Logical_Operator_out5405_out1 <= Logical_Operator_out1295_out1 XOR Logical_Operator_out1311_out1;

  Logical_Operator_out5406_out1 <= Logical_Operator_out1296_out1 XOR Logical_Operator_out1312_out1;

  Logical_Operator_out5407_out1 <= Logical_Operator_out272_out1 XOR Logical_Operator_out288_out1;

  Logical_Operator_out5408_out1 <= in544 XOR in576;

  Logical_Operator_out5409_out1 <= Logical_Operator_out4385_out1 XOR Logical_Operator_out4401_out1;

  Logical_Operator_out5410_out1 <= Logical_Operator_out4386_out1 XOR Logical_Operator_out4402_out1;

  Logical_Operator_out5411_out1 <= Logical_Operator_out4387_out1 XOR Logical_Operator_out4403_out1;

  Logical_Operator_out5412_out1 <= Logical_Operator_out4388_out1 XOR Logical_Operator_out4404_out1;

  Logical_Operator_out5413_out1 <= Logical_Operator_out4389_out1 XOR Logical_Operator_out4405_out1;

  Logical_Operator_out5414_out1 <= Logical_Operator_out4390_out1 XOR Logical_Operator_out4406_out1;

  Logical_Operator_out5415_out1 <= Logical_Operator_out4391_out1 XOR Logical_Operator_out4407_out1;

  Logical_Operator_out5416_out1 <= Logical_Operator_out4392_out1 XOR Logical_Operator_out4408_out1;

  Logical_Operator_out5417_out1 <= Logical_Operator_out4393_out1 XOR Logical_Operator_out4409_out1;

  Logical_Operator_out5418_out1 <= Logical_Operator_out4394_out1 XOR Logical_Operator_out4410_out1;

  Logical_Operator_out5419_out1 <= Logical_Operator_out4395_out1 XOR Logical_Operator_out4411_out1;

  Logical_Operator_out5420_out1 <= Logical_Operator_out4396_out1 XOR Logical_Operator_out4412_out1;

  Logical_Operator_out5421_out1 <= Logical_Operator_out4397_out1 XOR Logical_Operator_out4413_out1;

  Logical_Operator_out5422_out1 <= Logical_Operator_out4398_out1 XOR Logical_Operator_out4414_out1;

  Logical_Operator_out5423_out1 <= Logical_Operator_out4399_out1 XOR Logical_Operator_out4415_out1;

  Logical_Operator_out5424_out1 <= Logical_Operator_out4400_out1 XOR Logical_Operator_out4416_out1;

  Logical_Operator_out5425_out1 <= Logical_Operator_out3369_out1 XOR Logical_Operator_out3385_out1;

  Logical_Operator_out5426_out1 <= Logical_Operator_out3370_out1 XOR Logical_Operator_out3386_out1;

  Logical_Operator_out5427_out1 <= Logical_Operator_out3371_out1 XOR Logical_Operator_out3387_out1;

  Logical_Operator_out5428_out1 <= Logical_Operator_out3372_out1 XOR Logical_Operator_out3388_out1;

  Logical_Operator_out5429_out1 <= Logical_Operator_out3373_out1 XOR Logical_Operator_out3389_out1;

  Logical_Operator_out5430_out1 <= Logical_Operator_out3374_out1 XOR Logical_Operator_out3390_out1;

  Logical_Operator_out5431_out1 <= Logical_Operator_out3375_out1 XOR Logical_Operator_out3391_out1;

  Logical_Operator_out5432_out1 <= Logical_Operator_out3376_out1 XOR Logical_Operator_out3392_out1;

  Logical_Operator_out5433_out1 <= Logical_Operator_out2349_out1 XOR Logical_Operator_out2365_out1;

  Logical_Operator_out5434_out1 <= Logical_Operator_out2350_out1 XOR Logical_Operator_out2366_out1;

  Logical_Operator_out5435_out1 <= Logical_Operator_out2351_out1 XOR Logical_Operator_out2367_out1;

  Logical_Operator_out5436_out1 <= Logical_Operator_out2352_out1 XOR Logical_Operator_out2368_out1;

  Logical_Operator_out5437_out1 <= Logical_Operator_out1327_out1 XOR Logical_Operator_out1343_out1;

  Logical_Operator_out5438_out1 <= Logical_Operator_out1328_out1 XOR Logical_Operator_out1344_out1;

  Logical_Operator_out5439_out1 <= Logical_Operator_out304_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out5440_out1 <= in608 XOR in640;

  Logical_Operator_out5441_out1 <= Logical_Operator_out4417_out1 XOR Logical_Operator_out4433_out1;

  Logical_Operator_out5442_out1 <= Logical_Operator_out4418_out1 XOR Logical_Operator_out4434_out1;

  Logical_Operator_out5443_out1 <= Logical_Operator_out4419_out1 XOR Logical_Operator_out4435_out1;

  Logical_Operator_out5444_out1 <= Logical_Operator_out4420_out1 XOR Logical_Operator_out4436_out1;

  Logical_Operator_out5445_out1 <= Logical_Operator_out4421_out1 XOR Logical_Operator_out4437_out1;

  Logical_Operator_out5446_out1 <= Logical_Operator_out4422_out1 XOR Logical_Operator_out4438_out1;

  Logical_Operator_out5447_out1 <= Logical_Operator_out4423_out1 XOR Logical_Operator_out4439_out1;

  Logical_Operator_out5448_out1 <= Logical_Operator_out4424_out1 XOR Logical_Operator_out4440_out1;

  Logical_Operator_out5449_out1 <= Logical_Operator_out4425_out1 XOR Logical_Operator_out4441_out1;

  Logical_Operator_out5450_out1 <= Logical_Operator_out4426_out1 XOR Logical_Operator_out4442_out1;

  Logical_Operator_out5451_out1 <= Logical_Operator_out4427_out1 XOR Logical_Operator_out4443_out1;

  Logical_Operator_out5452_out1 <= Logical_Operator_out4428_out1 XOR Logical_Operator_out4444_out1;

  Logical_Operator_out5453_out1 <= Logical_Operator_out4429_out1 XOR Logical_Operator_out4445_out1;

  Logical_Operator_out5454_out1 <= Logical_Operator_out4430_out1 XOR Logical_Operator_out4446_out1;

  Logical_Operator_out5455_out1 <= Logical_Operator_out4431_out1 XOR Logical_Operator_out4447_out1;

  Logical_Operator_out5456_out1 <= Logical_Operator_out4432_out1 XOR Logical_Operator_out4448_out1;

  Logical_Operator_out5457_out1 <= Logical_Operator_out3401_out1 XOR Logical_Operator_out3417_out1;

  Logical_Operator_out5458_out1 <= Logical_Operator_out3402_out1 XOR Logical_Operator_out3418_out1;

  Logical_Operator_out5459_out1 <= Logical_Operator_out3403_out1 XOR Logical_Operator_out3419_out1;

  Logical_Operator_out5460_out1 <= Logical_Operator_out3404_out1 XOR Logical_Operator_out3420_out1;

  Logical_Operator_out5461_out1 <= Logical_Operator_out3405_out1 XOR Logical_Operator_out3421_out1;

  Logical_Operator_out5462_out1 <= Logical_Operator_out3406_out1 XOR Logical_Operator_out3422_out1;

  Logical_Operator_out5463_out1 <= Logical_Operator_out3407_out1 XOR Logical_Operator_out3423_out1;

  Logical_Operator_out5464_out1 <= Logical_Operator_out3408_out1 XOR Logical_Operator_out3424_out1;

  Logical_Operator_out5465_out1 <= Logical_Operator_out2381_out1 XOR Logical_Operator_out2397_out1;

  Logical_Operator_out5466_out1 <= Logical_Operator_out2382_out1 XOR Logical_Operator_out2398_out1;

  Logical_Operator_out5467_out1 <= Logical_Operator_out2383_out1 XOR Logical_Operator_out2399_out1;

  Logical_Operator_out5468_out1 <= Logical_Operator_out2384_out1 XOR Logical_Operator_out2400_out1;

  Logical_Operator_out5469_out1 <= Logical_Operator_out1359_out1 XOR Logical_Operator_out1375_out1;

  Logical_Operator_out5470_out1 <= Logical_Operator_out1360_out1 XOR Logical_Operator_out1376_out1;

  Logical_Operator_out5471_out1 <= Logical_Operator_out336_out1 XOR Logical_Operator_out352_out1;

  Logical_Operator_out5472_out1 <= in672 XOR in704;

  Logical_Operator_out5473_out1 <= Logical_Operator_out4449_out1 XOR Logical_Operator_out4465_out1;

  Logical_Operator_out5474_out1 <= Logical_Operator_out4450_out1 XOR Logical_Operator_out4466_out1;

  Logical_Operator_out5475_out1 <= Logical_Operator_out4451_out1 XOR Logical_Operator_out4467_out1;

  Logical_Operator_out5476_out1 <= Logical_Operator_out4452_out1 XOR Logical_Operator_out4468_out1;

  Logical_Operator_out5477_out1 <= Logical_Operator_out4453_out1 XOR Logical_Operator_out4469_out1;

  Logical_Operator_out5478_out1 <= Logical_Operator_out4454_out1 XOR Logical_Operator_out4470_out1;

  Logical_Operator_out5479_out1 <= Logical_Operator_out4455_out1 XOR Logical_Operator_out4471_out1;

  Logical_Operator_out5480_out1 <= Logical_Operator_out4456_out1 XOR Logical_Operator_out4472_out1;

  Logical_Operator_out5481_out1 <= Logical_Operator_out4457_out1 XOR Logical_Operator_out4473_out1;

  Logical_Operator_out5482_out1 <= Logical_Operator_out4458_out1 XOR Logical_Operator_out4474_out1;

  Logical_Operator_out5483_out1 <= Logical_Operator_out4459_out1 XOR Logical_Operator_out4475_out1;

  Logical_Operator_out5484_out1 <= Logical_Operator_out4460_out1 XOR Logical_Operator_out4476_out1;

  Logical_Operator_out5485_out1 <= Logical_Operator_out4461_out1 XOR Logical_Operator_out4477_out1;

  Logical_Operator_out5486_out1 <= Logical_Operator_out4462_out1 XOR Logical_Operator_out4478_out1;

  Logical_Operator_out5487_out1 <= Logical_Operator_out4463_out1 XOR Logical_Operator_out4479_out1;

  Logical_Operator_out5488_out1 <= Logical_Operator_out4464_out1 XOR Logical_Operator_out4480_out1;

  Logical_Operator_out5489_out1 <= Logical_Operator_out3433_out1 XOR Logical_Operator_out3449_out1;

  Logical_Operator_out5490_out1 <= Logical_Operator_out3434_out1 XOR Logical_Operator_out3450_out1;

  Logical_Operator_out5491_out1 <= Logical_Operator_out3435_out1 XOR Logical_Operator_out3451_out1;

  Logical_Operator_out5492_out1 <= Logical_Operator_out3436_out1 XOR Logical_Operator_out3452_out1;

  Logical_Operator_out5493_out1 <= Logical_Operator_out3437_out1 XOR Logical_Operator_out3453_out1;

  Logical_Operator_out5494_out1 <= Logical_Operator_out3438_out1 XOR Logical_Operator_out3454_out1;

  Logical_Operator_out5495_out1 <= Logical_Operator_out3439_out1 XOR Logical_Operator_out3455_out1;

  Logical_Operator_out5496_out1 <= Logical_Operator_out3440_out1 XOR Logical_Operator_out3456_out1;

  Logical_Operator_out5497_out1 <= Logical_Operator_out2413_out1 XOR Logical_Operator_out2429_out1;

  Logical_Operator_out5498_out1 <= Logical_Operator_out2414_out1 XOR Logical_Operator_out2430_out1;

  Logical_Operator_out5499_out1 <= Logical_Operator_out2415_out1 XOR Logical_Operator_out2431_out1;

  Logical_Operator_out5500_out1 <= Logical_Operator_out2416_out1 XOR Logical_Operator_out2432_out1;

  Logical_Operator_out5501_out1 <= Logical_Operator_out1391_out1 XOR Logical_Operator_out1407_out1;

  Logical_Operator_out5502_out1 <= Logical_Operator_out1392_out1 XOR Logical_Operator_out1408_out1;

  Logical_Operator_out5503_out1 <= Logical_Operator_out368_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out5504_out1 <= in736 XOR in768;

  Logical_Operator_out5505_out1 <= Logical_Operator_out4481_out1 XOR Logical_Operator_out4497_out1;

  Logical_Operator_out5506_out1 <= Logical_Operator_out4482_out1 XOR Logical_Operator_out4498_out1;

  Logical_Operator_out5507_out1 <= Logical_Operator_out4483_out1 XOR Logical_Operator_out4499_out1;

  Logical_Operator_out5508_out1 <= Logical_Operator_out4484_out1 XOR Logical_Operator_out4500_out1;

  Logical_Operator_out5509_out1 <= Logical_Operator_out4485_out1 XOR Logical_Operator_out4501_out1;

  Logical_Operator_out5510_out1 <= Logical_Operator_out4486_out1 XOR Logical_Operator_out4502_out1;

  Logical_Operator_out5511_out1 <= Logical_Operator_out4487_out1 XOR Logical_Operator_out4503_out1;

  Logical_Operator_out5512_out1 <= Logical_Operator_out4488_out1 XOR Logical_Operator_out4504_out1;

  Logical_Operator_out5513_out1 <= Logical_Operator_out4489_out1 XOR Logical_Operator_out4505_out1;

  Logical_Operator_out5514_out1 <= Logical_Operator_out4490_out1 XOR Logical_Operator_out4506_out1;

  Logical_Operator_out5515_out1 <= Logical_Operator_out4491_out1 XOR Logical_Operator_out4507_out1;

  Logical_Operator_out5516_out1 <= Logical_Operator_out4492_out1 XOR Logical_Operator_out4508_out1;

  Logical_Operator_out5517_out1 <= Logical_Operator_out4493_out1 XOR Logical_Operator_out4509_out1;

  Logical_Operator_out5518_out1 <= Logical_Operator_out4494_out1 XOR Logical_Operator_out4510_out1;

  Logical_Operator_out5519_out1 <= Logical_Operator_out4495_out1 XOR Logical_Operator_out4511_out1;

  Logical_Operator_out5520_out1 <= Logical_Operator_out4496_out1 XOR Logical_Operator_out4512_out1;

  Logical_Operator_out5521_out1 <= Logical_Operator_out3465_out1 XOR Logical_Operator_out3481_out1;

  Logical_Operator_out5522_out1 <= Logical_Operator_out3466_out1 XOR Logical_Operator_out3482_out1;

  Logical_Operator_out5523_out1 <= Logical_Operator_out3467_out1 XOR Logical_Operator_out3483_out1;

  Logical_Operator_out5524_out1 <= Logical_Operator_out3468_out1 XOR Logical_Operator_out3484_out1;

  Logical_Operator_out5525_out1 <= Logical_Operator_out3469_out1 XOR Logical_Operator_out3485_out1;

  Logical_Operator_out5526_out1 <= Logical_Operator_out3470_out1 XOR Logical_Operator_out3486_out1;

  Logical_Operator_out5527_out1 <= Logical_Operator_out3471_out1 XOR Logical_Operator_out3487_out1;

  Logical_Operator_out5528_out1 <= Logical_Operator_out3472_out1 XOR Logical_Operator_out3488_out1;

  Logical_Operator_out5529_out1 <= Logical_Operator_out2445_out1 XOR Logical_Operator_out2461_out1;

  Logical_Operator_out5530_out1 <= Logical_Operator_out2446_out1 XOR Logical_Operator_out2462_out1;

  Logical_Operator_out5531_out1 <= Logical_Operator_out2447_out1 XOR Logical_Operator_out2463_out1;

  Logical_Operator_out5532_out1 <= Logical_Operator_out2448_out1 XOR Logical_Operator_out2464_out1;

  Logical_Operator_out5533_out1 <= Logical_Operator_out1423_out1 XOR Logical_Operator_out1439_out1;

  Logical_Operator_out5534_out1 <= Logical_Operator_out1424_out1 XOR Logical_Operator_out1440_out1;

  Logical_Operator_out5535_out1 <= Logical_Operator_out400_out1 XOR Logical_Operator_out416_out1;

  Logical_Operator_out5536_out1 <= in800 XOR in832;

  Logical_Operator_out5537_out1 <= Logical_Operator_out4513_out1 XOR Logical_Operator_out4529_out1;

  Logical_Operator_out5538_out1 <= Logical_Operator_out4514_out1 XOR Logical_Operator_out4530_out1;

  Logical_Operator_out5539_out1 <= Logical_Operator_out4515_out1 XOR Logical_Operator_out4531_out1;

  Logical_Operator_out5540_out1 <= Logical_Operator_out4516_out1 XOR Logical_Operator_out4532_out1;

  Logical_Operator_out5541_out1 <= Logical_Operator_out4517_out1 XOR Logical_Operator_out4533_out1;

  Logical_Operator_out5542_out1 <= Logical_Operator_out4518_out1 XOR Logical_Operator_out4534_out1;

  Logical_Operator_out5543_out1 <= Logical_Operator_out4519_out1 XOR Logical_Operator_out4535_out1;

  Logical_Operator_out5544_out1 <= Logical_Operator_out4520_out1 XOR Logical_Operator_out4536_out1;

  Logical_Operator_out5545_out1 <= Logical_Operator_out4521_out1 XOR Logical_Operator_out4537_out1;

  Logical_Operator_out5546_out1 <= Logical_Operator_out4522_out1 XOR Logical_Operator_out4538_out1;

  Logical_Operator_out5547_out1 <= Logical_Operator_out4523_out1 XOR Logical_Operator_out4539_out1;

  Logical_Operator_out5548_out1 <= Logical_Operator_out4524_out1 XOR Logical_Operator_out4540_out1;

  Logical_Operator_out5549_out1 <= Logical_Operator_out4525_out1 XOR Logical_Operator_out4541_out1;

  Logical_Operator_out5550_out1 <= Logical_Operator_out4526_out1 XOR Logical_Operator_out4542_out1;

  Logical_Operator_out5551_out1 <= Logical_Operator_out4527_out1 XOR Logical_Operator_out4543_out1;

  Logical_Operator_out5552_out1 <= Logical_Operator_out4528_out1 XOR Logical_Operator_out4544_out1;

  Logical_Operator_out5553_out1 <= Logical_Operator_out3497_out1 XOR Logical_Operator_out3513_out1;

  Logical_Operator_out5554_out1 <= Logical_Operator_out3498_out1 XOR Logical_Operator_out3514_out1;

  Logical_Operator_out5555_out1 <= Logical_Operator_out3499_out1 XOR Logical_Operator_out3515_out1;

  Logical_Operator_out5556_out1 <= Logical_Operator_out3500_out1 XOR Logical_Operator_out3516_out1;

  Logical_Operator_out5557_out1 <= Logical_Operator_out3501_out1 XOR Logical_Operator_out3517_out1;

  Logical_Operator_out5558_out1 <= Logical_Operator_out3502_out1 XOR Logical_Operator_out3518_out1;

  Logical_Operator_out5559_out1 <= Logical_Operator_out3503_out1 XOR Logical_Operator_out3519_out1;

  Logical_Operator_out5560_out1 <= Logical_Operator_out3504_out1 XOR Logical_Operator_out3520_out1;

  Logical_Operator_out5561_out1 <= Logical_Operator_out2477_out1 XOR Logical_Operator_out2493_out1;

  Logical_Operator_out5562_out1 <= Logical_Operator_out2478_out1 XOR Logical_Operator_out2494_out1;

  Logical_Operator_out5563_out1 <= Logical_Operator_out2479_out1 XOR Logical_Operator_out2495_out1;

  Logical_Operator_out5564_out1 <= Logical_Operator_out2480_out1 XOR Logical_Operator_out2496_out1;

  Logical_Operator_out5565_out1 <= Logical_Operator_out1455_out1 XOR Logical_Operator_out1471_out1;

  Logical_Operator_out5566_out1 <= Logical_Operator_out1456_out1 XOR Logical_Operator_out1472_out1;

  Logical_Operator_out5567_out1 <= Logical_Operator_out432_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out5568_out1 <= in864 XOR in896;

  Logical_Operator_out5569_out1 <= Logical_Operator_out4545_out1 XOR Logical_Operator_out4561_out1;

  Logical_Operator_out5570_out1 <= Logical_Operator_out4546_out1 XOR Logical_Operator_out4562_out1;

  Logical_Operator_out5571_out1 <= Logical_Operator_out4547_out1 XOR Logical_Operator_out4563_out1;

  Logical_Operator_out5572_out1 <= Logical_Operator_out4548_out1 XOR Logical_Operator_out4564_out1;

  Logical_Operator_out5573_out1 <= Logical_Operator_out4549_out1 XOR Logical_Operator_out4565_out1;

  Logical_Operator_out5574_out1 <= Logical_Operator_out4550_out1 XOR Logical_Operator_out4566_out1;

  Logical_Operator_out5575_out1 <= Logical_Operator_out4551_out1 XOR Logical_Operator_out4567_out1;

  Logical_Operator_out5576_out1 <= Logical_Operator_out4552_out1 XOR Logical_Operator_out4568_out1;

  Logical_Operator_out5577_out1 <= Logical_Operator_out4553_out1 XOR Logical_Operator_out4569_out1;

  Logical_Operator_out5578_out1 <= Logical_Operator_out4554_out1 XOR Logical_Operator_out4570_out1;

  Logical_Operator_out5579_out1 <= Logical_Operator_out4555_out1 XOR Logical_Operator_out4571_out1;

  Logical_Operator_out5580_out1 <= Logical_Operator_out4556_out1 XOR Logical_Operator_out4572_out1;

  Logical_Operator_out5581_out1 <= Logical_Operator_out4557_out1 XOR Logical_Operator_out4573_out1;

  Logical_Operator_out5582_out1 <= Logical_Operator_out4558_out1 XOR Logical_Operator_out4574_out1;

  Logical_Operator_out5583_out1 <= Logical_Operator_out4559_out1 XOR Logical_Operator_out4575_out1;

  Logical_Operator_out5584_out1 <= Logical_Operator_out4560_out1 XOR Logical_Operator_out4576_out1;

  Logical_Operator_out5585_out1 <= Logical_Operator_out3529_out1 XOR Logical_Operator_out3545_out1;

  Logical_Operator_out5586_out1 <= Logical_Operator_out3530_out1 XOR Logical_Operator_out3546_out1;

  Logical_Operator_out5587_out1 <= Logical_Operator_out3531_out1 XOR Logical_Operator_out3547_out1;

  Logical_Operator_out5588_out1 <= Logical_Operator_out3532_out1 XOR Logical_Operator_out3548_out1;

  Logical_Operator_out5589_out1 <= Logical_Operator_out3533_out1 XOR Logical_Operator_out3549_out1;

  Logical_Operator_out5590_out1 <= Logical_Operator_out3534_out1 XOR Logical_Operator_out3550_out1;

  Logical_Operator_out5591_out1 <= Logical_Operator_out3535_out1 XOR Logical_Operator_out3551_out1;

  Logical_Operator_out5592_out1 <= Logical_Operator_out3536_out1 XOR Logical_Operator_out3552_out1;

  Logical_Operator_out5593_out1 <= Logical_Operator_out2509_out1 XOR Logical_Operator_out2525_out1;

  Logical_Operator_out5594_out1 <= Logical_Operator_out2510_out1 XOR Logical_Operator_out2526_out1;

  Logical_Operator_out5595_out1 <= Logical_Operator_out2511_out1 XOR Logical_Operator_out2527_out1;

  Logical_Operator_out5596_out1 <= Logical_Operator_out2512_out1 XOR Logical_Operator_out2528_out1;

  Logical_Operator_out5597_out1 <= Logical_Operator_out1487_out1 XOR Logical_Operator_out1503_out1;

  Logical_Operator_out5598_out1 <= Logical_Operator_out1488_out1 XOR Logical_Operator_out1504_out1;

  Logical_Operator_out5599_out1 <= Logical_Operator_out464_out1 XOR Logical_Operator_out480_out1;

  Logical_Operator_out5600_out1 <= in928 XOR in960;

  Logical_Operator_out5601_out1 <= Logical_Operator_out4577_out1 XOR Logical_Operator_out4593_out1;

  Logical_Operator_out5602_out1 <= Logical_Operator_out4578_out1 XOR Logical_Operator_out4594_out1;

  Logical_Operator_out5603_out1 <= Logical_Operator_out4579_out1 XOR Logical_Operator_out4595_out1;

  Logical_Operator_out5604_out1 <= Logical_Operator_out4580_out1 XOR Logical_Operator_out4596_out1;

  Logical_Operator_out5605_out1 <= Logical_Operator_out4581_out1 XOR Logical_Operator_out4597_out1;

  Logical_Operator_out5606_out1 <= Logical_Operator_out4582_out1 XOR Logical_Operator_out4598_out1;

  Logical_Operator_out5607_out1 <= Logical_Operator_out4583_out1 XOR Logical_Operator_out4599_out1;

  Logical_Operator_out5608_out1 <= Logical_Operator_out4584_out1 XOR Logical_Operator_out4600_out1;

  Logical_Operator_out5609_out1 <= Logical_Operator_out4585_out1 XOR Logical_Operator_out4601_out1;

  Logical_Operator_out5610_out1 <= Logical_Operator_out4586_out1 XOR Logical_Operator_out4602_out1;

  Logical_Operator_out5611_out1 <= Logical_Operator_out4587_out1 XOR Logical_Operator_out4603_out1;

  Logical_Operator_out5612_out1 <= Logical_Operator_out4588_out1 XOR Logical_Operator_out4604_out1;

  Logical_Operator_out5613_out1 <= Logical_Operator_out4589_out1 XOR Logical_Operator_out4605_out1;

  Logical_Operator_out5614_out1 <= Logical_Operator_out4590_out1 XOR Logical_Operator_out4606_out1;

  Logical_Operator_out5615_out1 <= Logical_Operator_out4591_out1 XOR Logical_Operator_out4607_out1;

  Logical_Operator_out5616_out1 <= Logical_Operator_out4592_out1 XOR Logical_Operator_out4608_out1;

  Logical_Operator_out5617_out1 <= Logical_Operator_out3561_out1 XOR Logical_Operator_out3577_out1;

  Logical_Operator_out5618_out1 <= Logical_Operator_out3562_out1 XOR Logical_Operator_out3578_out1;

  Logical_Operator_out5619_out1 <= Logical_Operator_out3563_out1 XOR Logical_Operator_out3579_out1;

  Logical_Operator_out5620_out1 <= Logical_Operator_out3564_out1 XOR Logical_Operator_out3580_out1;

  Logical_Operator_out5621_out1 <= Logical_Operator_out3565_out1 XOR Logical_Operator_out3581_out1;

  Logical_Operator_out5622_out1 <= Logical_Operator_out3566_out1 XOR Logical_Operator_out3582_out1;

  Logical_Operator_out5623_out1 <= Logical_Operator_out3567_out1 XOR Logical_Operator_out3583_out1;

  Logical_Operator_out5624_out1 <= Logical_Operator_out3568_out1 XOR Logical_Operator_out3584_out1;

  Logical_Operator_out5625_out1 <= Logical_Operator_out2541_out1 XOR Logical_Operator_out2557_out1;

  Logical_Operator_out5626_out1 <= Logical_Operator_out2542_out1 XOR Logical_Operator_out2558_out1;

  Logical_Operator_out5627_out1 <= Logical_Operator_out2543_out1 XOR Logical_Operator_out2559_out1;

  Logical_Operator_out5628_out1 <= Logical_Operator_out2544_out1 XOR Logical_Operator_out2560_out1;

  Logical_Operator_out5629_out1 <= Logical_Operator_out1519_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out5630_out1 <= Logical_Operator_out1520_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out5631_out1 <= Logical_Operator_out496_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out5632_out1 <= in992 XOR in1024;

  Logical_Operator_out5633_out1 <= Logical_Operator_out4609_out1 XOR Logical_Operator_out4625_out1;

  Logical_Operator_out5634_out1 <= Logical_Operator_out4610_out1 XOR Logical_Operator_out4626_out1;

  Logical_Operator_out5635_out1 <= Logical_Operator_out4611_out1 XOR Logical_Operator_out4627_out1;

  Logical_Operator_out5636_out1 <= Logical_Operator_out4612_out1 XOR Logical_Operator_out4628_out1;

  Logical_Operator_out5637_out1 <= Logical_Operator_out4613_out1 XOR Logical_Operator_out4629_out1;

  Logical_Operator_out5638_out1 <= Logical_Operator_out4614_out1 XOR Logical_Operator_out4630_out1;

  Logical_Operator_out5639_out1 <= Logical_Operator_out4615_out1 XOR Logical_Operator_out4631_out1;

  Logical_Operator_out5640_out1 <= Logical_Operator_out4616_out1 XOR Logical_Operator_out4632_out1;

  Logical_Operator_out5641_out1 <= Logical_Operator_out4617_out1 XOR Logical_Operator_out4633_out1;

  Logical_Operator_out5642_out1 <= Logical_Operator_out4618_out1 XOR Logical_Operator_out4634_out1;

  Logical_Operator_out5643_out1 <= Logical_Operator_out4619_out1 XOR Logical_Operator_out4635_out1;

  Logical_Operator_out5644_out1 <= Logical_Operator_out4620_out1 XOR Logical_Operator_out4636_out1;

  Logical_Operator_out5645_out1 <= Logical_Operator_out4621_out1 XOR Logical_Operator_out4637_out1;

  Logical_Operator_out5646_out1 <= Logical_Operator_out4622_out1 XOR Logical_Operator_out4638_out1;

  Logical_Operator_out5647_out1 <= Logical_Operator_out4623_out1 XOR Logical_Operator_out4639_out1;

  Logical_Operator_out5648_out1 <= Logical_Operator_out4624_out1 XOR Logical_Operator_out4640_out1;

  Logical_Operator_out5649_out1 <= Logical_Operator_out3593_out1 XOR Logical_Operator_out3609_out1;

  Logical_Operator_out5650_out1 <= Logical_Operator_out3594_out1 XOR Logical_Operator_out3610_out1;

  Logical_Operator_out5651_out1 <= Logical_Operator_out3595_out1 XOR Logical_Operator_out3611_out1;

  Logical_Operator_out5652_out1 <= Logical_Operator_out3596_out1 XOR Logical_Operator_out3612_out1;

  Logical_Operator_out5653_out1 <= Logical_Operator_out3597_out1 XOR Logical_Operator_out3613_out1;

  Logical_Operator_out5654_out1 <= Logical_Operator_out3598_out1 XOR Logical_Operator_out3614_out1;

  Logical_Operator_out5655_out1 <= Logical_Operator_out3599_out1 XOR Logical_Operator_out3615_out1;

  Logical_Operator_out5656_out1 <= Logical_Operator_out3600_out1 XOR Logical_Operator_out3616_out1;

  Logical_Operator_out5657_out1 <= Logical_Operator_out2573_out1 XOR Logical_Operator_out2589_out1;

  Logical_Operator_out5658_out1 <= Logical_Operator_out2574_out1 XOR Logical_Operator_out2590_out1;

  Logical_Operator_out5659_out1 <= Logical_Operator_out2575_out1 XOR Logical_Operator_out2591_out1;

  Logical_Operator_out5660_out1 <= Logical_Operator_out2576_out1 XOR Logical_Operator_out2592_out1;

  Logical_Operator_out5661_out1 <= Logical_Operator_out1551_out1 XOR Logical_Operator_out1567_out1;

  Logical_Operator_out5662_out1 <= Logical_Operator_out1552_out1 XOR Logical_Operator_out1568_out1;

  Logical_Operator_out5663_out1 <= Logical_Operator_out528_out1 XOR Logical_Operator_out544_out1;

  Logical_Operator_out5664_out1 <= in1056 XOR in1088;

  Logical_Operator_out5665_out1 <= Logical_Operator_out4641_out1 XOR Logical_Operator_out4657_out1;

  Logical_Operator_out5666_out1 <= Logical_Operator_out4642_out1 XOR Logical_Operator_out4658_out1;

  Logical_Operator_out5667_out1 <= Logical_Operator_out4643_out1 XOR Logical_Operator_out4659_out1;

  Logical_Operator_out5668_out1 <= Logical_Operator_out4644_out1 XOR Logical_Operator_out4660_out1;

  Logical_Operator_out5669_out1 <= Logical_Operator_out4645_out1 XOR Logical_Operator_out4661_out1;

  Logical_Operator_out5670_out1 <= Logical_Operator_out4646_out1 XOR Logical_Operator_out4662_out1;

  Logical_Operator_out5671_out1 <= Logical_Operator_out4647_out1 XOR Logical_Operator_out4663_out1;

  Logical_Operator_out5672_out1 <= Logical_Operator_out4648_out1 XOR Logical_Operator_out4664_out1;

  Logical_Operator_out5673_out1 <= Logical_Operator_out4649_out1 XOR Logical_Operator_out4665_out1;

  Logical_Operator_out5674_out1 <= Logical_Operator_out4650_out1 XOR Logical_Operator_out4666_out1;

  Logical_Operator_out5675_out1 <= Logical_Operator_out4651_out1 XOR Logical_Operator_out4667_out1;

  Logical_Operator_out5676_out1 <= Logical_Operator_out4652_out1 XOR Logical_Operator_out4668_out1;

  Logical_Operator_out5677_out1 <= Logical_Operator_out4653_out1 XOR Logical_Operator_out4669_out1;

  Logical_Operator_out5678_out1 <= Logical_Operator_out4654_out1 XOR Logical_Operator_out4670_out1;

  Logical_Operator_out5679_out1 <= Logical_Operator_out4655_out1 XOR Logical_Operator_out4671_out1;

  Logical_Operator_out5680_out1 <= Logical_Operator_out4656_out1 XOR Logical_Operator_out4672_out1;

  Logical_Operator_out5681_out1 <= Logical_Operator_out3625_out1 XOR Logical_Operator_out3641_out1;

  Logical_Operator_out5682_out1 <= Logical_Operator_out3626_out1 XOR Logical_Operator_out3642_out1;

  Logical_Operator_out5683_out1 <= Logical_Operator_out3627_out1 XOR Logical_Operator_out3643_out1;

  Logical_Operator_out5684_out1 <= Logical_Operator_out3628_out1 XOR Logical_Operator_out3644_out1;

  Logical_Operator_out5685_out1 <= Logical_Operator_out3629_out1 XOR Logical_Operator_out3645_out1;

  Logical_Operator_out5686_out1 <= Logical_Operator_out3630_out1 XOR Logical_Operator_out3646_out1;

  Logical_Operator_out5687_out1 <= Logical_Operator_out3631_out1 XOR Logical_Operator_out3647_out1;

  Logical_Operator_out5688_out1 <= Logical_Operator_out3632_out1 XOR Logical_Operator_out3648_out1;

  Logical_Operator_out5689_out1 <= Logical_Operator_out2605_out1 XOR Logical_Operator_out2621_out1;

  Logical_Operator_out5690_out1 <= Logical_Operator_out2606_out1 XOR Logical_Operator_out2622_out1;

  Logical_Operator_out5691_out1 <= Logical_Operator_out2607_out1 XOR Logical_Operator_out2623_out1;

  Logical_Operator_out5692_out1 <= Logical_Operator_out2608_out1 XOR Logical_Operator_out2624_out1;

  Logical_Operator_out5693_out1 <= Logical_Operator_out1583_out1 XOR Logical_Operator_out1599_out1;

  Logical_Operator_out5694_out1 <= Logical_Operator_out1584_out1 XOR Logical_Operator_out1600_out1;

  Logical_Operator_out5695_out1 <= Logical_Operator_out560_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out5696_out1 <= in1120 XOR in1152;

  Logical_Operator_out5697_out1 <= Logical_Operator_out4673_out1 XOR Logical_Operator_out4689_out1;

  Logical_Operator_out5698_out1 <= Logical_Operator_out4674_out1 XOR Logical_Operator_out4690_out1;

  Logical_Operator_out5699_out1 <= Logical_Operator_out4675_out1 XOR Logical_Operator_out4691_out1;

  Logical_Operator_out5700_out1 <= Logical_Operator_out4676_out1 XOR Logical_Operator_out4692_out1;

  Logical_Operator_out5701_out1 <= Logical_Operator_out4677_out1 XOR Logical_Operator_out4693_out1;

  Logical_Operator_out5702_out1 <= Logical_Operator_out4678_out1 XOR Logical_Operator_out4694_out1;

  Logical_Operator_out5703_out1 <= Logical_Operator_out4679_out1 XOR Logical_Operator_out4695_out1;

  Logical_Operator_out5704_out1 <= Logical_Operator_out4680_out1 XOR Logical_Operator_out4696_out1;

  Logical_Operator_out5705_out1 <= Logical_Operator_out4681_out1 XOR Logical_Operator_out4697_out1;

  Logical_Operator_out5706_out1 <= Logical_Operator_out4682_out1 XOR Logical_Operator_out4698_out1;

  Logical_Operator_out5707_out1 <= Logical_Operator_out4683_out1 XOR Logical_Operator_out4699_out1;

  Logical_Operator_out5708_out1 <= Logical_Operator_out4684_out1 XOR Logical_Operator_out4700_out1;

  Logical_Operator_out5709_out1 <= Logical_Operator_out4685_out1 XOR Logical_Operator_out4701_out1;

  Logical_Operator_out5710_out1 <= Logical_Operator_out4686_out1 XOR Logical_Operator_out4702_out1;

  Logical_Operator_out5711_out1 <= Logical_Operator_out4687_out1 XOR Logical_Operator_out4703_out1;

  Logical_Operator_out5712_out1 <= Logical_Operator_out4688_out1 XOR Logical_Operator_out4704_out1;

  Logical_Operator_out5713_out1 <= Logical_Operator_out3657_out1 XOR Logical_Operator_out3673_out1;

  Logical_Operator_out5714_out1 <= Logical_Operator_out3658_out1 XOR Logical_Operator_out3674_out1;

  Logical_Operator_out5715_out1 <= Logical_Operator_out3659_out1 XOR Logical_Operator_out3675_out1;

  Logical_Operator_out5716_out1 <= Logical_Operator_out3660_out1 XOR Logical_Operator_out3676_out1;

  Logical_Operator_out5717_out1 <= Logical_Operator_out3661_out1 XOR Logical_Operator_out3677_out1;

  Logical_Operator_out5718_out1 <= Logical_Operator_out3662_out1 XOR Logical_Operator_out3678_out1;

  Logical_Operator_out5719_out1 <= Logical_Operator_out3663_out1 XOR Logical_Operator_out3679_out1;

  Logical_Operator_out5720_out1 <= Logical_Operator_out3664_out1 XOR Logical_Operator_out3680_out1;

  Logical_Operator_out5721_out1 <= Logical_Operator_out2637_out1 XOR Logical_Operator_out2653_out1;

  Logical_Operator_out5722_out1 <= Logical_Operator_out2638_out1 XOR Logical_Operator_out2654_out1;

  Logical_Operator_out5723_out1 <= Logical_Operator_out2639_out1 XOR Logical_Operator_out2655_out1;

  Logical_Operator_out5724_out1 <= Logical_Operator_out2640_out1 XOR Logical_Operator_out2656_out1;

  Logical_Operator_out5725_out1 <= Logical_Operator_out1615_out1 XOR Logical_Operator_out1631_out1;

  Logical_Operator_out5726_out1 <= Logical_Operator_out1616_out1 XOR Logical_Operator_out1632_out1;

  Logical_Operator_out5727_out1 <= Logical_Operator_out592_out1 XOR Logical_Operator_out608_out1;

  Logical_Operator_out5728_out1 <= in1184 XOR in1216;

  Logical_Operator_out5729_out1 <= Logical_Operator_out4705_out1 XOR Logical_Operator_out4721_out1;

  Logical_Operator_out5730_out1 <= Logical_Operator_out4706_out1 XOR Logical_Operator_out4722_out1;

  Logical_Operator_out5731_out1 <= Logical_Operator_out4707_out1 XOR Logical_Operator_out4723_out1;

  Logical_Operator_out5732_out1 <= Logical_Operator_out4708_out1 XOR Logical_Operator_out4724_out1;

  Logical_Operator_out5733_out1 <= Logical_Operator_out4709_out1 XOR Logical_Operator_out4725_out1;

  Logical_Operator_out5734_out1 <= Logical_Operator_out4710_out1 XOR Logical_Operator_out4726_out1;

  Logical_Operator_out5735_out1 <= Logical_Operator_out4711_out1 XOR Logical_Operator_out4727_out1;

  Logical_Operator_out5736_out1 <= Logical_Operator_out4712_out1 XOR Logical_Operator_out4728_out1;

  Logical_Operator_out5737_out1 <= Logical_Operator_out4713_out1 XOR Logical_Operator_out4729_out1;

  Logical_Operator_out5738_out1 <= Logical_Operator_out4714_out1 XOR Logical_Operator_out4730_out1;

  Logical_Operator_out5739_out1 <= Logical_Operator_out4715_out1 XOR Logical_Operator_out4731_out1;

  Logical_Operator_out5740_out1 <= Logical_Operator_out4716_out1 XOR Logical_Operator_out4732_out1;

  Logical_Operator_out5741_out1 <= Logical_Operator_out4717_out1 XOR Logical_Operator_out4733_out1;

  Logical_Operator_out5742_out1 <= Logical_Operator_out4718_out1 XOR Logical_Operator_out4734_out1;

  Logical_Operator_out5743_out1 <= Logical_Operator_out4719_out1 XOR Logical_Operator_out4735_out1;

  Logical_Operator_out5744_out1 <= Logical_Operator_out4720_out1 XOR Logical_Operator_out4736_out1;

  Logical_Operator_out5745_out1 <= Logical_Operator_out3689_out1 XOR Logical_Operator_out3705_out1;

  Logical_Operator_out5746_out1 <= Logical_Operator_out3690_out1 XOR Logical_Operator_out3706_out1;

  Logical_Operator_out5747_out1 <= Logical_Operator_out3691_out1 XOR Logical_Operator_out3707_out1;

  Logical_Operator_out5748_out1 <= Logical_Operator_out3692_out1 XOR Logical_Operator_out3708_out1;

  Logical_Operator_out5749_out1 <= Logical_Operator_out3693_out1 XOR Logical_Operator_out3709_out1;

  Logical_Operator_out5750_out1 <= Logical_Operator_out3694_out1 XOR Logical_Operator_out3710_out1;

  Logical_Operator_out5751_out1 <= Logical_Operator_out3695_out1 XOR Logical_Operator_out3711_out1;

  Logical_Operator_out5752_out1 <= Logical_Operator_out3696_out1 XOR Logical_Operator_out3712_out1;

  Logical_Operator_out5753_out1 <= Logical_Operator_out2669_out1 XOR Logical_Operator_out2685_out1;

  Logical_Operator_out5754_out1 <= Logical_Operator_out2670_out1 XOR Logical_Operator_out2686_out1;

  Logical_Operator_out5755_out1 <= Logical_Operator_out2671_out1 XOR Logical_Operator_out2687_out1;

  Logical_Operator_out5756_out1 <= Logical_Operator_out2672_out1 XOR Logical_Operator_out2688_out1;

  Logical_Operator_out5757_out1 <= Logical_Operator_out1647_out1 XOR Logical_Operator_out1663_out1;

  Logical_Operator_out5758_out1 <= Logical_Operator_out1648_out1 XOR Logical_Operator_out1664_out1;

  Logical_Operator_out5759_out1 <= Logical_Operator_out624_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out5760_out1 <= in1248 XOR in1280;

  Logical_Operator_out5761_out1 <= Logical_Operator_out4737_out1 XOR Logical_Operator_out4753_out1;

  Logical_Operator_out5762_out1 <= Logical_Operator_out4738_out1 XOR Logical_Operator_out4754_out1;

  Logical_Operator_out5763_out1 <= Logical_Operator_out4739_out1 XOR Logical_Operator_out4755_out1;

  Logical_Operator_out5764_out1 <= Logical_Operator_out4740_out1 XOR Logical_Operator_out4756_out1;

  Logical_Operator_out5765_out1 <= Logical_Operator_out4741_out1 XOR Logical_Operator_out4757_out1;

  Logical_Operator_out5766_out1 <= Logical_Operator_out4742_out1 XOR Logical_Operator_out4758_out1;

  Logical_Operator_out5767_out1 <= Logical_Operator_out4743_out1 XOR Logical_Operator_out4759_out1;

  Logical_Operator_out5768_out1 <= Logical_Operator_out4744_out1 XOR Logical_Operator_out4760_out1;

  Logical_Operator_out5769_out1 <= Logical_Operator_out4745_out1 XOR Logical_Operator_out4761_out1;

  Logical_Operator_out5770_out1 <= Logical_Operator_out4746_out1 XOR Logical_Operator_out4762_out1;

  Logical_Operator_out5771_out1 <= Logical_Operator_out4747_out1 XOR Logical_Operator_out4763_out1;

  Logical_Operator_out5772_out1 <= Logical_Operator_out4748_out1 XOR Logical_Operator_out4764_out1;

  Logical_Operator_out5773_out1 <= Logical_Operator_out4749_out1 XOR Logical_Operator_out4765_out1;

  Logical_Operator_out5774_out1 <= Logical_Operator_out4750_out1 XOR Logical_Operator_out4766_out1;

  Logical_Operator_out5775_out1 <= Logical_Operator_out4751_out1 XOR Logical_Operator_out4767_out1;

  Logical_Operator_out5776_out1 <= Logical_Operator_out4752_out1 XOR Logical_Operator_out4768_out1;

  Logical_Operator_out5777_out1 <= Logical_Operator_out3721_out1 XOR Logical_Operator_out3737_out1;

  Logical_Operator_out5778_out1 <= Logical_Operator_out3722_out1 XOR Logical_Operator_out3738_out1;

  Logical_Operator_out5779_out1 <= Logical_Operator_out3723_out1 XOR Logical_Operator_out3739_out1;

  Logical_Operator_out5780_out1 <= Logical_Operator_out3724_out1 XOR Logical_Operator_out3740_out1;

  Logical_Operator_out5781_out1 <= Logical_Operator_out3725_out1 XOR Logical_Operator_out3741_out1;

  Logical_Operator_out5782_out1 <= Logical_Operator_out3726_out1 XOR Logical_Operator_out3742_out1;

  Logical_Operator_out5783_out1 <= Logical_Operator_out3727_out1 XOR Logical_Operator_out3743_out1;

  Logical_Operator_out5784_out1 <= Logical_Operator_out3728_out1 XOR Logical_Operator_out3744_out1;

  Logical_Operator_out5785_out1 <= Logical_Operator_out2701_out1 XOR Logical_Operator_out2717_out1;

  Logical_Operator_out5786_out1 <= Logical_Operator_out2702_out1 XOR Logical_Operator_out2718_out1;

  Logical_Operator_out5787_out1 <= Logical_Operator_out2703_out1 XOR Logical_Operator_out2719_out1;

  Logical_Operator_out5788_out1 <= Logical_Operator_out2704_out1 XOR Logical_Operator_out2720_out1;

  Logical_Operator_out5789_out1 <= Logical_Operator_out1679_out1 XOR Logical_Operator_out1695_out1;

  Logical_Operator_out5790_out1 <= Logical_Operator_out1680_out1 XOR Logical_Operator_out1696_out1;

  Logical_Operator_out5791_out1 <= Logical_Operator_out656_out1 XOR Logical_Operator_out672_out1;

  Logical_Operator_out5792_out1 <= in1312 XOR in1344;

  Logical_Operator_out5793_out1 <= Logical_Operator_out4769_out1 XOR Logical_Operator_out4785_out1;

  Logical_Operator_out5794_out1 <= Logical_Operator_out4770_out1 XOR Logical_Operator_out4786_out1;

  Logical_Operator_out5795_out1 <= Logical_Operator_out4771_out1 XOR Logical_Operator_out4787_out1;

  Logical_Operator_out5796_out1 <= Logical_Operator_out4772_out1 XOR Logical_Operator_out4788_out1;

  Logical_Operator_out5797_out1 <= Logical_Operator_out4773_out1 XOR Logical_Operator_out4789_out1;

  Logical_Operator_out5798_out1 <= Logical_Operator_out4774_out1 XOR Logical_Operator_out4790_out1;

  Logical_Operator_out5799_out1 <= Logical_Operator_out4775_out1 XOR Logical_Operator_out4791_out1;

  Logical_Operator_out5800_out1 <= Logical_Operator_out4776_out1 XOR Logical_Operator_out4792_out1;

  Logical_Operator_out5801_out1 <= Logical_Operator_out4777_out1 XOR Logical_Operator_out4793_out1;

  Logical_Operator_out5802_out1 <= Logical_Operator_out4778_out1 XOR Logical_Operator_out4794_out1;

  Logical_Operator_out5803_out1 <= Logical_Operator_out4779_out1 XOR Logical_Operator_out4795_out1;

  Logical_Operator_out5804_out1 <= Logical_Operator_out4780_out1 XOR Logical_Operator_out4796_out1;

  Logical_Operator_out5805_out1 <= Logical_Operator_out4781_out1 XOR Logical_Operator_out4797_out1;

  Logical_Operator_out5806_out1 <= Logical_Operator_out4782_out1 XOR Logical_Operator_out4798_out1;

  Logical_Operator_out5807_out1 <= Logical_Operator_out4783_out1 XOR Logical_Operator_out4799_out1;

  Logical_Operator_out5808_out1 <= Logical_Operator_out4784_out1 XOR Logical_Operator_out4800_out1;

  Logical_Operator_out5809_out1 <= Logical_Operator_out3753_out1 XOR Logical_Operator_out3769_out1;

  Logical_Operator_out5810_out1 <= Logical_Operator_out3754_out1 XOR Logical_Operator_out3770_out1;

  Logical_Operator_out5811_out1 <= Logical_Operator_out3755_out1 XOR Logical_Operator_out3771_out1;

  Logical_Operator_out5812_out1 <= Logical_Operator_out3756_out1 XOR Logical_Operator_out3772_out1;

  Logical_Operator_out5813_out1 <= Logical_Operator_out3757_out1 XOR Logical_Operator_out3773_out1;

  Logical_Operator_out5814_out1 <= Logical_Operator_out3758_out1 XOR Logical_Operator_out3774_out1;

  Logical_Operator_out5815_out1 <= Logical_Operator_out3759_out1 XOR Logical_Operator_out3775_out1;

  Logical_Operator_out5816_out1 <= Logical_Operator_out3760_out1 XOR Logical_Operator_out3776_out1;

  Logical_Operator_out5817_out1 <= Logical_Operator_out2733_out1 XOR Logical_Operator_out2749_out1;

  Logical_Operator_out5818_out1 <= Logical_Operator_out2734_out1 XOR Logical_Operator_out2750_out1;

  Logical_Operator_out5819_out1 <= Logical_Operator_out2735_out1 XOR Logical_Operator_out2751_out1;

  Logical_Operator_out5820_out1 <= Logical_Operator_out2736_out1 XOR Logical_Operator_out2752_out1;

  Logical_Operator_out5821_out1 <= Logical_Operator_out1711_out1 XOR Logical_Operator_out1727_out1;

  Logical_Operator_out5822_out1 <= Logical_Operator_out1712_out1 XOR Logical_Operator_out1728_out1;

  Logical_Operator_out5823_out1 <= Logical_Operator_out688_out1 XOR Logical_Operator_out704_out1;

  Logical_Operator_out5824_out1 <= in1376 XOR in1408;

  Logical_Operator_out5825_out1 <= Logical_Operator_out4801_out1 XOR Logical_Operator_out4817_out1;

  Logical_Operator_out5826_out1 <= Logical_Operator_out4802_out1 XOR Logical_Operator_out4818_out1;

  Logical_Operator_out5827_out1 <= Logical_Operator_out4803_out1 XOR Logical_Operator_out4819_out1;

  Logical_Operator_out5828_out1 <= Logical_Operator_out4804_out1 XOR Logical_Operator_out4820_out1;

  Logical_Operator_out5829_out1 <= Logical_Operator_out4805_out1 XOR Logical_Operator_out4821_out1;

  Logical_Operator_out5830_out1 <= Logical_Operator_out4806_out1 XOR Logical_Operator_out4822_out1;

  Logical_Operator_out5831_out1 <= Logical_Operator_out4807_out1 XOR Logical_Operator_out4823_out1;

  Logical_Operator_out5832_out1 <= Logical_Operator_out4808_out1 XOR Logical_Operator_out4824_out1;

  Logical_Operator_out5833_out1 <= Logical_Operator_out4809_out1 XOR Logical_Operator_out4825_out1;

  Logical_Operator_out5834_out1 <= Logical_Operator_out4810_out1 XOR Logical_Operator_out4826_out1;

  Logical_Operator_out5835_out1 <= Logical_Operator_out4811_out1 XOR Logical_Operator_out4827_out1;

  Logical_Operator_out5836_out1 <= Logical_Operator_out4812_out1 XOR Logical_Operator_out4828_out1;

  Logical_Operator_out5837_out1 <= Logical_Operator_out4813_out1 XOR Logical_Operator_out4829_out1;

  Logical_Operator_out5838_out1 <= Logical_Operator_out4814_out1 XOR Logical_Operator_out4830_out1;

  Logical_Operator_out5839_out1 <= Logical_Operator_out4815_out1 XOR Logical_Operator_out4831_out1;

  Logical_Operator_out5840_out1 <= Logical_Operator_out4816_out1 XOR Logical_Operator_out4832_out1;

  Logical_Operator_out5841_out1 <= Logical_Operator_out3785_out1 XOR Logical_Operator_out3801_out1;

  Logical_Operator_out5842_out1 <= Logical_Operator_out3786_out1 XOR Logical_Operator_out3802_out1;

  Logical_Operator_out5843_out1 <= Logical_Operator_out3787_out1 XOR Logical_Operator_out3803_out1;

  Logical_Operator_out5844_out1 <= Logical_Operator_out3788_out1 XOR Logical_Operator_out3804_out1;

  Logical_Operator_out5845_out1 <= Logical_Operator_out3789_out1 XOR Logical_Operator_out3805_out1;

  Logical_Operator_out5846_out1 <= Logical_Operator_out3790_out1 XOR Logical_Operator_out3806_out1;

  Logical_Operator_out5847_out1 <= Logical_Operator_out3791_out1 XOR Logical_Operator_out3807_out1;

  Logical_Operator_out5848_out1 <= Logical_Operator_out3792_out1 XOR Logical_Operator_out3808_out1;

  Logical_Operator_out5849_out1 <= Logical_Operator_out2765_out1 XOR Logical_Operator_out2781_out1;

  Logical_Operator_out5850_out1 <= Logical_Operator_out2766_out1 XOR Logical_Operator_out2782_out1;

  Logical_Operator_out5851_out1 <= Logical_Operator_out2767_out1 XOR Logical_Operator_out2783_out1;

  Logical_Operator_out5852_out1 <= Logical_Operator_out2768_out1 XOR Logical_Operator_out2784_out1;

  Logical_Operator_out5853_out1 <= Logical_Operator_out1743_out1 XOR Logical_Operator_out1759_out1;

  Logical_Operator_out5854_out1 <= Logical_Operator_out1744_out1 XOR Logical_Operator_out1760_out1;

  Logical_Operator_out5855_out1 <= Logical_Operator_out720_out1 XOR Logical_Operator_out736_out1;

  Logical_Operator_out5856_out1 <= in1440 XOR in1472;

  Logical_Operator_out5857_out1 <= Logical_Operator_out4833_out1 XOR Logical_Operator_out4849_out1;

  Logical_Operator_out5858_out1 <= Logical_Operator_out4834_out1 XOR Logical_Operator_out4850_out1;

  Logical_Operator_out5859_out1 <= Logical_Operator_out4835_out1 XOR Logical_Operator_out4851_out1;

  Logical_Operator_out5860_out1 <= Logical_Operator_out4836_out1 XOR Logical_Operator_out4852_out1;

  Logical_Operator_out5861_out1 <= Logical_Operator_out4837_out1 XOR Logical_Operator_out4853_out1;

  Logical_Operator_out5862_out1 <= Logical_Operator_out4838_out1 XOR Logical_Operator_out4854_out1;

  Logical_Operator_out5863_out1 <= Logical_Operator_out4839_out1 XOR Logical_Operator_out4855_out1;

  Logical_Operator_out5864_out1 <= Logical_Operator_out4840_out1 XOR Logical_Operator_out4856_out1;

  Logical_Operator_out5865_out1 <= Logical_Operator_out4841_out1 XOR Logical_Operator_out4857_out1;

  Logical_Operator_out5866_out1 <= Logical_Operator_out4842_out1 XOR Logical_Operator_out4858_out1;

  Logical_Operator_out5867_out1 <= Logical_Operator_out4843_out1 XOR Logical_Operator_out4859_out1;

  Logical_Operator_out5868_out1 <= Logical_Operator_out4844_out1 XOR Logical_Operator_out4860_out1;

  Logical_Operator_out5869_out1 <= Logical_Operator_out4845_out1 XOR Logical_Operator_out4861_out1;

  Logical_Operator_out5870_out1 <= Logical_Operator_out4846_out1 XOR Logical_Operator_out4862_out1;

  Logical_Operator_out5871_out1 <= Logical_Operator_out4847_out1 XOR Logical_Operator_out4863_out1;

  Logical_Operator_out5872_out1 <= Logical_Operator_out4848_out1 XOR Logical_Operator_out4864_out1;

  Logical_Operator_out5873_out1 <= Logical_Operator_out3817_out1 XOR Logical_Operator_out3833_out1;

  Logical_Operator_out5874_out1 <= Logical_Operator_out3818_out1 XOR Logical_Operator_out3834_out1;

  Logical_Operator_out5875_out1 <= Logical_Operator_out3819_out1 XOR Logical_Operator_out3835_out1;

  Logical_Operator_out5876_out1 <= Logical_Operator_out3820_out1 XOR Logical_Operator_out3836_out1;

  Logical_Operator_out5877_out1 <= Logical_Operator_out3821_out1 XOR Logical_Operator_out3837_out1;

  Logical_Operator_out5878_out1 <= Logical_Operator_out3822_out1 XOR Logical_Operator_out3838_out1;

  Logical_Operator_out5879_out1 <= Logical_Operator_out3823_out1 XOR Logical_Operator_out3839_out1;

  Logical_Operator_out5880_out1 <= Logical_Operator_out3824_out1 XOR Logical_Operator_out3840_out1;

  Logical_Operator_out5881_out1 <= Logical_Operator_out2797_out1 XOR Logical_Operator_out2813_out1;

  Logical_Operator_out5882_out1 <= Logical_Operator_out2798_out1 XOR Logical_Operator_out2814_out1;

  Logical_Operator_out5883_out1 <= Logical_Operator_out2799_out1 XOR Logical_Operator_out2815_out1;

  Logical_Operator_out5884_out1 <= Logical_Operator_out2800_out1 XOR Logical_Operator_out2816_out1;

  Logical_Operator_out5885_out1 <= Logical_Operator_out1775_out1 XOR Logical_Operator_out1791_out1;

  Logical_Operator_out5886_out1 <= Logical_Operator_out1776_out1 XOR Logical_Operator_out1792_out1;

  Logical_Operator_out5887_out1 <= Logical_Operator_out752_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out5888_out1 <= in1504 XOR in1536;

  Logical_Operator_out5889_out1 <= Logical_Operator_out4865_out1 XOR Logical_Operator_out4881_out1;

  Logical_Operator_out5890_out1 <= Logical_Operator_out4866_out1 XOR Logical_Operator_out4882_out1;

  Logical_Operator_out5891_out1 <= Logical_Operator_out4867_out1 XOR Logical_Operator_out4883_out1;

  Logical_Operator_out5892_out1 <= Logical_Operator_out4868_out1 XOR Logical_Operator_out4884_out1;

  Logical_Operator_out5893_out1 <= Logical_Operator_out4869_out1 XOR Logical_Operator_out4885_out1;

  Logical_Operator_out5894_out1 <= Logical_Operator_out4870_out1 XOR Logical_Operator_out4886_out1;

  Logical_Operator_out5895_out1 <= Logical_Operator_out4871_out1 XOR Logical_Operator_out4887_out1;

  Logical_Operator_out5896_out1 <= Logical_Operator_out4872_out1 XOR Logical_Operator_out4888_out1;

  Logical_Operator_out5897_out1 <= Logical_Operator_out4873_out1 XOR Logical_Operator_out4889_out1;

  Logical_Operator_out5898_out1 <= Logical_Operator_out4874_out1 XOR Logical_Operator_out4890_out1;

  Logical_Operator_out5899_out1 <= Logical_Operator_out4875_out1 XOR Logical_Operator_out4891_out1;

  Logical_Operator_out5900_out1 <= Logical_Operator_out4876_out1 XOR Logical_Operator_out4892_out1;

  Logical_Operator_out5901_out1 <= Logical_Operator_out4877_out1 XOR Logical_Operator_out4893_out1;

  Logical_Operator_out5902_out1 <= Logical_Operator_out4878_out1 XOR Logical_Operator_out4894_out1;

  Logical_Operator_out5903_out1 <= Logical_Operator_out4879_out1 XOR Logical_Operator_out4895_out1;

  Logical_Operator_out5904_out1 <= Logical_Operator_out4880_out1 XOR Logical_Operator_out4896_out1;

  Logical_Operator_out5905_out1 <= Logical_Operator_out3849_out1 XOR Logical_Operator_out3865_out1;

  Logical_Operator_out5906_out1 <= Logical_Operator_out3850_out1 XOR Logical_Operator_out3866_out1;

  Logical_Operator_out5907_out1 <= Logical_Operator_out3851_out1 XOR Logical_Operator_out3867_out1;

  Logical_Operator_out5908_out1 <= Logical_Operator_out3852_out1 XOR Logical_Operator_out3868_out1;

  Logical_Operator_out5909_out1 <= Logical_Operator_out3853_out1 XOR Logical_Operator_out3869_out1;

  Logical_Operator_out5910_out1 <= Logical_Operator_out3854_out1 XOR Logical_Operator_out3870_out1;

  Logical_Operator_out5911_out1 <= Logical_Operator_out3855_out1 XOR Logical_Operator_out3871_out1;

  Logical_Operator_out5912_out1 <= Logical_Operator_out3856_out1 XOR Logical_Operator_out3872_out1;

  Logical_Operator_out5913_out1 <= Logical_Operator_out2829_out1 XOR Logical_Operator_out2845_out1;

  Logical_Operator_out5914_out1 <= Logical_Operator_out2830_out1 XOR Logical_Operator_out2846_out1;

  Logical_Operator_out5915_out1 <= Logical_Operator_out2831_out1 XOR Logical_Operator_out2847_out1;

  Logical_Operator_out5916_out1 <= Logical_Operator_out2832_out1 XOR Logical_Operator_out2848_out1;

  Logical_Operator_out5917_out1 <= Logical_Operator_out1807_out1 XOR Logical_Operator_out1823_out1;

  Logical_Operator_out5918_out1 <= Logical_Operator_out1808_out1 XOR Logical_Operator_out1824_out1;

  Logical_Operator_out5919_out1 <= Logical_Operator_out784_out1 XOR Logical_Operator_out800_out1;

  Logical_Operator_out5920_out1 <= in1568 XOR in1600;

  Logical_Operator_out5921_out1 <= Logical_Operator_out4897_out1 XOR Logical_Operator_out4913_out1;

  Logical_Operator_out5922_out1 <= Logical_Operator_out4898_out1 XOR Logical_Operator_out4914_out1;

  Logical_Operator_out5923_out1 <= Logical_Operator_out4899_out1 XOR Logical_Operator_out4915_out1;

  Logical_Operator_out5924_out1 <= Logical_Operator_out4900_out1 XOR Logical_Operator_out4916_out1;

  Logical_Operator_out5925_out1 <= Logical_Operator_out4901_out1 XOR Logical_Operator_out4917_out1;

  Logical_Operator_out5926_out1 <= Logical_Operator_out4902_out1 XOR Logical_Operator_out4918_out1;

  Logical_Operator_out5927_out1 <= Logical_Operator_out4903_out1 XOR Logical_Operator_out4919_out1;

  Logical_Operator_out5928_out1 <= Logical_Operator_out4904_out1 XOR Logical_Operator_out4920_out1;

  Logical_Operator_out5929_out1 <= Logical_Operator_out4905_out1 XOR Logical_Operator_out4921_out1;

  Logical_Operator_out5930_out1 <= Logical_Operator_out4906_out1 XOR Logical_Operator_out4922_out1;

  Logical_Operator_out5931_out1 <= Logical_Operator_out4907_out1 XOR Logical_Operator_out4923_out1;

  Logical_Operator_out5932_out1 <= Logical_Operator_out4908_out1 XOR Logical_Operator_out4924_out1;

  Logical_Operator_out5933_out1 <= Logical_Operator_out4909_out1 XOR Logical_Operator_out4925_out1;

  Logical_Operator_out5934_out1 <= Logical_Operator_out4910_out1 XOR Logical_Operator_out4926_out1;

  Logical_Operator_out5935_out1 <= Logical_Operator_out4911_out1 XOR Logical_Operator_out4927_out1;

  Logical_Operator_out5936_out1 <= Logical_Operator_out4912_out1 XOR Logical_Operator_out4928_out1;

  Logical_Operator_out5937_out1 <= Logical_Operator_out3881_out1 XOR Logical_Operator_out3897_out1;

  Logical_Operator_out5938_out1 <= Logical_Operator_out3882_out1 XOR Logical_Operator_out3898_out1;

  Logical_Operator_out5939_out1 <= Logical_Operator_out3883_out1 XOR Logical_Operator_out3899_out1;

  Logical_Operator_out5940_out1 <= Logical_Operator_out3884_out1 XOR Logical_Operator_out3900_out1;

  Logical_Operator_out5941_out1 <= Logical_Operator_out3885_out1 XOR Logical_Operator_out3901_out1;

  Logical_Operator_out5942_out1 <= Logical_Operator_out3886_out1 XOR Logical_Operator_out3902_out1;

  Logical_Operator_out5943_out1 <= Logical_Operator_out3887_out1 XOR Logical_Operator_out3903_out1;

  Logical_Operator_out5944_out1 <= Logical_Operator_out3888_out1 XOR Logical_Operator_out3904_out1;

  Logical_Operator_out5945_out1 <= Logical_Operator_out2861_out1 XOR Logical_Operator_out2877_out1;

  Logical_Operator_out5946_out1 <= Logical_Operator_out2862_out1 XOR Logical_Operator_out2878_out1;

  Logical_Operator_out5947_out1 <= Logical_Operator_out2863_out1 XOR Logical_Operator_out2879_out1;

  Logical_Operator_out5948_out1 <= Logical_Operator_out2864_out1 XOR Logical_Operator_out2880_out1;

  Logical_Operator_out5949_out1 <= Logical_Operator_out1839_out1 XOR Logical_Operator_out1855_out1;

  Logical_Operator_out5950_out1 <= Logical_Operator_out1840_out1 XOR Logical_Operator_out1856_out1;

  Logical_Operator_out5951_out1 <= Logical_Operator_out816_out1 XOR Logical_Operator_out832_out1;

  Logical_Operator_out5952_out1 <= in1632 XOR in1664;

  Logical_Operator_out5953_out1 <= Logical_Operator_out4929_out1 XOR Logical_Operator_out4945_out1;

  Logical_Operator_out5954_out1 <= Logical_Operator_out4930_out1 XOR Logical_Operator_out4946_out1;

  Logical_Operator_out5955_out1 <= Logical_Operator_out4931_out1 XOR Logical_Operator_out4947_out1;

  Logical_Operator_out5956_out1 <= Logical_Operator_out4932_out1 XOR Logical_Operator_out4948_out1;

  Logical_Operator_out5957_out1 <= Logical_Operator_out4933_out1 XOR Logical_Operator_out4949_out1;

  Logical_Operator_out5958_out1 <= Logical_Operator_out4934_out1 XOR Logical_Operator_out4950_out1;

  Logical_Operator_out5959_out1 <= Logical_Operator_out4935_out1 XOR Logical_Operator_out4951_out1;

  Logical_Operator_out5960_out1 <= Logical_Operator_out4936_out1 XOR Logical_Operator_out4952_out1;

  Logical_Operator_out5961_out1 <= Logical_Operator_out4937_out1 XOR Logical_Operator_out4953_out1;

  Logical_Operator_out5962_out1 <= Logical_Operator_out4938_out1 XOR Logical_Operator_out4954_out1;

  Logical_Operator_out5963_out1 <= Logical_Operator_out4939_out1 XOR Logical_Operator_out4955_out1;

  Logical_Operator_out5964_out1 <= Logical_Operator_out4940_out1 XOR Logical_Operator_out4956_out1;

  Logical_Operator_out5965_out1 <= Logical_Operator_out4941_out1 XOR Logical_Operator_out4957_out1;

  Logical_Operator_out5966_out1 <= Logical_Operator_out4942_out1 XOR Logical_Operator_out4958_out1;

  Logical_Operator_out5967_out1 <= Logical_Operator_out4943_out1 XOR Logical_Operator_out4959_out1;

  Logical_Operator_out5968_out1 <= Logical_Operator_out4944_out1 XOR Logical_Operator_out4960_out1;

  Logical_Operator_out5969_out1 <= Logical_Operator_out3913_out1 XOR Logical_Operator_out3929_out1;

  Logical_Operator_out5970_out1 <= Logical_Operator_out3914_out1 XOR Logical_Operator_out3930_out1;

  Logical_Operator_out5971_out1 <= Logical_Operator_out3915_out1 XOR Logical_Operator_out3931_out1;

  Logical_Operator_out5972_out1 <= Logical_Operator_out3916_out1 XOR Logical_Operator_out3932_out1;

  Logical_Operator_out5973_out1 <= Logical_Operator_out3917_out1 XOR Logical_Operator_out3933_out1;

  Logical_Operator_out5974_out1 <= Logical_Operator_out3918_out1 XOR Logical_Operator_out3934_out1;

  Logical_Operator_out5975_out1 <= Logical_Operator_out3919_out1 XOR Logical_Operator_out3935_out1;

  Logical_Operator_out5976_out1 <= Logical_Operator_out3920_out1 XOR Logical_Operator_out3936_out1;

  Logical_Operator_out5977_out1 <= Logical_Operator_out2893_out1 XOR Logical_Operator_out2909_out1;

  Logical_Operator_out5978_out1 <= Logical_Operator_out2894_out1 XOR Logical_Operator_out2910_out1;

  Logical_Operator_out5979_out1 <= Logical_Operator_out2895_out1 XOR Logical_Operator_out2911_out1;

  Logical_Operator_out5980_out1 <= Logical_Operator_out2896_out1 XOR Logical_Operator_out2912_out1;

  Logical_Operator_out5981_out1 <= Logical_Operator_out1871_out1 XOR Logical_Operator_out1887_out1;

  Logical_Operator_out5982_out1 <= Logical_Operator_out1872_out1 XOR Logical_Operator_out1888_out1;

  Logical_Operator_out5983_out1 <= Logical_Operator_out848_out1 XOR Logical_Operator_out864_out1;

  Logical_Operator_out5984_out1 <= in1696 XOR in1728;

  Logical_Operator_out5985_out1 <= Logical_Operator_out4961_out1 XOR Logical_Operator_out4977_out1;

  Logical_Operator_out5986_out1 <= Logical_Operator_out4962_out1 XOR Logical_Operator_out4978_out1;

  Logical_Operator_out5987_out1 <= Logical_Operator_out4963_out1 XOR Logical_Operator_out4979_out1;

  Logical_Operator_out5988_out1 <= Logical_Operator_out4964_out1 XOR Logical_Operator_out4980_out1;

  Logical_Operator_out5989_out1 <= Logical_Operator_out4965_out1 XOR Logical_Operator_out4981_out1;

  Logical_Operator_out5990_out1 <= Logical_Operator_out4966_out1 XOR Logical_Operator_out4982_out1;

  Logical_Operator_out5991_out1 <= Logical_Operator_out4967_out1 XOR Logical_Operator_out4983_out1;

  Logical_Operator_out5992_out1 <= Logical_Operator_out4968_out1 XOR Logical_Operator_out4984_out1;

  Logical_Operator_out5993_out1 <= Logical_Operator_out4969_out1 XOR Logical_Operator_out4985_out1;

  Logical_Operator_out5994_out1 <= Logical_Operator_out4970_out1 XOR Logical_Operator_out4986_out1;

  Logical_Operator_out5995_out1 <= Logical_Operator_out4971_out1 XOR Logical_Operator_out4987_out1;

  Logical_Operator_out5996_out1 <= Logical_Operator_out4972_out1 XOR Logical_Operator_out4988_out1;

  Logical_Operator_out5997_out1 <= Logical_Operator_out4973_out1 XOR Logical_Operator_out4989_out1;

  Logical_Operator_out5998_out1 <= Logical_Operator_out4974_out1 XOR Logical_Operator_out4990_out1;

  Logical_Operator_out5999_out1 <= Logical_Operator_out4975_out1 XOR Logical_Operator_out4991_out1;

  Logical_Operator_out6000_out1 <= Logical_Operator_out4976_out1 XOR Logical_Operator_out4992_out1;

  Logical_Operator_out6001_out1 <= Logical_Operator_out3945_out1 XOR Logical_Operator_out3961_out1;

  Logical_Operator_out6002_out1 <= Logical_Operator_out3946_out1 XOR Logical_Operator_out3962_out1;

  Logical_Operator_out6003_out1 <= Logical_Operator_out3947_out1 XOR Logical_Operator_out3963_out1;

  Logical_Operator_out6004_out1 <= Logical_Operator_out3948_out1 XOR Logical_Operator_out3964_out1;

  Logical_Operator_out6005_out1 <= Logical_Operator_out3949_out1 XOR Logical_Operator_out3965_out1;

  Logical_Operator_out6006_out1 <= Logical_Operator_out3950_out1 XOR Logical_Operator_out3966_out1;

  Logical_Operator_out6007_out1 <= Logical_Operator_out3951_out1 XOR Logical_Operator_out3967_out1;

  Logical_Operator_out6008_out1 <= Logical_Operator_out3952_out1 XOR Logical_Operator_out3968_out1;

  Logical_Operator_out6009_out1 <= Logical_Operator_out2925_out1 XOR Logical_Operator_out2941_out1;

  Logical_Operator_out6010_out1 <= Logical_Operator_out2926_out1 XOR Logical_Operator_out2942_out1;

  Logical_Operator_out6011_out1 <= Logical_Operator_out2927_out1 XOR Logical_Operator_out2943_out1;

  Logical_Operator_out6012_out1 <= Logical_Operator_out2928_out1 XOR Logical_Operator_out2944_out1;

  Logical_Operator_out6013_out1 <= Logical_Operator_out1903_out1 XOR Logical_Operator_out1919_out1;

  Logical_Operator_out6014_out1 <= Logical_Operator_out1904_out1 XOR Logical_Operator_out1920_out1;

  Logical_Operator_out6015_out1 <= Logical_Operator_out880_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out6016_out1 <= in1760 XOR in1792;

  Logical_Operator_out6017_out1 <= Logical_Operator_out4993_out1 XOR Logical_Operator_out5009_out1;

  Logical_Operator_out6018_out1 <= Logical_Operator_out4994_out1 XOR Logical_Operator_out5010_out1;

  Logical_Operator_out6019_out1 <= Logical_Operator_out4995_out1 XOR Logical_Operator_out5011_out1;

  Logical_Operator_out6020_out1 <= Logical_Operator_out4996_out1 XOR Logical_Operator_out5012_out1;

  Logical_Operator_out6021_out1 <= Logical_Operator_out4997_out1 XOR Logical_Operator_out5013_out1;

  Logical_Operator_out6022_out1 <= Logical_Operator_out4998_out1 XOR Logical_Operator_out5014_out1;

  Logical_Operator_out6023_out1 <= Logical_Operator_out4999_out1 XOR Logical_Operator_out5015_out1;

  Logical_Operator_out6024_out1 <= Logical_Operator_out5000_out1 XOR Logical_Operator_out5016_out1;

  Logical_Operator_out6025_out1 <= Logical_Operator_out5001_out1 XOR Logical_Operator_out5017_out1;

  Logical_Operator_out6026_out1 <= Logical_Operator_out5002_out1 XOR Logical_Operator_out5018_out1;

  Logical_Operator_out6027_out1 <= Logical_Operator_out5003_out1 XOR Logical_Operator_out5019_out1;

  Logical_Operator_out6028_out1 <= Logical_Operator_out5004_out1 XOR Logical_Operator_out5020_out1;

  Logical_Operator_out6029_out1 <= Logical_Operator_out5005_out1 XOR Logical_Operator_out5021_out1;

  Logical_Operator_out6030_out1 <= Logical_Operator_out5006_out1 XOR Logical_Operator_out5022_out1;

  Logical_Operator_out6031_out1 <= Logical_Operator_out5007_out1 XOR Logical_Operator_out5023_out1;

  Logical_Operator_out6032_out1 <= Logical_Operator_out5008_out1 XOR Logical_Operator_out5024_out1;

  Logical_Operator_out6033_out1 <= Logical_Operator_out3977_out1 XOR Logical_Operator_out3993_out1;

  Logical_Operator_out6034_out1 <= Logical_Operator_out3978_out1 XOR Logical_Operator_out3994_out1;

  Logical_Operator_out6035_out1 <= Logical_Operator_out3979_out1 XOR Logical_Operator_out3995_out1;

  Logical_Operator_out6036_out1 <= Logical_Operator_out3980_out1 XOR Logical_Operator_out3996_out1;

  Logical_Operator_out6037_out1 <= Logical_Operator_out3981_out1 XOR Logical_Operator_out3997_out1;

  Logical_Operator_out6038_out1 <= Logical_Operator_out3982_out1 XOR Logical_Operator_out3998_out1;

  Logical_Operator_out6039_out1 <= Logical_Operator_out3983_out1 XOR Logical_Operator_out3999_out1;

  Logical_Operator_out6040_out1 <= Logical_Operator_out3984_out1 XOR Logical_Operator_out4000_out1;

  Logical_Operator_out6041_out1 <= Logical_Operator_out2957_out1 XOR Logical_Operator_out2973_out1;

  Logical_Operator_out6042_out1 <= Logical_Operator_out2958_out1 XOR Logical_Operator_out2974_out1;

  Logical_Operator_out6043_out1 <= Logical_Operator_out2959_out1 XOR Logical_Operator_out2975_out1;

  Logical_Operator_out6044_out1 <= Logical_Operator_out2960_out1 XOR Logical_Operator_out2976_out1;

  Logical_Operator_out6045_out1 <= Logical_Operator_out1935_out1 XOR Logical_Operator_out1951_out1;

  Logical_Operator_out6046_out1 <= Logical_Operator_out1936_out1 XOR Logical_Operator_out1952_out1;

  Logical_Operator_out6047_out1 <= Logical_Operator_out912_out1 XOR Logical_Operator_out928_out1;

  Logical_Operator_out6048_out1 <= in1824 XOR in1856;

  Logical_Operator_out6049_out1 <= Logical_Operator_out5025_out1 XOR Logical_Operator_out5041_out1;

  Logical_Operator_out6050_out1 <= Logical_Operator_out5026_out1 XOR Logical_Operator_out5042_out1;

  Logical_Operator_out6051_out1 <= Logical_Operator_out5027_out1 XOR Logical_Operator_out5043_out1;

  Logical_Operator_out6052_out1 <= Logical_Operator_out5028_out1 XOR Logical_Operator_out5044_out1;

  Logical_Operator_out6053_out1 <= Logical_Operator_out5029_out1 XOR Logical_Operator_out5045_out1;

  Logical_Operator_out6054_out1 <= Logical_Operator_out5030_out1 XOR Logical_Operator_out5046_out1;

  Logical_Operator_out6055_out1 <= Logical_Operator_out5031_out1 XOR Logical_Operator_out5047_out1;

  Logical_Operator_out6056_out1 <= Logical_Operator_out5032_out1 XOR Logical_Operator_out5048_out1;

  Logical_Operator_out6057_out1 <= Logical_Operator_out5033_out1 XOR Logical_Operator_out5049_out1;

  Logical_Operator_out6058_out1 <= Logical_Operator_out5034_out1 XOR Logical_Operator_out5050_out1;

  Logical_Operator_out6059_out1 <= Logical_Operator_out5035_out1 XOR Logical_Operator_out5051_out1;

  Logical_Operator_out6060_out1 <= Logical_Operator_out5036_out1 XOR Logical_Operator_out5052_out1;

  Logical_Operator_out6061_out1 <= Logical_Operator_out5037_out1 XOR Logical_Operator_out5053_out1;

  Logical_Operator_out6062_out1 <= Logical_Operator_out5038_out1 XOR Logical_Operator_out5054_out1;

  Logical_Operator_out6063_out1 <= Logical_Operator_out5039_out1 XOR Logical_Operator_out5055_out1;

  Logical_Operator_out6064_out1 <= Logical_Operator_out5040_out1 XOR Logical_Operator_out5056_out1;

  Logical_Operator_out6065_out1 <= Logical_Operator_out4009_out1 XOR Logical_Operator_out4025_out1;

  Logical_Operator_out6066_out1 <= Logical_Operator_out4010_out1 XOR Logical_Operator_out4026_out1;

  Logical_Operator_out6067_out1 <= Logical_Operator_out4011_out1 XOR Logical_Operator_out4027_out1;

  Logical_Operator_out6068_out1 <= Logical_Operator_out4012_out1 XOR Logical_Operator_out4028_out1;

  Logical_Operator_out6069_out1 <= Logical_Operator_out4013_out1 XOR Logical_Operator_out4029_out1;

  Logical_Operator_out6070_out1 <= Logical_Operator_out4014_out1 XOR Logical_Operator_out4030_out1;

  Logical_Operator_out6071_out1 <= Logical_Operator_out4015_out1 XOR Logical_Operator_out4031_out1;

  Logical_Operator_out6072_out1 <= Logical_Operator_out4016_out1 XOR Logical_Operator_out4032_out1;

  Logical_Operator_out6073_out1 <= Logical_Operator_out2989_out1 XOR Logical_Operator_out3005_out1;

  Logical_Operator_out6074_out1 <= Logical_Operator_out2990_out1 XOR Logical_Operator_out3006_out1;

  Logical_Operator_out6075_out1 <= Logical_Operator_out2991_out1 XOR Logical_Operator_out3007_out1;

  Logical_Operator_out6076_out1 <= Logical_Operator_out2992_out1 XOR Logical_Operator_out3008_out1;

  Logical_Operator_out6077_out1 <= Logical_Operator_out1967_out1 XOR Logical_Operator_out1983_out1;

  Logical_Operator_out6078_out1 <= Logical_Operator_out1968_out1 XOR Logical_Operator_out1984_out1;

  Logical_Operator_out6079_out1 <= Logical_Operator_out944_out1 XOR Logical_Operator_out960_out1;

  Logical_Operator_out6080_out1 <= in1888 XOR in1920;

  Logical_Operator_out6081_out1 <= Logical_Operator_out5057_out1 XOR Logical_Operator_out5073_out1;

  Logical_Operator_out6082_out1 <= Logical_Operator_out5058_out1 XOR Logical_Operator_out5074_out1;

  Logical_Operator_out6083_out1 <= Logical_Operator_out5059_out1 XOR Logical_Operator_out5075_out1;

  Logical_Operator_out6084_out1 <= Logical_Operator_out5060_out1 XOR Logical_Operator_out5076_out1;

  Logical_Operator_out6085_out1 <= Logical_Operator_out5061_out1 XOR Logical_Operator_out5077_out1;

  Logical_Operator_out6086_out1 <= Logical_Operator_out5062_out1 XOR Logical_Operator_out5078_out1;

  Logical_Operator_out6087_out1 <= Logical_Operator_out5063_out1 XOR Logical_Operator_out5079_out1;

  Logical_Operator_out6088_out1 <= Logical_Operator_out5064_out1 XOR Logical_Operator_out5080_out1;

  Logical_Operator_out6089_out1 <= Logical_Operator_out5065_out1 XOR Logical_Operator_out5081_out1;

  Logical_Operator_out6090_out1 <= Logical_Operator_out5066_out1 XOR Logical_Operator_out5082_out1;

  Logical_Operator_out6091_out1 <= Logical_Operator_out5067_out1 XOR Logical_Operator_out5083_out1;

  Logical_Operator_out6092_out1 <= Logical_Operator_out5068_out1 XOR Logical_Operator_out5084_out1;

  Logical_Operator_out6093_out1 <= Logical_Operator_out5069_out1 XOR Logical_Operator_out5085_out1;

  Logical_Operator_out6094_out1 <= Logical_Operator_out5070_out1 XOR Logical_Operator_out5086_out1;

  Logical_Operator_out6095_out1 <= Logical_Operator_out5071_out1 XOR Logical_Operator_out5087_out1;

  Logical_Operator_out6096_out1 <= Logical_Operator_out5072_out1 XOR Logical_Operator_out5088_out1;

  Logical_Operator_out6097_out1 <= Logical_Operator_out4041_out1 XOR Logical_Operator_out4057_out1;

  Logical_Operator_out6098_out1 <= Logical_Operator_out4042_out1 XOR Logical_Operator_out4058_out1;

  Logical_Operator_out6099_out1 <= Logical_Operator_out4043_out1 XOR Logical_Operator_out4059_out1;

  Logical_Operator_out6100_out1 <= Logical_Operator_out4044_out1 XOR Logical_Operator_out4060_out1;

  Logical_Operator_out6101_out1 <= Logical_Operator_out4045_out1 XOR Logical_Operator_out4061_out1;

  Logical_Operator_out6102_out1 <= Logical_Operator_out4046_out1 XOR Logical_Operator_out4062_out1;

  Logical_Operator_out6103_out1 <= Logical_Operator_out4047_out1 XOR Logical_Operator_out4063_out1;

  Logical_Operator_out6104_out1 <= Logical_Operator_out4048_out1 XOR Logical_Operator_out4064_out1;

  Logical_Operator_out6105_out1 <= Logical_Operator_out3021_out1 XOR Logical_Operator_out3037_out1;

  Logical_Operator_out6106_out1 <= Logical_Operator_out3022_out1 XOR Logical_Operator_out3038_out1;

  Logical_Operator_out6107_out1 <= Logical_Operator_out3023_out1 XOR Logical_Operator_out3039_out1;

  Logical_Operator_out6108_out1 <= Logical_Operator_out3024_out1 XOR Logical_Operator_out3040_out1;

  Logical_Operator_out6109_out1 <= Logical_Operator_out1999_out1 XOR Logical_Operator_out2015_out1;

  Logical_Operator_out6110_out1 <= Logical_Operator_out2000_out1 XOR Logical_Operator_out2016_out1;

  Logical_Operator_out6111_out1 <= Logical_Operator_out976_out1 XOR Logical_Operator_out992_out1;

  Logical_Operator_out6112_out1 <= in1952 XOR in1984;

  Logical_Operator_out6113_out1 <= Logical_Operator_out5089_out1 XOR Logical_Operator_out5105_out1;

  Logical_Operator_out6114_out1 <= Logical_Operator_out5090_out1 XOR Logical_Operator_out5106_out1;

  Logical_Operator_out6115_out1 <= Logical_Operator_out5091_out1 XOR Logical_Operator_out5107_out1;

  Logical_Operator_out6116_out1 <= Logical_Operator_out5092_out1 XOR Logical_Operator_out5108_out1;

  Logical_Operator_out6117_out1 <= Logical_Operator_out5093_out1 XOR Logical_Operator_out5109_out1;

  Logical_Operator_out6118_out1 <= Logical_Operator_out5094_out1 XOR Logical_Operator_out5110_out1;

  Logical_Operator_out6119_out1 <= Logical_Operator_out5095_out1 XOR Logical_Operator_out5111_out1;

  Logical_Operator_out6120_out1 <= Logical_Operator_out5096_out1 XOR Logical_Operator_out5112_out1;

  Logical_Operator_out6121_out1 <= Logical_Operator_out5097_out1 XOR Logical_Operator_out5113_out1;

  Logical_Operator_out6122_out1 <= Logical_Operator_out5098_out1 XOR Logical_Operator_out5114_out1;

  Logical_Operator_out6123_out1 <= Logical_Operator_out5099_out1 XOR Logical_Operator_out5115_out1;

  Logical_Operator_out6124_out1 <= Logical_Operator_out5100_out1 XOR Logical_Operator_out5116_out1;

  Logical_Operator_out6125_out1 <= Logical_Operator_out5101_out1 XOR Logical_Operator_out5117_out1;

  Logical_Operator_out6126_out1 <= Logical_Operator_out5102_out1 XOR Logical_Operator_out5118_out1;

  Logical_Operator_out6127_out1 <= Logical_Operator_out5103_out1 XOR Logical_Operator_out5119_out1;

  Logical_Operator_out6128_out1 <= Logical_Operator_out5104_out1 XOR Logical_Operator_out5120_out1;

  Logical_Operator_out6129_out1 <= Logical_Operator_out4073_out1 XOR Logical_Operator_out4089_out1;

  Logical_Operator_out6130_out1 <= Logical_Operator_out4074_out1 XOR Logical_Operator_out4090_out1;

  Logical_Operator_out6131_out1 <= Logical_Operator_out4075_out1 XOR Logical_Operator_out4091_out1;

  Logical_Operator_out6132_out1 <= Logical_Operator_out4076_out1 XOR Logical_Operator_out4092_out1;

  Logical_Operator_out6133_out1 <= Logical_Operator_out4077_out1 XOR Logical_Operator_out4093_out1;

  Logical_Operator_out6134_out1 <= Logical_Operator_out4078_out1 XOR Logical_Operator_out4094_out1;

  Logical_Operator_out6135_out1 <= Logical_Operator_out4079_out1 XOR Logical_Operator_out4095_out1;

  Logical_Operator_out6136_out1 <= Logical_Operator_out4080_out1 XOR Logical_Operator_out4096_out1;

  Logical_Operator_out6137_out1 <= Logical_Operator_out3053_out1 XOR Logical_Operator_out3069_out1;

  Logical_Operator_out6138_out1 <= Logical_Operator_out3054_out1 XOR Logical_Operator_out3070_out1;

  Logical_Operator_out6139_out1 <= Logical_Operator_out3055_out1 XOR Logical_Operator_out3071_out1;

  Logical_Operator_out6140_out1 <= Logical_Operator_out3056_out1 XOR Logical_Operator_out3072_out1;

  Logical_Operator_out6141_out1 <= Logical_Operator_out2031_out1 XOR Logical_Operator_out2047_out1;

  Logical_Operator_out6142_out1 <= Logical_Operator_out2032_out1 XOR Logical_Operator_out2048_out1;

  Logical_Operator_out6143_out1 <= Logical_Operator_out1008_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out6144_out1 <= in2016 XOR in2048;

  Logical_Operator_out6145_out1 <= Logical_Operator_out5121_out1 XOR Logical_Operator_out5153_out1;

  Logical_Operator_out6146_out1 <= Logical_Operator_out5122_out1 XOR Logical_Operator_out5154_out1;

  Logical_Operator_out6147_out1 <= Logical_Operator_out5123_out1 XOR Logical_Operator_out5155_out1;

  Logical_Operator_out6148_out1 <= Logical_Operator_out5124_out1 XOR Logical_Operator_out5156_out1;

  Logical_Operator_out6149_out1 <= Logical_Operator_out5125_out1 XOR Logical_Operator_out5157_out1;

  Logical_Operator_out6150_out1 <= Logical_Operator_out5126_out1 XOR Logical_Operator_out5158_out1;

  Logical_Operator_out6151_out1 <= Logical_Operator_out5127_out1 XOR Logical_Operator_out5159_out1;

  Logical_Operator_out6152_out1 <= Logical_Operator_out5128_out1 XOR Logical_Operator_out5160_out1;

  Logical_Operator_out6153_out1 <= Logical_Operator_out5129_out1 XOR Logical_Operator_out5161_out1;

  Logical_Operator_out6154_out1 <= Logical_Operator_out5130_out1 XOR Logical_Operator_out5162_out1;

  Logical_Operator_out6155_out1 <= Logical_Operator_out5131_out1 XOR Logical_Operator_out5163_out1;

  Logical_Operator_out6156_out1 <= Logical_Operator_out5132_out1 XOR Logical_Operator_out5164_out1;

  Logical_Operator_out6157_out1 <= Logical_Operator_out5133_out1 XOR Logical_Operator_out5165_out1;

  Logical_Operator_out6158_out1 <= Logical_Operator_out5134_out1 XOR Logical_Operator_out5166_out1;

  Logical_Operator_out6159_out1 <= Logical_Operator_out5135_out1 XOR Logical_Operator_out5167_out1;

  Logical_Operator_out6160_out1 <= Logical_Operator_out5136_out1 XOR Logical_Operator_out5168_out1;

  Logical_Operator_out6161_out1 <= Logical_Operator_out5137_out1 XOR Logical_Operator_out5169_out1;

  Logical_Operator_out6162_out1 <= Logical_Operator_out5138_out1 XOR Logical_Operator_out5170_out1;

  Logical_Operator_out6163_out1 <= Logical_Operator_out5139_out1 XOR Logical_Operator_out5171_out1;

  Logical_Operator_out6164_out1 <= Logical_Operator_out5140_out1 XOR Logical_Operator_out5172_out1;

  Logical_Operator_out6165_out1 <= Logical_Operator_out5141_out1 XOR Logical_Operator_out5173_out1;

  Logical_Operator_out6166_out1 <= Logical_Operator_out5142_out1 XOR Logical_Operator_out5174_out1;

  Logical_Operator_out6167_out1 <= Logical_Operator_out5143_out1 XOR Logical_Operator_out5175_out1;

  Logical_Operator_out6168_out1 <= Logical_Operator_out5144_out1 XOR Logical_Operator_out5176_out1;

  Logical_Operator_out6169_out1 <= Logical_Operator_out5145_out1 XOR Logical_Operator_out5177_out1;

  Logical_Operator_out6170_out1 <= Logical_Operator_out5146_out1 XOR Logical_Operator_out5178_out1;

  Logical_Operator_out6171_out1 <= Logical_Operator_out5147_out1 XOR Logical_Operator_out5179_out1;

  Logical_Operator_out6172_out1 <= Logical_Operator_out5148_out1 XOR Logical_Operator_out5180_out1;

  Logical_Operator_out6173_out1 <= Logical_Operator_out5149_out1 XOR Logical_Operator_out5181_out1;

  Logical_Operator_out6174_out1 <= Logical_Operator_out5150_out1 XOR Logical_Operator_out5182_out1;

  Logical_Operator_out6175_out1 <= Logical_Operator_out5151_out1 XOR Logical_Operator_out5183_out1;

  Logical_Operator_out6176_out1 <= Logical_Operator_out5152_out1 XOR Logical_Operator_out5184_out1;

  Logical_Operator_out6177_out1 <= Logical_Operator_out4113_out1 XOR Logical_Operator_out4145_out1;

  Logical_Operator_out6178_out1 <= Logical_Operator_out4114_out1 XOR Logical_Operator_out4146_out1;

  Logical_Operator_out6179_out1 <= Logical_Operator_out4115_out1 XOR Logical_Operator_out4147_out1;

  Logical_Operator_out6180_out1 <= Logical_Operator_out4116_out1 XOR Logical_Operator_out4148_out1;

  Logical_Operator_out6181_out1 <= Logical_Operator_out4117_out1 XOR Logical_Operator_out4149_out1;

  Logical_Operator_out6182_out1 <= Logical_Operator_out4118_out1 XOR Logical_Operator_out4150_out1;

  Logical_Operator_out6183_out1 <= Logical_Operator_out4119_out1 XOR Logical_Operator_out4151_out1;

  Logical_Operator_out6184_out1 <= Logical_Operator_out4120_out1 XOR Logical_Operator_out4152_out1;

  Logical_Operator_out6185_out1 <= Logical_Operator_out4121_out1 XOR Logical_Operator_out4153_out1;

  Logical_Operator_out6186_out1 <= Logical_Operator_out4122_out1 XOR Logical_Operator_out4154_out1;

  Logical_Operator_out6187_out1 <= Logical_Operator_out4123_out1 XOR Logical_Operator_out4155_out1;

  Logical_Operator_out6188_out1 <= Logical_Operator_out4124_out1 XOR Logical_Operator_out4156_out1;

  Logical_Operator_out6189_out1 <= Logical_Operator_out4125_out1 XOR Logical_Operator_out4157_out1;

  Logical_Operator_out6190_out1 <= Logical_Operator_out4126_out1 XOR Logical_Operator_out4158_out1;

  Logical_Operator_out6191_out1 <= Logical_Operator_out4127_out1 XOR Logical_Operator_out4159_out1;

  Logical_Operator_out6192_out1 <= Logical_Operator_out4128_out1 XOR Logical_Operator_out4160_out1;

  Logical_Operator_out6193_out1 <= Logical_Operator_out3097_out1 XOR Logical_Operator_out3129_out1;

  Logical_Operator_out6194_out1 <= Logical_Operator_out3098_out1 XOR Logical_Operator_out3130_out1;

  Logical_Operator_out6195_out1 <= Logical_Operator_out3099_out1 XOR Logical_Operator_out3131_out1;

  Logical_Operator_out6196_out1 <= Logical_Operator_out3100_out1 XOR Logical_Operator_out3132_out1;

  Logical_Operator_out6197_out1 <= Logical_Operator_out3101_out1 XOR Logical_Operator_out3133_out1;

  Logical_Operator_out6198_out1 <= Logical_Operator_out3102_out1 XOR Logical_Operator_out3134_out1;

  Logical_Operator_out6199_out1 <= Logical_Operator_out3103_out1 XOR Logical_Operator_out3135_out1;

  Logical_Operator_out6200_out1 <= Logical_Operator_out3104_out1 XOR Logical_Operator_out3136_out1;

  Logical_Operator_out6201_out1 <= Logical_Operator_out2077_out1 XOR Logical_Operator_out2109_out1;

  Logical_Operator_out6202_out1 <= Logical_Operator_out2078_out1 XOR Logical_Operator_out2110_out1;

  Logical_Operator_out6203_out1 <= Logical_Operator_out2079_out1 XOR Logical_Operator_out2111_out1;

  Logical_Operator_out6204_out1 <= Logical_Operator_out2080_out1 XOR Logical_Operator_out2112_out1;

  Logical_Operator_out6205_out1 <= Logical_Operator_out1055_out1 XOR Logical_Operator_out1087_out1;

  Logical_Operator_out6206_out1 <= Logical_Operator_out1056_out1 XOR Logical_Operator_out1088_out1;

  Logical_Operator_out6207_out1 <= Logical_Operator_out32_out1 XOR Logical_Operator_out64_out1;

  Logical_Operator_out6208_out1 <= in64 XOR in128;

  Logical_Operator_out6209_out1 <= Logical_Operator_out5185_out1 XOR Logical_Operator_out5217_out1;

  Logical_Operator_out6210_out1 <= Logical_Operator_out5186_out1 XOR Logical_Operator_out5218_out1;

  Logical_Operator_out6211_out1 <= Logical_Operator_out5187_out1 XOR Logical_Operator_out5219_out1;

  Logical_Operator_out6212_out1 <= Logical_Operator_out5188_out1 XOR Logical_Operator_out5220_out1;

  Logical_Operator_out6213_out1 <= Logical_Operator_out5189_out1 XOR Logical_Operator_out5221_out1;

  Logical_Operator_out6214_out1 <= Logical_Operator_out5190_out1 XOR Logical_Operator_out5222_out1;

  Logical_Operator_out6215_out1 <= Logical_Operator_out5191_out1 XOR Logical_Operator_out5223_out1;

  Logical_Operator_out6216_out1 <= Logical_Operator_out5192_out1 XOR Logical_Operator_out5224_out1;

  Logical_Operator_out6217_out1 <= Logical_Operator_out5193_out1 XOR Logical_Operator_out5225_out1;

  Logical_Operator_out6218_out1 <= Logical_Operator_out5194_out1 XOR Logical_Operator_out5226_out1;

  Logical_Operator_out6219_out1 <= Logical_Operator_out5195_out1 XOR Logical_Operator_out5227_out1;

  Logical_Operator_out6220_out1 <= Logical_Operator_out5196_out1 XOR Logical_Operator_out5228_out1;

  Logical_Operator_out6221_out1 <= Logical_Operator_out5197_out1 XOR Logical_Operator_out5229_out1;

  Logical_Operator_out6222_out1 <= Logical_Operator_out5198_out1 XOR Logical_Operator_out5230_out1;

  Logical_Operator_out6223_out1 <= Logical_Operator_out5199_out1 XOR Logical_Operator_out5231_out1;

  Logical_Operator_out6224_out1 <= Logical_Operator_out5200_out1 XOR Logical_Operator_out5232_out1;

  Logical_Operator_out6225_out1 <= Logical_Operator_out5201_out1 XOR Logical_Operator_out5233_out1;

  Logical_Operator_out6226_out1 <= Logical_Operator_out5202_out1 XOR Logical_Operator_out5234_out1;

  Logical_Operator_out6227_out1 <= Logical_Operator_out5203_out1 XOR Logical_Operator_out5235_out1;

  Logical_Operator_out6228_out1 <= Logical_Operator_out5204_out1 XOR Logical_Operator_out5236_out1;

  Logical_Operator_out6229_out1 <= Logical_Operator_out5205_out1 XOR Logical_Operator_out5237_out1;

  Logical_Operator_out6230_out1 <= Logical_Operator_out5206_out1 XOR Logical_Operator_out5238_out1;

  Logical_Operator_out6231_out1 <= Logical_Operator_out5207_out1 XOR Logical_Operator_out5239_out1;

  Logical_Operator_out6232_out1 <= Logical_Operator_out5208_out1 XOR Logical_Operator_out5240_out1;

  Logical_Operator_out6233_out1 <= Logical_Operator_out5209_out1 XOR Logical_Operator_out5241_out1;

  Logical_Operator_out6234_out1 <= Logical_Operator_out5210_out1 XOR Logical_Operator_out5242_out1;

  Logical_Operator_out6235_out1 <= Logical_Operator_out5211_out1 XOR Logical_Operator_out5243_out1;

  Logical_Operator_out6236_out1 <= Logical_Operator_out5212_out1 XOR Logical_Operator_out5244_out1;

  Logical_Operator_out6237_out1 <= Logical_Operator_out5213_out1 XOR Logical_Operator_out5245_out1;

  Logical_Operator_out6238_out1 <= Logical_Operator_out5214_out1 XOR Logical_Operator_out5246_out1;

  Logical_Operator_out6239_out1 <= Logical_Operator_out5215_out1 XOR Logical_Operator_out5247_out1;

  Logical_Operator_out6240_out1 <= Logical_Operator_out5216_out1 XOR Logical_Operator_out5248_out1;

  Logical_Operator_out6241_out1 <= Logical_Operator_out4177_out1 XOR Logical_Operator_out4209_out1;

  Logical_Operator_out6242_out1 <= Logical_Operator_out4178_out1 XOR Logical_Operator_out4210_out1;

  Logical_Operator_out6243_out1 <= Logical_Operator_out4179_out1 XOR Logical_Operator_out4211_out1;

  Logical_Operator_out6244_out1 <= Logical_Operator_out4180_out1 XOR Logical_Operator_out4212_out1;

  Logical_Operator_out6245_out1 <= Logical_Operator_out4181_out1 XOR Logical_Operator_out4213_out1;

  Logical_Operator_out6246_out1 <= Logical_Operator_out4182_out1 XOR Logical_Operator_out4214_out1;

  Logical_Operator_out6247_out1 <= Logical_Operator_out4183_out1 XOR Logical_Operator_out4215_out1;

  Logical_Operator_out6248_out1 <= Logical_Operator_out4184_out1 XOR Logical_Operator_out4216_out1;

  Logical_Operator_out6249_out1 <= Logical_Operator_out4185_out1 XOR Logical_Operator_out4217_out1;

  Logical_Operator_out6250_out1 <= Logical_Operator_out4186_out1 XOR Logical_Operator_out4218_out1;

  Logical_Operator_out6251_out1 <= Logical_Operator_out4187_out1 XOR Logical_Operator_out4219_out1;

  Logical_Operator_out6252_out1 <= Logical_Operator_out4188_out1 XOR Logical_Operator_out4220_out1;

  Logical_Operator_out6253_out1 <= Logical_Operator_out4189_out1 XOR Logical_Operator_out4221_out1;

  Logical_Operator_out6254_out1 <= Logical_Operator_out4190_out1 XOR Logical_Operator_out4222_out1;

  Logical_Operator_out6255_out1 <= Logical_Operator_out4191_out1 XOR Logical_Operator_out4223_out1;

  Logical_Operator_out6256_out1 <= Logical_Operator_out4192_out1 XOR Logical_Operator_out4224_out1;

  Logical_Operator_out6257_out1 <= Logical_Operator_out3161_out1 XOR Logical_Operator_out3193_out1;

  Logical_Operator_out6258_out1 <= Logical_Operator_out3162_out1 XOR Logical_Operator_out3194_out1;

  Logical_Operator_out6259_out1 <= Logical_Operator_out3163_out1 XOR Logical_Operator_out3195_out1;

  Logical_Operator_out6260_out1 <= Logical_Operator_out3164_out1 XOR Logical_Operator_out3196_out1;

  Logical_Operator_out6261_out1 <= Logical_Operator_out3165_out1 XOR Logical_Operator_out3197_out1;

  Logical_Operator_out6262_out1 <= Logical_Operator_out3166_out1 XOR Logical_Operator_out3198_out1;

  Logical_Operator_out6263_out1 <= Logical_Operator_out3167_out1 XOR Logical_Operator_out3199_out1;

  Logical_Operator_out6264_out1 <= Logical_Operator_out3168_out1 XOR Logical_Operator_out3200_out1;

  Logical_Operator_out6265_out1 <= Logical_Operator_out2141_out1 XOR Logical_Operator_out2173_out1;

  Logical_Operator_out6266_out1 <= Logical_Operator_out2142_out1 XOR Logical_Operator_out2174_out1;

  Logical_Operator_out6267_out1 <= Logical_Operator_out2143_out1 XOR Logical_Operator_out2175_out1;

  Logical_Operator_out6268_out1 <= Logical_Operator_out2144_out1 XOR Logical_Operator_out2176_out1;

  Logical_Operator_out6269_out1 <= Logical_Operator_out1119_out1 XOR Logical_Operator_out1151_out1;

  Logical_Operator_out6270_out1 <= Logical_Operator_out1120_out1 XOR Logical_Operator_out1152_out1;

  Logical_Operator_out6271_out1 <= Logical_Operator_out96_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out6272_out1 <= in192 XOR in256;

  Logical_Operator_out6273_out1 <= Logical_Operator_out5249_out1 XOR Logical_Operator_out5281_out1;

  Logical_Operator_out6274_out1 <= Logical_Operator_out5250_out1 XOR Logical_Operator_out5282_out1;

  Logical_Operator_out6275_out1 <= Logical_Operator_out5251_out1 XOR Logical_Operator_out5283_out1;

  Logical_Operator_out6276_out1 <= Logical_Operator_out5252_out1 XOR Logical_Operator_out5284_out1;

  Logical_Operator_out6277_out1 <= Logical_Operator_out5253_out1 XOR Logical_Operator_out5285_out1;

  Logical_Operator_out6278_out1 <= Logical_Operator_out5254_out1 XOR Logical_Operator_out5286_out1;

  Logical_Operator_out6279_out1 <= Logical_Operator_out5255_out1 XOR Logical_Operator_out5287_out1;

  Logical_Operator_out6280_out1 <= Logical_Operator_out5256_out1 XOR Logical_Operator_out5288_out1;

  Logical_Operator_out6281_out1 <= Logical_Operator_out5257_out1 XOR Logical_Operator_out5289_out1;

  Logical_Operator_out6282_out1 <= Logical_Operator_out5258_out1 XOR Logical_Operator_out5290_out1;

  Logical_Operator_out6283_out1 <= Logical_Operator_out5259_out1 XOR Logical_Operator_out5291_out1;

  Logical_Operator_out6284_out1 <= Logical_Operator_out5260_out1 XOR Logical_Operator_out5292_out1;

  Logical_Operator_out6285_out1 <= Logical_Operator_out5261_out1 XOR Logical_Operator_out5293_out1;

  Logical_Operator_out6286_out1 <= Logical_Operator_out5262_out1 XOR Logical_Operator_out5294_out1;

  Logical_Operator_out6287_out1 <= Logical_Operator_out5263_out1 XOR Logical_Operator_out5295_out1;

  Logical_Operator_out6288_out1 <= Logical_Operator_out5264_out1 XOR Logical_Operator_out5296_out1;

  Logical_Operator_out6289_out1 <= Logical_Operator_out5265_out1 XOR Logical_Operator_out5297_out1;

  Logical_Operator_out6290_out1 <= Logical_Operator_out5266_out1 XOR Logical_Operator_out5298_out1;

  Logical_Operator_out6291_out1 <= Logical_Operator_out5267_out1 XOR Logical_Operator_out5299_out1;

  Logical_Operator_out6292_out1 <= Logical_Operator_out5268_out1 XOR Logical_Operator_out5300_out1;

  Logical_Operator_out6293_out1 <= Logical_Operator_out5269_out1 XOR Logical_Operator_out5301_out1;

  Logical_Operator_out6294_out1 <= Logical_Operator_out5270_out1 XOR Logical_Operator_out5302_out1;

  Logical_Operator_out6295_out1 <= Logical_Operator_out5271_out1 XOR Logical_Operator_out5303_out1;

  Logical_Operator_out6296_out1 <= Logical_Operator_out5272_out1 XOR Logical_Operator_out5304_out1;

  Logical_Operator_out6297_out1 <= Logical_Operator_out5273_out1 XOR Logical_Operator_out5305_out1;

  Logical_Operator_out6298_out1 <= Logical_Operator_out5274_out1 XOR Logical_Operator_out5306_out1;

  Logical_Operator_out6299_out1 <= Logical_Operator_out5275_out1 XOR Logical_Operator_out5307_out1;

  Logical_Operator_out6300_out1 <= Logical_Operator_out5276_out1 XOR Logical_Operator_out5308_out1;

  Logical_Operator_out6301_out1 <= Logical_Operator_out5277_out1 XOR Logical_Operator_out5309_out1;

  Logical_Operator_out6302_out1 <= Logical_Operator_out5278_out1 XOR Logical_Operator_out5310_out1;

  Logical_Operator_out6303_out1 <= Logical_Operator_out5279_out1 XOR Logical_Operator_out5311_out1;

  Logical_Operator_out6304_out1 <= Logical_Operator_out5280_out1 XOR Logical_Operator_out5312_out1;

  Logical_Operator_out6305_out1 <= Logical_Operator_out4241_out1 XOR Logical_Operator_out4273_out1;

  Logical_Operator_out6306_out1 <= Logical_Operator_out4242_out1 XOR Logical_Operator_out4274_out1;

  Logical_Operator_out6307_out1 <= Logical_Operator_out4243_out1 XOR Logical_Operator_out4275_out1;

  Logical_Operator_out6308_out1 <= Logical_Operator_out4244_out1 XOR Logical_Operator_out4276_out1;

  Logical_Operator_out6309_out1 <= Logical_Operator_out4245_out1 XOR Logical_Operator_out4277_out1;

  Logical_Operator_out6310_out1 <= Logical_Operator_out4246_out1 XOR Logical_Operator_out4278_out1;

  Logical_Operator_out6311_out1 <= Logical_Operator_out4247_out1 XOR Logical_Operator_out4279_out1;

  Logical_Operator_out6312_out1 <= Logical_Operator_out4248_out1 XOR Logical_Operator_out4280_out1;

  Logical_Operator_out6313_out1 <= Logical_Operator_out4249_out1 XOR Logical_Operator_out4281_out1;

  Logical_Operator_out6314_out1 <= Logical_Operator_out4250_out1 XOR Logical_Operator_out4282_out1;

  Logical_Operator_out6315_out1 <= Logical_Operator_out4251_out1 XOR Logical_Operator_out4283_out1;

  Logical_Operator_out6316_out1 <= Logical_Operator_out4252_out1 XOR Logical_Operator_out4284_out1;

  Logical_Operator_out6317_out1 <= Logical_Operator_out4253_out1 XOR Logical_Operator_out4285_out1;

  Logical_Operator_out6318_out1 <= Logical_Operator_out4254_out1 XOR Logical_Operator_out4286_out1;

  Logical_Operator_out6319_out1 <= Logical_Operator_out4255_out1 XOR Logical_Operator_out4287_out1;

  Logical_Operator_out6320_out1 <= Logical_Operator_out4256_out1 XOR Logical_Operator_out4288_out1;

  Logical_Operator_out6321_out1 <= Logical_Operator_out3225_out1 XOR Logical_Operator_out3257_out1;

  Logical_Operator_out6322_out1 <= Logical_Operator_out3226_out1 XOR Logical_Operator_out3258_out1;

  Logical_Operator_out6323_out1 <= Logical_Operator_out3227_out1 XOR Logical_Operator_out3259_out1;

  Logical_Operator_out6324_out1 <= Logical_Operator_out3228_out1 XOR Logical_Operator_out3260_out1;

  Logical_Operator_out6325_out1 <= Logical_Operator_out3229_out1 XOR Logical_Operator_out3261_out1;

  Logical_Operator_out6326_out1 <= Logical_Operator_out3230_out1 XOR Logical_Operator_out3262_out1;

  Logical_Operator_out6327_out1 <= Logical_Operator_out3231_out1 XOR Logical_Operator_out3263_out1;

  Logical_Operator_out6328_out1 <= Logical_Operator_out3232_out1 XOR Logical_Operator_out3264_out1;

  Logical_Operator_out6329_out1 <= Logical_Operator_out2205_out1 XOR Logical_Operator_out2237_out1;

  Logical_Operator_out6330_out1 <= Logical_Operator_out2206_out1 XOR Logical_Operator_out2238_out1;

  Logical_Operator_out6331_out1 <= Logical_Operator_out2207_out1 XOR Logical_Operator_out2239_out1;

  Logical_Operator_out6332_out1 <= Logical_Operator_out2208_out1 XOR Logical_Operator_out2240_out1;

  Logical_Operator_out6333_out1 <= Logical_Operator_out1183_out1 XOR Logical_Operator_out1215_out1;

  Logical_Operator_out6334_out1 <= Logical_Operator_out1184_out1 XOR Logical_Operator_out1216_out1;

  Logical_Operator_out6335_out1 <= Logical_Operator_out160_out1 XOR Logical_Operator_out192_out1;

  Logical_Operator_out6336_out1 <= in320 XOR in384;

  Logical_Operator_out6337_out1 <= Logical_Operator_out5313_out1 XOR Logical_Operator_out5345_out1;

  Logical_Operator_out6338_out1 <= Logical_Operator_out5314_out1 XOR Logical_Operator_out5346_out1;

  Logical_Operator_out6339_out1 <= Logical_Operator_out5315_out1 XOR Logical_Operator_out5347_out1;

  Logical_Operator_out6340_out1 <= Logical_Operator_out5316_out1 XOR Logical_Operator_out5348_out1;

  Logical_Operator_out6341_out1 <= Logical_Operator_out5317_out1 XOR Logical_Operator_out5349_out1;

  Logical_Operator_out6342_out1 <= Logical_Operator_out5318_out1 XOR Logical_Operator_out5350_out1;

  Logical_Operator_out6343_out1 <= Logical_Operator_out5319_out1 XOR Logical_Operator_out5351_out1;

  Logical_Operator_out6344_out1 <= Logical_Operator_out5320_out1 XOR Logical_Operator_out5352_out1;

  Logical_Operator_out6345_out1 <= Logical_Operator_out5321_out1 XOR Logical_Operator_out5353_out1;

  Logical_Operator_out6346_out1 <= Logical_Operator_out5322_out1 XOR Logical_Operator_out5354_out1;

  Logical_Operator_out6347_out1 <= Logical_Operator_out5323_out1 XOR Logical_Operator_out5355_out1;

  Logical_Operator_out6348_out1 <= Logical_Operator_out5324_out1 XOR Logical_Operator_out5356_out1;

  Logical_Operator_out6349_out1 <= Logical_Operator_out5325_out1 XOR Logical_Operator_out5357_out1;

  Logical_Operator_out6350_out1 <= Logical_Operator_out5326_out1 XOR Logical_Operator_out5358_out1;

  Logical_Operator_out6351_out1 <= Logical_Operator_out5327_out1 XOR Logical_Operator_out5359_out1;

  Logical_Operator_out6352_out1 <= Logical_Operator_out5328_out1 XOR Logical_Operator_out5360_out1;

  Logical_Operator_out6353_out1 <= Logical_Operator_out5329_out1 XOR Logical_Operator_out5361_out1;

  Logical_Operator_out6354_out1 <= Logical_Operator_out5330_out1 XOR Logical_Operator_out5362_out1;

  Logical_Operator_out6355_out1 <= Logical_Operator_out5331_out1 XOR Logical_Operator_out5363_out1;

  Logical_Operator_out6356_out1 <= Logical_Operator_out5332_out1 XOR Logical_Operator_out5364_out1;

  Logical_Operator_out6357_out1 <= Logical_Operator_out5333_out1 XOR Logical_Operator_out5365_out1;

  Logical_Operator_out6358_out1 <= Logical_Operator_out5334_out1 XOR Logical_Operator_out5366_out1;

  Logical_Operator_out6359_out1 <= Logical_Operator_out5335_out1 XOR Logical_Operator_out5367_out1;

  Logical_Operator_out6360_out1 <= Logical_Operator_out5336_out1 XOR Logical_Operator_out5368_out1;

  Logical_Operator_out6361_out1 <= Logical_Operator_out5337_out1 XOR Logical_Operator_out5369_out1;

  Logical_Operator_out6362_out1 <= Logical_Operator_out5338_out1 XOR Logical_Operator_out5370_out1;

  Logical_Operator_out6363_out1 <= Logical_Operator_out5339_out1 XOR Logical_Operator_out5371_out1;

  Logical_Operator_out6364_out1 <= Logical_Operator_out5340_out1 XOR Logical_Operator_out5372_out1;

  Logical_Operator_out6365_out1 <= Logical_Operator_out5341_out1 XOR Logical_Operator_out5373_out1;

  Logical_Operator_out6366_out1 <= Logical_Operator_out5342_out1 XOR Logical_Operator_out5374_out1;

  Logical_Operator_out6367_out1 <= Logical_Operator_out5343_out1 XOR Logical_Operator_out5375_out1;

  Logical_Operator_out6368_out1 <= Logical_Operator_out5344_out1 XOR Logical_Operator_out5376_out1;

  Logical_Operator_out6369_out1 <= Logical_Operator_out4305_out1 XOR Logical_Operator_out4337_out1;

  Logical_Operator_out6370_out1 <= Logical_Operator_out4306_out1 XOR Logical_Operator_out4338_out1;

  Logical_Operator_out6371_out1 <= Logical_Operator_out4307_out1 XOR Logical_Operator_out4339_out1;

  Logical_Operator_out6372_out1 <= Logical_Operator_out4308_out1 XOR Logical_Operator_out4340_out1;

  Logical_Operator_out6373_out1 <= Logical_Operator_out4309_out1 XOR Logical_Operator_out4341_out1;

  Logical_Operator_out6374_out1 <= Logical_Operator_out4310_out1 XOR Logical_Operator_out4342_out1;

  Logical_Operator_out6375_out1 <= Logical_Operator_out4311_out1 XOR Logical_Operator_out4343_out1;

  Logical_Operator_out6376_out1 <= Logical_Operator_out4312_out1 XOR Logical_Operator_out4344_out1;

  Logical_Operator_out6377_out1 <= Logical_Operator_out4313_out1 XOR Logical_Operator_out4345_out1;

  Logical_Operator_out6378_out1 <= Logical_Operator_out4314_out1 XOR Logical_Operator_out4346_out1;

  Logical_Operator_out6379_out1 <= Logical_Operator_out4315_out1 XOR Logical_Operator_out4347_out1;

  Logical_Operator_out6380_out1 <= Logical_Operator_out4316_out1 XOR Logical_Operator_out4348_out1;

  Logical_Operator_out6381_out1 <= Logical_Operator_out4317_out1 XOR Logical_Operator_out4349_out1;

  Logical_Operator_out6382_out1 <= Logical_Operator_out4318_out1 XOR Logical_Operator_out4350_out1;

  Logical_Operator_out6383_out1 <= Logical_Operator_out4319_out1 XOR Logical_Operator_out4351_out1;

  Logical_Operator_out6384_out1 <= Logical_Operator_out4320_out1 XOR Logical_Operator_out4352_out1;

  Logical_Operator_out6385_out1 <= Logical_Operator_out3289_out1 XOR Logical_Operator_out3321_out1;

  Logical_Operator_out6386_out1 <= Logical_Operator_out3290_out1 XOR Logical_Operator_out3322_out1;

  Logical_Operator_out6387_out1 <= Logical_Operator_out3291_out1 XOR Logical_Operator_out3323_out1;

  Logical_Operator_out6388_out1 <= Logical_Operator_out3292_out1 XOR Logical_Operator_out3324_out1;

  Logical_Operator_out6389_out1 <= Logical_Operator_out3293_out1 XOR Logical_Operator_out3325_out1;

  Logical_Operator_out6390_out1 <= Logical_Operator_out3294_out1 XOR Logical_Operator_out3326_out1;

  Logical_Operator_out6391_out1 <= Logical_Operator_out3295_out1 XOR Logical_Operator_out3327_out1;

  Logical_Operator_out6392_out1 <= Logical_Operator_out3296_out1 XOR Logical_Operator_out3328_out1;

  Logical_Operator_out6393_out1 <= Logical_Operator_out2269_out1 XOR Logical_Operator_out2301_out1;

  Logical_Operator_out6394_out1 <= Logical_Operator_out2270_out1 XOR Logical_Operator_out2302_out1;

  Logical_Operator_out6395_out1 <= Logical_Operator_out2271_out1 XOR Logical_Operator_out2303_out1;

  Logical_Operator_out6396_out1 <= Logical_Operator_out2272_out1 XOR Logical_Operator_out2304_out1;

  Logical_Operator_out6397_out1 <= Logical_Operator_out1247_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out6398_out1 <= Logical_Operator_out1248_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out6399_out1 <= Logical_Operator_out224_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out6400_out1 <= in448 XOR in512;

  Logical_Operator_out6401_out1 <= Logical_Operator_out5377_out1 XOR Logical_Operator_out5409_out1;

  Logical_Operator_out6402_out1 <= Logical_Operator_out5378_out1 XOR Logical_Operator_out5410_out1;

  Logical_Operator_out6403_out1 <= Logical_Operator_out5379_out1 XOR Logical_Operator_out5411_out1;

  Logical_Operator_out6404_out1 <= Logical_Operator_out5380_out1 XOR Logical_Operator_out5412_out1;

  Logical_Operator_out6405_out1 <= Logical_Operator_out5381_out1 XOR Logical_Operator_out5413_out1;

  Logical_Operator_out6406_out1 <= Logical_Operator_out5382_out1 XOR Logical_Operator_out5414_out1;

  Logical_Operator_out6407_out1 <= Logical_Operator_out5383_out1 XOR Logical_Operator_out5415_out1;

  Logical_Operator_out6408_out1 <= Logical_Operator_out5384_out1 XOR Logical_Operator_out5416_out1;

  Logical_Operator_out6409_out1 <= Logical_Operator_out5385_out1 XOR Logical_Operator_out5417_out1;

  Logical_Operator_out6410_out1 <= Logical_Operator_out5386_out1 XOR Logical_Operator_out5418_out1;

  Logical_Operator_out6411_out1 <= Logical_Operator_out5387_out1 XOR Logical_Operator_out5419_out1;

  Logical_Operator_out6412_out1 <= Logical_Operator_out5388_out1 XOR Logical_Operator_out5420_out1;

  Logical_Operator_out6413_out1 <= Logical_Operator_out5389_out1 XOR Logical_Operator_out5421_out1;

  Logical_Operator_out6414_out1 <= Logical_Operator_out5390_out1 XOR Logical_Operator_out5422_out1;

  Logical_Operator_out6415_out1 <= Logical_Operator_out5391_out1 XOR Logical_Operator_out5423_out1;

  Logical_Operator_out6416_out1 <= Logical_Operator_out5392_out1 XOR Logical_Operator_out5424_out1;

  Logical_Operator_out6417_out1 <= Logical_Operator_out5393_out1 XOR Logical_Operator_out5425_out1;

  Logical_Operator_out6418_out1 <= Logical_Operator_out5394_out1 XOR Logical_Operator_out5426_out1;

  Logical_Operator_out6419_out1 <= Logical_Operator_out5395_out1 XOR Logical_Operator_out5427_out1;

  Logical_Operator_out6420_out1 <= Logical_Operator_out5396_out1 XOR Logical_Operator_out5428_out1;

  Logical_Operator_out6421_out1 <= Logical_Operator_out5397_out1 XOR Logical_Operator_out5429_out1;

  Logical_Operator_out6422_out1 <= Logical_Operator_out5398_out1 XOR Logical_Operator_out5430_out1;

  Logical_Operator_out6423_out1 <= Logical_Operator_out5399_out1 XOR Logical_Operator_out5431_out1;

  Logical_Operator_out6424_out1 <= Logical_Operator_out5400_out1 XOR Logical_Operator_out5432_out1;

  Logical_Operator_out6425_out1 <= Logical_Operator_out5401_out1 XOR Logical_Operator_out5433_out1;

  Logical_Operator_out6426_out1 <= Logical_Operator_out5402_out1 XOR Logical_Operator_out5434_out1;

  Logical_Operator_out6427_out1 <= Logical_Operator_out5403_out1 XOR Logical_Operator_out5435_out1;

  Logical_Operator_out6428_out1 <= Logical_Operator_out5404_out1 XOR Logical_Operator_out5436_out1;

  Logical_Operator_out6429_out1 <= Logical_Operator_out5405_out1 XOR Logical_Operator_out5437_out1;

  Logical_Operator_out6430_out1 <= Logical_Operator_out5406_out1 XOR Logical_Operator_out5438_out1;

  Logical_Operator_out6431_out1 <= Logical_Operator_out5407_out1 XOR Logical_Operator_out5439_out1;

  Logical_Operator_out6432_out1 <= Logical_Operator_out5408_out1 XOR Logical_Operator_out5440_out1;

  Logical_Operator_out6433_out1 <= Logical_Operator_out4369_out1 XOR Logical_Operator_out4401_out1;

  Logical_Operator_out6434_out1 <= Logical_Operator_out4370_out1 XOR Logical_Operator_out4402_out1;

  Logical_Operator_out6435_out1 <= Logical_Operator_out4371_out1 XOR Logical_Operator_out4403_out1;

  Logical_Operator_out6436_out1 <= Logical_Operator_out4372_out1 XOR Logical_Operator_out4404_out1;

  Logical_Operator_out6437_out1 <= Logical_Operator_out4373_out1 XOR Logical_Operator_out4405_out1;

  Logical_Operator_out6438_out1 <= Logical_Operator_out4374_out1 XOR Logical_Operator_out4406_out1;

  Logical_Operator_out6439_out1 <= Logical_Operator_out4375_out1 XOR Logical_Operator_out4407_out1;

  Logical_Operator_out6440_out1 <= Logical_Operator_out4376_out1 XOR Logical_Operator_out4408_out1;

  Logical_Operator_out6441_out1 <= Logical_Operator_out4377_out1 XOR Logical_Operator_out4409_out1;

  Logical_Operator_out6442_out1 <= Logical_Operator_out4378_out1 XOR Logical_Operator_out4410_out1;

  Logical_Operator_out6443_out1 <= Logical_Operator_out4379_out1 XOR Logical_Operator_out4411_out1;

  Logical_Operator_out6444_out1 <= Logical_Operator_out4380_out1 XOR Logical_Operator_out4412_out1;

  Logical_Operator_out6445_out1 <= Logical_Operator_out4381_out1 XOR Logical_Operator_out4413_out1;

  Logical_Operator_out6446_out1 <= Logical_Operator_out4382_out1 XOR Logical_Operator_out4414_out1;

  Logical_Operator_out6447_out1 <= Logical_Operator_out4383_out1 XOR Logical_Operator_out4415_out1;

  Logical_Operator_out6448_out1 <= Logical_Operator_out4384_out1 XOR Logical_Operator_out4416_out1;

  Logical_Operator_out6449_out1 <= Logical_Operator_out3353_out1 XOR Logical_Operator_out3385_out1;

  Logical_Operator_out6450_out1 <= Logical_Operator_out3354_out1 XOR Logical_Operator_out3386_out1;

  Logical_Operator_out6451_out1 <= Logical_Operator_out3355_out1 XOR Logical_Operator_out3387_out1;

  Logical_Operator_out6452_out1 <= Logical_Operator_out3356_out1 XOR Logical_Operator_out3388_out1;

  Logical_Operator_out6453_out1 <= Logical_Operator_out3357_out1 XOR Logical_Operator_out3389_out1;

  Logical_Operator_out6454_out1 <= Logical_Operator_out3358_out1 XOR Logical_Operator_out3390_out1;

  Logical_Operator_out6455_out1 <= Logical_Operator_out3359_out1 XOR Logical_Operator_out3391_out1;

  Logical_Operator_out6456_out1 <= Logical_Operator_out3360_out1 XOR Logical_Operator_out3392_out1;

  Logical_Operator_out6457_out1 <= Logical_Operator_out2333_out1 XOR Logical_Operator_out2365_out1;

  Logical_Operator_out6458_out1 <= Logical_Operator_out2334_out1 XOR Logical_Operator_out2366_out1;

  Logical_Operator_out6459_out1 <= Logical_Operator_out2335_out1 XOR Logical_Operator_out2367_out1;

  Logical_Operator_out6460_out1 <= Logical_Operator_out2336_out1 XOR Logical_Operator_out2368_out1;

  Logical_Operator_out6461_out1 <= Logical_Operator_out1311_out1 XOR Logical_Operator_out1343_out1;

  Logical_Operator_out6462_out1 <= Logical_Operator_out1312_out1 XOR Logical_Operator_out1344_out1;

  Logical_Operator_out6463_out1 <= Logical_Operator_out288_out1 XOR Logical_Operator_out320_out1;

  Logical_Operator_out6464_out1 <= in576 XOR in640;

  Logical_Operator_out6465_out1 <= Logical_Operator_out5441_out1 XOR Logical_Operator_out5473_out1;

  Logical_Operator_out6466_out1 <= Logical_Operator_out5442_out1 XOR Logical_Operator_out5474_out1;

  Logical_Operator_out6467_out1 <= Logical_Operator_out5443_out1 XOR Logical_Operator_out5475_out1;

  Logical_Operator_out6468_out1 <= Logical_Operator_out5444_out1 XOR Logical_Operator_out5476_out1;

  Logical_Operator_out6469_out1 <= Logical_Operator_out5445_out1 XOR Logical_Operator_out5477_out1;

  Logical_Operator_out6470_out1 <= Logical_Operator_out5446_out1 XOR Logical_Operator_out5478_out1;

  Logical_Operator_out6471_out1 <= Logical_Operator_out5447_out1 XOR Logical_Operator_out5479_out1;

  Logical_Operator_out6472_out1 <= Logical_Operator_out5448_out1 XOR Logical_Operator_out5480_out1;

  Logical_Operator_out6473_out1 <= Logical_Operator_out5449_out1 XOR Logical_Operator_out5481_out1;

  Logical_Operator_out6474_out1 <= Logical_Operator_out5450_out1 XOR Logical_Operator_out5482_out1;

  Logical_Operator_out6475_out1 <= Logical_Operator_out5451_out1 XOR Logical_Operator_out5483_out1;

  Logical_Operator_out6476_out1 <= Logical_Operator_out5452_out1 XOR Logical_Operator_out5484_out1;

  Logical_Operator_out6477_out1 <= Logical_Operator_out5453_out1 XOR Logical_Operator_out5485_out1;

  Logical_Operator_out6478_out1 <= Logical_Operator_out5454_out1 XOR Logical_Operator_out5486_out1;

  Logical_Operator_out6479_out1 <= Logical_Operator_out5455_out1 XOR Logical_Operator_out5487_out1;

  Logical_Operator_out6480_out1 <= Logical_Operator_out5456_out1 XOR Logical_Operator_out5488_out1;

  Logical_Operator_out6481_out1 <= Logical_Operator_out5457_out1 XOR Logical_Operator_out5489_out1;

  Logical_Operator_out6482_out1 <= Logical_Operator_out5458_out1 XOR Logical_Operator_out5490_out1;

  Logical_Operator_out6483_out1 <= Logical_Operator_out5459_out1 XOR Logical_Operator_out5491_out1;

  Logical_Operator_out6484_out1 <= Logical_Operator_out5460_out1 XOR Logical_Operator_out5492_out1;

  Logical_Operator_out6485_out1 <= Logical_Operator_out5461_out1 XOR Logical_Operator_out5493_out1;

  Logical_Operator_out6486_out1 <= Logical_Operator_out5462_out1 XOR Logical_Operator_out5494_out1;

  Logical_Operator_out6487_out1 <= Logical_Operator_out5463_out1 XOR Logical_Operator_out5495_out1;

  Logical_Operator_out6488_out1 <= Logical_Operator_out5464_out1 XOR Logical_Operator_out5496_out1;

  Logical_Operator_out6489_out1 <= Logical_Operator_out5465_out1 XOR Logical_Operator_out5497_out1;

  Logical_Operator_out6490_out1 <= Logical_Operator_out5466_out1 XOR Logical_Operator_out5498_out1;

  Logical_Operator_out6491_out1 <= Logical_Operator_out5467_out1 XOR Logical_Operator_out5499_out1;

  Logical_Operator_out6492_out1 <= Logical_Operator_out5468_out1 XOR Logical_Operator_out5500_out1;

  Logical_Operator_out6493_out1 <= Logical_Operator_out5469_out1 XOR Logical_Operator_out5501_out1;

  Logical_Operator_out6494_out1 <= Logical_Operator_out5470_out1 XOR Logical_Operator_out5502_out1;

  Logical_Operator_out6495_out1 <= Logical_Operator_out5471_out1 XOR Logical_Operator_out5503_out1;

  Logical_Operator_out6496_out1 <= Logical_Operator_out5472_out1 XOR Logical_Operator_out5504_out1;

  Logical_Operator_out6497_out1 <= Logical_Operator_out4433_out1 XOR Logical_Operator_out4465_out1;

  Logical_Operator_out6498_out1 <= Logical_Operator_out4434_out1 XOR Logical_Operator_out4466_out1;

  Logical_Operator_out6499_out1 <= Logical_Operator_out4435_out1 XOR Logical_Operator_out4467_out1;

  Logical_Operator_out6500_out1 <= Logical_Operator_out4436_out1 XOR Logical_Operator_out4468_out1;

  Logical_Operator_out6501_out1 <= Logical_Operator_out4437_out1 XOR Logical_Operator_out4469_out1;

  Logical_Operator_out6502_out1 <= Logical_Operator_out4438_out1 XOR Logical_Operator_out4470_out1;

  Logical_Operator_out6503_out1 <= Logical_Operator_out4439_out1 XOR Logical_Operator_out4471_out1;

  Logical_Operator_out6504_out1 <= Logical_Operator_out4440_out1 XOR Logical_Operator_out4472_out1;

  Logical_Operator_out6505_out1 <= Logical_Operator_out4441_out1 XOR Logical_Operator_out4473_out1;

  Logical_Operator_out6506_out1 <= Logical_Operator_out4442_out1 XOR Logical_Operator_out4474_out1;

  Logical_Operator_out6507_out1 <= Logical_Operator_out4443_out1 XOR Logical_Operator_out4475_out1;

  Logical_Operator_out6508_out1 <= Logical_Operator_out4444_out1 XOR Logical_Operator_out4476_out1;

  Logical_Operator_out6509_out1 <= Logical_Operator_out4445_out1 XOR Logical_Operator_out4477_out1;

  Logical_Operator_out6510_out1 <= Logical_Operator_out4446_out1 XOR Logical_Operator_out4478_out1;

  Logical_Operator_out6511_out1 <= Logical_Operator_out4447_out1 XOR Logical_Operator_out4479_out1;

  Logical_Operator_out6512_out1 <= Logical_Operator_out4448_out1 XOR Logical_Operator_out4480_out1;

  Logical_Operator_out6513_out1 <= Logical_Operator_out3417_out1 XOR Logical_Operator_out3449_out1;

  Logical_Operator_out6514_out1 <= Logical_Operator_out3418_out1 XOR Logical_Operator_out3450_out1;

  Logical_Operator_out6515_out1 <= Logical_Operator_out3419_out1 XOR Logical_Operator_out3451_out1;

  Logical_Operator_out6516_out1 <= Logical_Operator_out3420_out1 XOR Logical_Operator_out3452_out1;

  Logical_Operator_out6517_out1 <= Logical_Operator_out3421_out1 XOR Logical_Operator_out3453_out1;

  Logical_Operator_out6518_out1 <= Logical_Operator_out3422_out1 XOR Logical_Operator_out3454_out1;

  Logical_Operator_out6519_out1 <= Logical_Operator_out3423_out1 XOR Logical_Operator_out3455_out1;

  Logical_Operator_out6520_out1 <= Logical_Operator_out3424_out1 XOR Logical_Operator_out3456_out1;

  Logical_Operator_out6521_out1 <= Logical_Operator_out2397_out1 XOR Logical_Operator_out2429_out1;

  Logical_Operator_out6522_out1 <= Logical_Operator_out2398_out1 XOR Logical_Operator_out2430_out1;

  Logical_Operator_out6523_out1 <= Logical_Operator_out2399_out1 XOR Logical_Operator_out2431_out1;

  Logical_Operator_out6524_out1 <= Logical_Operator_out2400_out1 XOR Logical_Operator_out2432_out1;

  Logical_Operator_out6525_out1 <= Logical_Operator_out1375_out1 XOR Logical_Operator_out1407_out1;

  Logical_Operator_out6526_out1 <= Logical_Operator_out1376_out1 XOR Logical_Operator_out1408_out1;

  Logical_Operator_out6527_out1 <= Logical_Operator_out352_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out6528_out1 <= in704 XOR in768;

  Logical_Operator_out6529_out1 <= Logical_Operator_out5505_out1 XOR Logical_Operator_out5537_out1;

  Logical_Operator_out6530_out1 <= Logical_Operator_out5506_out1 XOR Logical_Operator_out5538_out1;

  Logical_Operator_out6531_out1 <= Logical_Operator_out5507_out1 XOR Logical_Operator_out5539_out1;

  Logical_Operator_out6532_out1 <= Logical_Operator_out5508_out1 XOR Logical_Operator_out5540_out1;

  Logical_Operator_out6533_out1 <= Logical_Operator_out5509_out1 XOR Logical_Operator_out5541_out1;

  Logical_Operator_out6534_out1 <= Logical_Operator_out5510_out1 XOR Logical_Operator_out5542_out1;

  Logical_Operator_out6535_out1 <= Logical_Operator_out5511_out1 XOR Logical_Operator_out5543_out1;

  Logical_Operator_out6536_out1 <= Logical_Operator_out5512_out1 XOR Logical_Operator_out5544_out1;

  Logical_Operator_out6537_out1 <= Logical_Operator_out5513_out1 XOR Logical_Operator_out5545_out1;

  Logical_Operator_out6538_out1 <= Logical_Operator_out5514_out1 XOR Logical_Operator_out5546_out1;

  Logical_Operator_out6539_out1 <= Logical_Operator_out5515_out1 XOR Logical_Operator_out5547_out1;

  Logical_Operator_out6540_out1 <= Logical_Operator_out5516_out1 XOR Logical_Operator_out5548_out1;

  Logical_Operator_out6541_out1 <= Logical_Operator_out5517_out1 XOR Logical_Operator_out5549_out1;

  Logical_Operator_out6542_out1 <= Logical_Operator_out5518_out1 XOR Logical_Operator_out5550_out1;

  Logical_Operator_out6543_out1 <= Logical_Operator_out5519_out1 XOR Logical_Operator_out5551_out1;

  Logical_Operator_out6544_out1 <= Logical_Operator_out5520_out1 XOR Logical_Operator_out5552_out1;

  Logical_Operator_out6545_out1 <= Logical_Operator_out5521_out1 XOR Logical_Operator_out5553_out1;

  Logical_Operator_out6546_out1 <= Logical_Operator_out5522_out1 XOR Logical_Operator_out5554_out1;

  Logical_Operator_out6547_out1 <= Logical_Operator_out5523_out1 XOR Logical_Operator_out5555_out1;

  Logical_Operator_out6548_out1 <= Logical_Operator_out5524_out1 XOR Logical_Operator_out5556_out1;

  Logical_Operator_out6549_out1 <= Logical_Operator_out5525_out1 XOR Logical_Operator_out5557_out1;

  Logical_Operator_out6550_out1 <= Logical_Operator_out5526_out1 XOR Logical_Operator_out5558_out1;

  Logical_Operator_out6551_out1 <= Logical_Operator_out5527_out1 XOR Logical_Operator_out5559_out1;

  Logical_Operator_out6552_out1 <= Logical_Operator_out5528_out1 XOR Logical_Operator_out5560_out1;

  Logical_Operator_out6553_out1 <= Logical_Operator_out5529_out1 XOR Logical_Operator_out5561_out1;

  Logical_Operator_out6554_out1 <= Logical_Operator_out5530_out1 XOR Logical_Operator_out5562_out1;

  Logical_Operator_out6555_out1 <= Logical_Operator_out5531_out1 XOR Logical_Operator_out5563_out1;

  Logical_Operator_out6556_out1 <= Logical_Operator_out5532_out1 XOR Logical_Operator_out5564_out1;

  Logical_Operator_out6557_out1 <= Logical_Operator_out5533_out1 XOR Logical_Operator_out5565_out1;

  Logical_Operator_out6558_out1 <= Logical_Operator_out5534_out1 XOR Logical_Operator_out5566_out1;

  Logical_Operator_out6559_out1 <= Logical_Operator_out5535_out1 XOR Logical_Operator_out5567_out1;

  Logical_Operator_out6560_out1 <= Logical_Operator_out5536_out1 XOR Logical_Operator_out5568_out1;

  Logical_Operator_out6561_out1 <= Logical_Operator_out4497_out1 XOR Logical_Operator_out4529_out1;

  Logical_Operator_out6562_out1 <= Logical_Operator_out4498_out1 XOR Logical_Operator_out4530_out1;

  Logical_Operator_out6563_out1 <= Logical_Operator_out4499_out1 XOR Logical_Operator_out4531_out1;

  Logical_Operator_out6564_out1 <= Logical_Operator_out4500_out1 XOR Logical_Operator_out4532_out1;

  Logical_Operator_out6565_out1 <= Logical_Operator_out4501_out1 XOR Logical_Operator_out4533_out1;

  Logical_Operator_out6566_out1 <= Logical_Operator_out4502_out1 XOR Logical_Operator_out4534_out1;

  Logical_Operator_out6567_out1 <= Logical_Operator_out4503_out1 XOR Logical_Operator_out4535_out1;

  Logical_Operator_out6568_out1 <= Logical_Operator_out4504_out1 XOR Logical_Operator_out4536_out1;

  Logical_Operator_out6569_out1 <= Logical_Operator_out4505_out1 XOR Logical_Operator_out4537_out1;

  Logical_Operator_out6570_out1 <= Logical_Operator_out4506_out1 XOR Logical_Operator_out4538_out1;

  Logical_Operator_out6571_out1 <= Logical_Operator_out4507_out1 XOR Logical_Operator_out4539_out1;

  Logical_Operator_out6572_out1 <= Logical_Operator_out4508_out1 XOR Logical_Operator_out4540_out1;

  Logical_Operator_out6573_out1 <= Logical_Operator_out4509_out1 XOR Logical_Operator_out4541_out1;

  Logical_Operator_out6574_out1 <= Logical_Operator_out4510_out1 XOR Logical_Operator_out4542_out1;

  Logical_Operator_out6575_out1 <= Logical_Operator_out4511_out1 XOR Logical_Operator_out4543_out1;

  Logical_Operator_out6576_out1 <= Logical_Operator_out4512_out1 XOR Logical_Operator_out4544_out1;

  Logical_Operator_out6577_out1 <= Logical_Operator_out3481_out1 XOR Logical_Operator_out3513_out1;

  Logical_Operator_out6578_out1 <= Logical_Operator_out3482_out1 XOR Logical_Operator_out3514_out1;

  Logical_Operator_out6579_out1 <= Logical_Operator_out3483_out1 XOR Logical_Operator_out3515_out1;

  Logical_Operator_out6580_out1 <= Logical_Operator_out3484_out1 XOR Logical_Operator_out3516_out1;

  Logical_Operator_out6581_out1 <= Logical_Operator_out3485_out1 XOR Logical_Operator_out3517_out1;

  Logical_Operator_out6582_out1 <= Logical_Operator_out3486_out1 XOR Logical_Operator_out3518_out1;

  Logical_Operator_out6583_out1 <= Logical_Operator_out3487_out1 XOR Logical_Operator_out3519_out1;

  Logical_Operator_out6584_out1 <= Logical_Operator_out3488_out1 XOR Logical_Operator_out3520_out1;

  Logical_Operator_out6585_out1 <= Logical_Operator_out2461_out1 XOR Logical_Operator_out2493_out1;

  Logical_Operator_out6586_out1 <= Logical_Operator_out2462_out1 XOR Logical_Operator_out2494_out1;

  Logical_Operator_out6587_out1 <= Logical_Operator_out2463_out1 XOR Logical_Operator_out2495_out1;

  Logical_Operator_out6588_out1 <= Logical_Operator_out2464_out1 XOR Logical_Operator_out2496_out1;

  Logical_Operator_out6589_out1 <= Logical_Operator_out1439_out1 XOR Logical_Operator_out1471_out1;

  Logical_Operator_out6590_out1 <= Logical_Operator_out1440_out1 XOR Logical_Operator_out1472_out1;

  Logical_Operator_out6591_out1 <= Logical_Operator_out416_out1 XOR Logical_Operator_out448_out1;

  Logical_Operator_out6592_out1 <= in832 XOR in896;

  Logical_Operator_out6593_out1 <= Logical_Operator_out5569_out1 XOR Logical_Operator_out5601_out1;

  Logical_Operator_out6594_out1 <= Logical_Operator_out5570_out1 XOR Logical_Operator_out5602_out1;

  Logical_Operator_out6595_out1 <= Logical_Operator_out5571_out1 XOR Logical_Operator_out5603_out1;

  Logical_Operator_out6596_out1 <= Logical_Operator_out5572_out1 XOR Logical_Operator_out5604_out1;

  Logical_Operator_out6597_out1 <= Logical_Operator_out5573_out1 XOR Logical_Operator_out5605_out1;

  Logical_Operator_out6598_out1 <= Logical_Operator_out5574_out1 XOR Logical_Operator_out5606_out1;

  Logical_Operator_out6599_out1 <= Logical_Operator_out5575_out1 XOR Logical_Operator_out5607_out1;

  Logical_Operator_out6600_out1 <= Logical_Operator_out5576_out1 XOR Logical_Operator_out5608_out1;

  Logical_Operator_out6601_out1 <= Logical_Operator_out5577_out1 XOR Logical_Operator_out5609_out1;

  Logical_Operator_out6602_out1 <= Logical_Operator_out5578_out1 XOR Logical_Operator_out5610_out1;

  Logical_Operator_out6603_out1 <= Logical_Operator_out5579_out1 XOR Logical_Operator_out5611_out1;

  Logical_Operator_out6604_out1 <= Logical_Operator_out5580_out1 XOR Logical_Operator_out5612_out1;

  Logical_Operator_out6605_out1 <= Logical_Operator_out5581_out1 XOR Logical_Operator_out5613_out1;

  Logical_Operator_out6606_out1 <= Logical_Operator_out5582_out1 XOR Logical_Operator_out5614_out1;

  Logical_Operator_out6607_out1 <= Logical_Operator_out5583_out1 XOR Logical_Operator_out5615_out1;

  Logical_Operator_out6608_out1 <= Logical_Operator_out5584_out1 XOR Logical_Operator_out5616_out1;

  Logical_Operator_out6609_out1 <= Logical_Operator_out5585_out1 XOR Logical_Operator_out5617_out1;

  Logical_Operator_out6610_out1 <= Logical_Operator_out5586_out1 XOR Logical_Operator_out5618_out1;

  Logical_Operator_out6611_out1 <= Logical_Operator_out5587_out1 XOR Logical_Operator_out5619_out1;

  Logical_Operator_out6612_out1 <= Logical_Operator_out5588_out1 XOR Logical_Operator_out5620_out1;

  Logical_Operator_out6613_out1 <= Logical_Operator_out5589_out1 XOR Logical_Operator_out5621_out1;

  Logical_Operator_out6614_out1 <= Logical_Operator_out5590_out1 XOR Logical_Operator_out5622_out1;

  Logical_Operator_out6615_out1 <= Logical_Operator_out5591_out1 XOR Logical_Operator_out5623_out1;

  Logical_Operator_out6616_out1 <= Logical_Operator_out5592_out1 XOR Logical_Operator_out5624_out1;

  Logical_Operator_out6617_out1 <= Logical_Operator_out5593_out1 XOR Logical_Operator_out5625_out1;

  Logical_Operator_out6618_out1 <= Logical_Operator_out5594_out1 XOR Logical_Operator_out5626_out1;

  Logical_Operator_out6619_out1 <= Logical_Operator_out5595_out1 XOR Logical_Operator_out5627_out1;

  Logical_Operator_out6620_out1 <= Logical_Operator_out5596_out1 XOR Logical_Operator_out5628_out1;

  Logical_Operator_out6621_out1 <= Logical_Operator_out5597_out1 XOR Logical_Operator_out5629_out1;

  Logical_Operator_out6622_out1 <= Logical_Operator_out5598_out1 XOR Logical_Operator_out5630_out1;

  Logical_Operator_out6623_out1 <= Logical_Operator_out5599_out1 XOR Logical_Operator_out5631_out1;

  Logical_Operator_out6624_out1 <= Logical_Operator_out5600_out1 XOR Logical_Operator_out5632_out1;

  Logical_Operator_out6625_out1 <= Logical_Operator_out4561_out1 XOR Logical_Operator_out4593_out1;

  Logical_Operator_out6626_out1 <= Logical_Operator_out4562_out1 XOR Logical_Operator_out4594_out1;

  Logical_Operator_out6627_out1 <= Logical_Operator_out4563_out1 XOR Logical_Operator_out4595_out1;

  Logical_Operator_out6628_out1 <= Logical_Operator_out4564_out1 XOR Logical_Operator_out4596_out1;

  Logical_Operator_out6629_out1 <= Logical_Operator_out4565_out1 XOR Logical_Operator_out4597_out1;

  Logical_Operator_out6630_out1 <= Logical_Operator_out4566_out1 XOR Logical_Operator_out4598_out1;

  Logical_Operator_out6631_out1 <= Logical_Operator_out4567_out1 XOR Logical_Operator_out4599_out1;

  Logical_Operator_out6632_out1 <= Logical_Operator_out4568_out1 XOR Logical_Operator_out4600_out1;

  Logical_Operator_out6633_out1 <= Logical_Operator_out4569_out1 XOR Logical_Operator_out4601_out1;

  Logical_Operator_out6634_out1 <= Logical_Operator_out4570_out1 XOR Logical_Operator_out4602_out1;

  Logical_Operator_out6635_out1 <= Logical_Operator_out4571_out1 XOR Logical_Operator_out4603_out1;

  Logical_Operator_out6636_out1 <= Logical_Operator_out4572_out1 XOR Logical_Operator_out4604_out1;

  Logical_Operator_out6637_out1 <= Logical_Operator_out4573_out1 XOR Logical_Operator_out4605_out1;

  Logical_Operator_out6638_out1 <= Logical_Operator_out4574_out1 XOR Logical_Operator_out4606_out1;

  Logical_Operator_out6639_out1 <= Logical_Operator_out4575_out1 XOR Logical_Operator_out4607_out1;

  Logical_Operator_out6640_out1 <= Logical_Operator_out4576_out1 XOR Logical_Operator_out4608_out1;

  Logical_Operator_out6641_out1 <= Logical_Operator_out3545_out1 XOR Logical_Operator_out3577_out1;

  Logical_Operator_out6642_out1 <= Logical_Operator_out3546_out1 XOR Logical_Operator_out3578_out1;

  Logical_Operator_out6643_out1 <= Logical_Operator_out3547_out1 XOR Logical_Operator_out3579_out1;

  Logical_Operator_out6644_out1 <= Logical_Operator_out3548_out1 XOR Logical_Operator_out3580_out1;

  Logical_Operator_out6645_out1 <= Logical_Operator_out3549_out1 XOR Logical_Operator_out3581_out1;

  Logical_Operator_out6646_out1 <= Logical_Operator_out3550_out1 XOR Logical_Operator_out3582_out1;

  Logical_Operator_out6647_out1 <= Logical_Operator_out3551_out1 XOR Logical_Operator_out3583_out1;

  Logical_Operator_out6648_out1 <= Logical_Operator_out3552_out1 XOR Logical_Operator_out3584_out1;

  Logical_Operator_out6649_out1 <= Logical_Operator_out2525_out1 XOR Logical_Operator_out2557_out1;

  Logical_Operator_out6650_out1 <= Logical_Operator_out2526_out1 XOR Logical_Operator_out2558_out1;

  Logical_Operator_out6651_out1 <= Logical_Operator_out2527_out1 XOR Logical_Operator_out2559_out1;

  Logical_Operator_out6652_out1 <= Logical_Operator_out2528_out1 XOR Logical_Operator_out2560_out1;

  Logical_Operator_out6653_out1 <= Logical_Operator_out1503_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out6654_out1 <= Logical_Operator_out1504_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out6655_out1 <= Logical_Operator_out480_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out6656_out1 <= in960 XOR in1024;

  Logical_Operator_out6657_out1 <= Logical_Operator_out5633_out1 XOR Logical_Operator_out5665_out1;

  Logical_Operator_out6658_out1 <= Logical_Operator_out5634_out1 XOR Logical_Operator_out5666_out1;

  Logical_Operator_out6659_out1 <= Logical_Operator_out5635_out1 XOR Logical_Operator_out5667_out1;

  Logical_Operator_out6660_out1 <= Logical_Operator_out5636_out1 XOR Logical_Operator_out5668_out1;

  Logical_Operator_out6661_out1 <= Logical_Operator_out5637_out1 XOR Logical_Operator_out5669_out1;

  Logical_Operator_out6662_out1 <= Logical_Operator_out5638_out1 XOR Logical_Operator_out5670_out1;

  Logical_Operator_out6663_out1 <= Logical_Operator_out5639_out1 XOR Logical_Operator_out5671_out1;

  Logical_Operator_out6664_out1 <= Logical_Operator_out5640_out1 XOR Logical_Operator_out5672_out1;

  Logical_Operator_out6665_out1 <= Logical_Operator_out5641_out1 XOR Logical_Operator_out5673_out1;

  Logical_Operator_out6666_out1 <= Logical_Operator_out5642_out1 XOR Logical_Operator_out5674_out1;

  Logical_Operator_out6667_out1 <= Logical_Operator_out5643_out1 XOR Logical_Operator_out5675_out1;

  Logical_Operator_out6668_out1 <= Logical_Operator_out5644_out1 XOR Logical_Operator_out5676_out1;

  Logical_Operator_out6669_out1 <= Logical_Operator_out5645_out1 XOR Logical_Operator_out5677_out1;

  Logical_Operator_out6670_out1 <= Logical_Operator_out5646_out1 XOR Logical_Operator_out5678_out1;

  Logical_Operator_out6671_out1 <= Logical_Operator_out5647_out1 XOR Logical_Operator_out5679_out1;

  Logical_Operator_out6672_out1 <= Logical_Operator_out5648_out1 XOR Logical_Operator_out5680_out1;

  Logical_Operator_out6673_out1 <= Logical_Operator_out5649_out1 XOR Logical_Operator_out5681_out1;

  Logical_Operator_out6674_out1 <= Logical_Operator_out5650_out1 XOR Logical_Operator_out5682_out1;

  Logical_Operator_out6675_out1 <= Logical_Operator_out5651_out1 XOR Logical_Operator_out5683_out1;

  Logical_Operator_out6676_out1 <= Logical_Operator_out5652_out1 XOR Logical_Operator_out5684_out1;

  Logical_Operator_out6677_out1 <= Logical_Operator_out5653_out1 XOR Logical_Operator_out5685_out1;

  Logical_Operator_out6678_out1 <= Logical_Operator_out5654_out1 XOR Logical_Operator_out5686_out1;

  Logical_Operator_out6679_out1 <= Logical_Operator_out5655_out1 XOR Logical_Operator_out5687_out1;

  Logical_Operator_out6680_out1 <= Logical_Operator_out5656_out1 XOR Logical_Operator_out5688_out1;

  Logical_Operator_out6681_out1 <= Logical_Operator_out5657_out1 XOR Logical_Operator_out5689_out1;

  Logical_Operator_out6682_out1 <= Logical_Operator_out5658_out1 XOR Logical_Operator_out5690_out1;

  Logical_Operator_out6683_out1 <= Logical_Operator_out5659_out1 XOR Logical_Operator_out5691_out1;

  Logical_Operator_out6684_out1 <= Logical_Operator_out5660_out1 XOR Logical_Operator_out5692_out1;

  Logical_Operator_out6685_out1 <= Logical_Operator_out5661_out1 XOR Logical_Operator_out5693_out1;

  Logical_Operator_out6686_out1 <= Logical_Operator_out5662_out1 XOR Logical_Operator_out5694_out1;

  Logical_Operator_out6687_out1 <= Logical_Operator_out5663_out1 XOR Logical_Operator_out5695_out1;

  Logical_Operator_out6688_out1 <= Logical_Operator_out5664_out1 XOR Logical_Operator_out5696_out1;

  Logical_Operator_out6689_out1 <= Logical_Operator_out4625_out1 XOR Logical_Operator_out4657_out1;

  Logical_Operator_out6690_out1 <= Logical_Operator_out4626_out1 XOR Logical_Operator_out4658_out1;

  Logical_Operator_out6691_out1 <= Logical_Operator_out4627_out1 XOR Logical_Operator_out4659_out1;

  Logical_Operator_out6692_out1 <= Logical_Operator_out4628_out1 XOR Logical_Operator_out4660_out1;

  Logical_Operator_out6693_out1 <= Logical_Operator_out4629_out1 XOR Logical_Operator_out4661_out1;

  Logical_Operator_out6694_out1 <= Logical_Operator_out4630_out1 XOR Logical_Operator_out4662_out1;

  Logical_Operator_out6695_out1 <= Logical_Operator_out4631_out1 XOR Logical_Operator_out4663_out1;

  Logical_Operator_out6696_out1 <= Logical_Operator_out4632_out1 XOR Logical_Operator_out4664_out1;

  Logical_Operator_out6697_out1 <= Logical_Operator_out4633_out1 XOR Logical_Operator_out4665_out1;

  Logical_Operator_out6698_out1 <= Logical_Operator_out4634_out1 XOR Logical_Operator_out4666_out1;

  Logical_Operator_out6699_out1 <= Logical_Operator_out4635_out1 XOR Logical_Operator_out4667_out1;

  Logical_Operator_out6700_out1 <= Logical_Operator_out4636_out1 XOR Logical_Operator_out4668_out1;

  Logical_Operator_out6701_out1 <= Logical_Operator_out4637_out1 XOR Logical_Operator_out4669_out1;

  Logical_Operator_out6702_out1 <= Logical_Operator_out4638_out1 XOR Logical_Operator_out4670_out1;

  Logical_Operator_out6703_out1 <= Logical_Operator_out4639_out1 XOR Logical_Operator_out4671_out1;

  Logical_Operator_out6704_out1 <= Logical_Operator_out4640_out1 XOR Logical_Operator_out4672_out1;

  Logical_Operator_out6705_out1 <= Logical_Operator_out3609_out1 XOR Logical_Operator_out3641_out1;

  Logical_Operator_out6706_out1 <= Logical_Operator_out3610_out1 XOR Logical_Operator_out3642_out1;

  Logical_Operator_out6707_out1 <= Logical_Operator_out3611_out1 XOR Logical_Operator_out3643_out1;

  Logical_Operator_out6708_out1 <= Logical_Operator_out3612_out1 XOR Logical_Operator_out3644_out1;

  Logical_Operator_out6709_out1 <= Logical_Operator_out3613_out1 XOR Logical_Operator_out3645_out1;

  Logical_Operator_out6710_out1 <= Logical_Operator_out3614_out1 XOR Logical_Operator_out3646_out1;

  Logical_Operator_out6711_out1 <= Logical_Operator_out3615_out1 XOR Logical_Operator_out3647_out1;

  Logical_Operator_out6712_out1 <= Logical_Operator_out3616_out1 XOR Logical_Operator_out3648_out1;

  Logical_Operator_out6713_out1 <= Logical_Operator_out2589_out1 XOR Logical_Operator_out2621_out1;

  Logical_Operator_out6714_out1 <= Logical_Operator_out2590_out1 XOR Logical_Operator_out2622_out1;

  Logical_Operator_out6715_out1 <= Logical_Operator_out2591_out1 XOR Logical_Operator_out2623_out1;

  Logical_Operator_out6716_out1 <= Logical_Operator_out2592_out1 XOR Logical_Operator_out2624_out1;

  Logical_Operator_out6717_out1 <= Logical_Operator_out1567_out1 XOR Logical_Operator_out1599_out1;

  Logical_Operator_out6718_out1 <= Logical_Operator_out1568_out1 XOR Logical_Operator_out1600_out1;

  Logical_Operator_out6719_out1 <= Logical_Operator_out544_out1 XOR Logical_Operator_out576_out1;

  Logical_Operator_out6720_out1 <= in1088 XOR in1152;

  Logical_Operator_out6721_out1 <= Logical_Operator_out5697_out1 XOR Logical_Operator_out5729_out1;

  Logical_Operator_out6722_out1 <= Logical_Operator_out5698_out1 XOR Logical_Operator_out5730_out1;

  Logical_Operator_out6723_out1 <= Logical_Operator_out5699_out1 XOR Logical_Operator_out5731_out1;

  Logical_Operator_out6724_out1 <= Logical_Operator_out5700_out1 XOR Logical_Operator_out5732_out1;

  Logical_Operator_out6725_out1 <= Logical_Operator_out5701_out1 XOR Logical_Operator_out5733_out1;

  Logical_Operator_out6726_out1 <= Logical_Operator_out5702_out1 XOR Logical_Operator_out5734_out1;

  Logical_Operator_out6727_out1 <= Logical_Operator_out5703_out1 XOR Logical_Operator_out5735_out1;

  Logical_Operator_out6728_out1 <= Logical_Operator_out5704_out1 XOR Logical_Operator_out5736_out1;

  Logical_Operator_out6729_out1 <= Logical_Operator_out5705_out1 XOR Logical_Operator_out5737_out1;

  Logical_Operator_out6730_out1 <= Logical_Operator_out5706_out1 XOR Logical_Operator_out5738_out1;

  Logical_Operator_out6731_out1 <= Logical_Operator_out5707_out1 XOR Logical_Operator_out5739_out1;

  Logical_Operator_out6732_out1 <= Logical_Operator_out5708_out1 XOR Logical_Operator_out5740_out1;

  Logical_Operator_out6733_out1 <= Logical_Operator_out5709_out1 XOR Logical_Operator_out5741_out1;

  Logical_Operator_out6734_out1 <= Logical_Operator_out5710_out1 XOR Logical_Operator_out5742_out1;

  Logical_Operator_out6735_out1 <= Logical_Operator_out5711_out1 XOR Logical_Operator_out5743_out1;

  Logical_Operator_out6736_out1 <= Logical_Operator_out5712_out1 XOR Logical_Operator_out5744_out1;

  Logical_Operator_out6737_out1 <= Logical_Operator_out5713_out1 XOR Logical_Operator_out5745_out1;

  Logical_Operator_out6738_out1 <= Logical_Operator_out5714_out1 XOR Logical_Operator_out5746_out1;

  Logical_Operator_out6739_out1 <= Logical_Operator_out5715_out1 XOR Logical_Operator_out5747_out1;

  Logical_Operator_out6740_out1 <= Logical_Operator_out5716_out1 XOR Logical_Operator_out5748_out1;

  Logical_Operator_out6741_out1 <= Logical_Operator_out5717_out1 XOR Logical_Operator_out5749_out1;

  Logical_Operator_out6742_out1 <= Logical_Operator_out5718_out1 XOR Logical_Operator_out5750_out1;

  Logical_Operator_out6743_out1 <= Logical_Operator_out5719_out1 XOR Logical_Operator_out5751_out1;

  Logical_Operator_out6744_out1 <= Logical_Operator_out5720_out1 XOR Logical_Operator_out5752_out1;

  Logical_Operator_out6745_out1 <= Logical_Operator_out5721_out1 XOR Logical_Operator_out5753_out1;

  Logical_Operator_out6746_out1 <= Logical_Operator_out5722_out1 XOR Logical_Operator_out5754_out1;

  Logical_Operator_out6747_out1 <= Logical_Operator_out5723_out1 XOR Logical_Operator_out5755_out1;

  Logical_Operator_out6748_out1 <= Logical_Operator_out5724_out1 XOR Logical_Operator_out5756_out1;

  Logical_Operator_out6749_out1 <= Logical_Operator_out5725_out1 XOR Logical_Operator_out5757_out1;

  Logical_Operator_out6750_out1 <= Logical_Operator_out5726_out1 XOR Logical_Operator_out5758_out1;

  Logical_Operator_out6751_out1 <= Logical_Operator_out5727_out1 XOR Logical_Operator_out5759_out1;

  Logical_Operator_out6752_out1 <= Logical_Operator_out5728_out1 XOR Logical_Operator_out5760_out1;

  Logical_Operator_out6753_out1 <= Logical_Operator_out4689_out1 XOR Logical_Operator_out4721_out1;

  Logical_Operator_out6754_out1 <= Logical_Operator_out4690_out1 XOR Logical_Operator_out4722_out1;

  Logical_Operator_out6755_out1 <= Logical_Operator_out4691_out1 XOR Logical_Operator_out4723_out1;

  Logical_Operator_out6756_out1 <= Logical_Operator_out4692_out1 XOR Logical_Operator_out4724_out1;

  Logical_Operator_out6757_out1 <= Logical_Operator_out4693_out1 XOR Logical_Operator_out4725_out1;

  Logical_Operator_out6758_out1 <= Logical_Operator_out4694_out1 XOR Logical_Operator_out4726_out1;

  Logical_Operator_out6759_out1 <= Logical_Operator_out4695_out1 XOR Logical_Operator_out4727_out1;

  Logical_Operator_out6760_out1 <= Logical_Operator_out4696_out1 XOR Logical_Operator_out4728_out1;

  Logical_Operator_out6761_out1 <= Logical_Operator_out4697_out1 XOR Logical_Operator_out4729_out1;

  Logical_Operator_out6762_out1 <= Logical_Operator_out4698_out1 XOR Logical_Operator_out4730_out1;

  Logical_Operator_out6763_out1 <= Logical_Operator_out4699_out1 XOR Logical_Operator_out4731_out1;

  Logical_Operator_out6764_out1 <= Logical_Operator_out4700_out1 XOR Logical_Operator_out4732_out1;

  Logical_Operator_out6765_out1 <= Logical_Operator_out4701_out1 XOR Logical_Operator_out4733_out1;

  Logical_Operator_out6766_out1 <= Logical_Operator_out4702_out1 XOR Logical_Operator_out4734_out1;

  Logical_Operator_out6767_out1 <= Logical_Operator_out4703_out1 XOR Logical_Operator_out4735_out1;

  Logical_Operator_out6768_out1 <= Logical_Operator_out4704_out1 XOR Logical_Operator_out4736_out1;

  Logical_Operator_out6769_out1 <= Logical_Operator_out3673_out1 XOR Logical_Operator_out3705_out1;

  Logical_Operator_out6770_out1 <= Logical_Operator_out3674_out1 XOR Logical_Operator_out3706_out1;

  Logical_Operator_out6771_out1 <= Logical_Operator_out3675_out1 XOR Logical_Operator_out3707_out1;

  Logical_Operator_out6772_out1 <= Logical_Operator_out3676_out1 XOR Logical_Operator_out3708_out1;

  Logical_Operator_out6773_out1 <= Logical_Operator_out3677_out1 XOR Logical_Operator_out3709_out1;

  Logical_Operator_out6774_out1 <= Logical_Operator_out3678_out1 XOR Logical_Operator_out3710_out1;

  Logical_Operator_out6775_out1 <= Logical_Operator_out3679_out1 XOR Logical_Operator_out3711_out1;

  Logical_Operator_out6776_out1 <= Logical_Operator_out3680_out1 XOR Logical_Operator_out3712_out1;

  Logical_Operator_out6777_out1 <= Logical_Operator_out2653_out1 XOR Logical_Operator_out2685_out1;

  Logical_Operator_out6778_out1 <= Logical_Operator_out2654_out1 XOR Logical_Operator_out2686_out1;

  Logical_Operator_out6779_out1 <= Logical_Operator_out2655_out1 XOR Logical_Operator_out2687_out1;

  Logical_Operator_out6780_out1 <= Logical_Operator_out2656_out1 XOR Logical_Operator_out2688_out1;

  Logical_Operator_out6781_out1 <= Logical_Operator_out1631_out1 XOR Logical_Operator_out1663_out1;

  Logical_Operator_out6782_out1 <= Logical_Operator_out1632_out1 XOR Logical_Operator_out1664_out1;

  Logical_Operator_out6783_out1 <= Logical_Operator_out608_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out6784_out1 <= in1216 XOR in1280;

  Logical_Operator_out6785_out1 <= Logical_Operator_out5761_out1 XOR Logical_Operator_out5793_out1;

  Logical_Operator_out6786_out1 <= Logical_Operator_out5762_out1 XOR Logical_Operator_out5794_out1;

  Logical_Operator_out6787_out1 <= Logical_Operator_out5763_out1 XOR Logical_Operator_out5795_out1;

  Logical_Operator_out6788_out1 <= Logical_Operator_out5764_out1 XOR Logical_Operator_out5796_out1;

  Logical_Operator_out6789_out1 <= Logical_Operator_out5765_out1 XOR Logical_Operator_out5797_out1;

  Logical_Operator_out6790_out1 <= Logical_Operator_out5766_out1 XOR Logical_Operator_out5798_out1;

  Logical_Operator_out6791_out1 <= Logical_Operator_out5767_out1 XOR Logical_Operator_out5799_out1;

  Logical_Operator_out6792_out1 <= Logical_Operator_out5768_out1 XOR Logical_Operator_out5800_out1;

  Logical_Operator_out6793_out1 <= Logical_Operator_out5769_out1 XOR Logical_Operator_out5801_out1;

  Logical_Operator_out6794_out1 <= Logical_Operator_out5770_out1 XOR Logical_Operator_out5802_out1;

  Logical_Operator_out6795_out1 <= Logical_Operator_out5771_out1 XOR Logical_Operator_out5803_out1;

  Logical_Operator_out6796_out1 <= Logical_Operator_out5772_out1 XOR Logical_Operator_out5804_out1;

  Logical_Operator_out6797_out1 <= Logical_Operator_out5773_out1 XOR Logical_Operator_out5805_out1;

  Logical_Operator_out6798_out1 <= Logical_Operator_out5774_out1 XOR Logical_Operator_out5806_out1;

  Logical_Operator_out6799_out1 <= Logical_Operator_out5775_out1 XOR Logical_Operator_out5807_out1;

  Logical_Operator_out6800_out1 <= Logical_Operator_out5776_out1 XOR Logical_Operator_out5808_out1;

  Logical_Operator_out6801_out1 <= Logical_Operator_out5777_out1 XOR Logical_Operator_out5809_out1;

  Logical_Operator_out6802_out1 <= Logical_Operator_out5778_out1 XOR Logical_Operator_out5810_out1;

  Logical_Operator_out6803_out1 <= Logical_Operator_out5779_out1 XOR Logical_Operator_out5811_out1;

  Logical_Operator_out6804_out1 <= Logical_Operator_out5780_out1 XOR Logical_Operator_out5812_out1;

  Logical_Operator_out6805_out1 <= Logical_Operator_out5781_out1 XOR Logical_Operator_out5813_out1;

  Logical_Operator_out6806_out1 <= Logical_Operator_out5782_out1 XOR Logical_Operator_out5814_out1;

  Logical_Operator_out6807_out1 <= Logical_Operator_out5783_out1 XOR Logical_Operator_out5815_out1;

  Logical_Operator_out6808_out1 <= Logical_Operator_out5784_out1 XOR Logical_Operator_out5816_out1;

  Logical_Operator_out6809_out1 <= Logical_Operator_out5785_out1 XOR Logical_Operator_out5817_out1;

  Logical_Operator_out6810_out1 <= Logical_Operator_out5786_out1 XOR Logical_Operator_out5818_out1;

  Logical_Operator_out6811_out1 <= Logical_Operator_out5787_out1 XOR Logical_Operator_out5819_out1;

  Logical_Operator_out6812_out1 <= Logical_Operator_out5788_out1 XOR Logical_Operator_out5820_out1;

  Logical_Operator_out6813_out1 <= Logical_Operator_out5789_out1 XOR Logical_Operator_out5821_out1;

  Logical_Operator_out6814_out1 <= Logical_Operator_out5790_out1 XOR Logical_Operator_out5822_out1;

  Logical_Operator_out6815_out1 <= Logical_Operator_out5791_out1 XOR Logical_Operator_out5823_out1;

  Logical_Operator_out6816_out1 <= Logical_Operator_out5792_out1 XOR Logical_Operator_out5824_out1;

  Logical_Operator_out6817_out1 <= Logical_Operator_out4753_out1 XOR Logical_Operator_out4785_out1;

  Logical_Operator_out6818_out1 <= Logical_Operator_out4754_out1 XOR Logical_Operator_out4786_out1;

  Logical_Operator_out6819_out1 <= Logical_Operator_out4755_out1 XOR Logical_Operator_out4787_out1;

  Logical_Operator_out6820_out1 <= Logical_Operator_out4756_out1 XOR Logical_Operator_out4788_out1;

  Logical_Operator_out6821_out1 <= Logical_Operator_out4757_out1 XOR Logical_Operator_out4789_out1;

  Logical_Operator_out6822_out1 <= Logical_Operator_out4758_out1 XOR Logical_Operator_out4790_out1;

  Logical_Operator_out6823_out1 <= Logical_Operator_out4759_out1 XOR Logical_Operator_out4791_out1;

  Logical_Operator_out6824_out1 <= Logical_Operator_out4760_out1 XOR Logical_Operator_out4792_out1;

  Logical_Operator_out6825_out1 <= Logical_Operator_out4761_out1 XOR Logical_Operator_out4793_out1;

  Logical_Operator_out6826_out1 <= Logical_Operator_out4762_out1 XOR Logical_Operator_out4794_out1;

  Logical_Operator_out6827_out1 <= Logical_Operator_out4763_out1 XOR Logical_Operator_out4795_out1;

  Logical_Operator_out6828_out1 <= Logical_Operator_out4764_out1 XOR Logical_Operator_out4796_out1;

  Logical_Operator_out6829_out1 <= Logical_Operator_out4765_out1 XOR Logical_Operator_out4797_out1;

  Logical_Operator_out6830_out1 <= Logical_Operator_out4766_out1 XOR Logical_Operator_out4798_out1;

  Logical_Operator_out6831_out1 <= Logical_Operator_out4767_out1 XOR Logical_Operator_out4799_out1;

  Logical_Operator_out6832_out1 <= Logical_Operator_out4768_out1 XOR Logical_Operator_out4800_out1;

  Logical_Operator_out6833_out1 <= Logical_Operator_out3737_out1 XOR Logical_Operator_out3769_out1;

  Logical_Operator_out6834_out1 <= Logical_Operator_out3738_out1 XOR Logical_Operator_out3770_out1;

  Logical_Operator_out6835_out1 <= Logical_Operator_out3739_out1 XOR Logical_Operator_out3771_out1;

  Logical_Operator_out6836_out1 <= Logical_Operator_out3740_out1 XOR Logical_Operator_out3772_out1;

  Logical_Operator_out6837_out1 <= Logical_Operator_out3741_out1 XOR Logical_Operator_out3773_out1;

  Logical_Operator_out6838_out1 <= Logical_Operator_out3742_out1 XOR Logical_Operator_out3774_out1;

  Logical_Operator_out6839_out1 <= Logical_Operator_out3743_out1 XOR Logical_Operator_out3775_out1;

  Logical_Operator_out6840_out1 <= Logical_Operator_out3744_out1 XOR Logical_Operator_out3776_out1;

  Logical_Operator_out6841_out1 <= Logical_Operator_out2717_out1 XOR Logical_Operator_out2749_out1;

  Logical_Operator_out6842_out1 <= Logical_Operator_out2718_out1 XOR Logical_Operator_out2750_out1;

  Logical_Operator_out6843_out1 <= Logical_Operator_out2719_out1 XOR Logical_Operator_out2751_out1;

  Logical_Operator_out6844_out1 <= Logical_Operator_out2720_out1 XOR Logical_Operator_out2752_out1;

  Logical_Operator_out6845_out1 <= Logical_Operator_out1695_out1 XOR Logical_Operator_out1727_out1;

  Logical_Operator_out6846_out1 <= Logical_Operator_out1696_out1 XOR Logical_Operator_out1728_out1;

  Logical_Operator_out6847_out1 <= Logical_Operator_out672_out1 XOR Logical_Operator_out704_out1;

  Logical_Operator_out6848_out1 <= in1344 XOR in1408;

  Logical_Operator_out6849_out1 <= Logical_Operator_out5825_out1 XOR Logical_Operator_out5857_out1;

  Logical_Operator_out6850_out1 <= Logical_Operator_out5826_out1 XOR Logical_Operator_out5858_out1;

  Logical_Operator_out6851_out1 <= Logical_Operator_out5827_out1 XOR Logical_Operator_out5859_out1;

  Logical_Operator_out6852_out1 <= Logical_Operator_out5828_out1 XOR Logical_Operator_out5860_out1;

  Logical_Operator_out6853_out1 <= Logical_Operator_out5829_out1 XOR Logical_Operator_out5861_out1;

  Logical_Operator_out6854_out1 <= Logical_Operator_out5830_out1 XOR Logical_Operator_out5862_out1;

  Logical_Operator_out6855_out1 <= Logical_Operator_out5831_out1 XOR Logical_Operator_out5863_out1;

  Logical_Operator_out6856_out1 <= Logical_Operator_out5832_out1 XOR Logical_Operator_out5864_out1;

  Logical_Operator_out6857_out1 <= Logical_Operator_out5833_out1 XOR Logical_Operator_out5865_out1;

  Logical_Operator_out6858_out1 <= Logical_Operator_out5834_out1 XOR Logical_Operator_out5866_out1;

  Logical_Operator_out6859_out1 <= Logical_Operator_out5835_out1 XOR Logical_Operator_out5867_out1;

  Logical_Operator_out6860_out1 <= Logical_Operator_out5836_out1 XOR Logical_Operator_out5868_out1;

  Logical_Operator_out6861_out1 <= Logical_Operator_out5837_out1 XOR Logical_Operator_out5869_out1;

  Logical_Operator_out6862_out1 <= Logical_Operator_out5838_out1 XOR Logical_Operator_out5870_out1;

  Logical_Operator_out6863_out1 <= Logical_Operator_out5839_out1 XOR Logical_Operator_out5871_out1;

  Logical_Operator_out6864_out1 <= Logical_Operator_out5840_out1 XOR Logical_Operator_out5872_out1;

  Logical_Operator_out6865_out1 <= Logical_Operator_out5841_out1 XOR Logical_Operator_out5873_out1;

  Logical_Operator_out6866_out1 <= Logical_Operator_out5842_out1 XOR Logical_Operator_out5874_out1;

  Logical_Operator_out6867_out1 <= Logical_Operator_out5843_out1 XOR Logical_Operator_out5875_out1;

  Logical_Operator_out6868_out1 <= Logical_Operator_out5844_out1 XOR Logical_Operator_out5876_out1;

  Logical_Operator_out6869_out1 <= Logical_Operator_out5845_out1 XOR Logical_Operator_out5877_out1;

  Logical_Operator_out6870_out1 <= Logical_Operator_out5846_out1 XOR Logical_Operator_out5878_out1;

  Logical_Operator_out6871_out1 <= Logical_Operator_out5847_out1 XOR Logical_Operator_out5879_out1;

  Logical_Operator_out6872_out1 <= Logical_Operator_out5848_out1 XOR Logical_Operator_out5880_out1;

  Logical_Operator_out6873_out1 <= Logical_Operator_out5849_out1 XOR Logical_Operator_out5881_out1;

  Logical_Operator_out6874_out1 <= Logical_Operator_out5850_out1 XOR Logical_Operator_out5882_out1;

  Logical_Operator_out6875_out1 <= Logical_Operator_out5851_out1 XOR Logical_Operator_out5883_out1;

  Logical_Operator_out6876_out1 <= Logical_Operator_out5852_out1 XOR Logical_Operator_out5884_out1;

  Logical_Operator_out6877_out1 <= Logical_Operator_out5853_out1 XOR Logical_Operator_out5885_out1;

  Logical_Operator_out6878_out1 <= Logical_Operator_out5854_out1 XOR Logical_Operator_out5886_out1;

  Logical_Operator_out6879_out1 <= Logical_Operator_out5855_out1 XOR Logical_Operator_out5887_out1;

  Logical_Operator_out6880_out1 <= Logical_Operator_out5856_out1 XOR Logical_Operator_out5888_out1;

  Logical_Operator_out6881_out1 <= Logical_Operator_out4817_out1 XOR Logical_Operator_out4849_out1;

  Logical_Operator_out6882_out1 <= Logical_Operator_out4818_out1 XOR Logical_Operator_out4850_out1;

  Logical_Operator_out6883_out1 <= Logical_Operator_out4819_out1 XOR Logical_Operator_out4851_out1;

  Logical_Operator_out6884_out1 <= Logical_Operator_out4820_out1 XOR Logical_Operator_out4852_out1;

  Logical_Operator_out6885_out1 <= Logical_Operator_out4821_out1 XOR Logical_Operator_out4853_out1;

  Logical_Operator_out6886_out1 <= Logical_Operator_out4822_out1 XOR Logical_Operator_out4854_out1;

  Logical_Operator_out6887_out1 <= Logical_Operator_out4823_out1 XOR Logical_Operator_out4855_out1;

  Logical_Operator_out6888_out1 <= Logical_Operator_out4824_out1 XOR Logical_Operator_out4856_out1;

  Logical_Operator_out6889_out1 <= Logical_Operator_out4825_out1 XOR Logical_Operator_out4857_out1;

  Logical_Operator_out6890_out1 <= Logical_Operator_out4826_out1 XOR Logical_Operator_out4858_out1;

  Logical_Operator_out6891_out1 <= Logical_Operator_out4827_out1 XOR Logical_Operator_out4859_out1;

  Logical_Operator_out6892_out1 <= Logical_Operator_out4828_out1 XOR Logical_Operator_out4860_out1;

  Logical_Operator_out6893_out1 <= Logical_Operator_out4829_out1 XOR Logical_Operator_out4861_out1;

  Logical_Operator_out6894_out1 <= Logical_Operator_out4830_out1 XOR Logical_Operator_out4862_out1;

  Logical_Operator_out6895_out1 <= Logical_Operator_out4831_out1 XOR Logical_Operator_out4863_out1;

  Logical_Operator_out6896_out1 <= Logical_Operator_out4832_out1 XOR Logical_Operator_out4864_out1;

  Logical_Operator_out6897_out1 <= Logical_Operator_out3801_out1 XOR Logical_Operator_out3833_out1;

  Logical_Operator_out6898_out1 <= Logical_Operator_out3802_out1 XOR Logical_Operator_out3834_out1;

  Logical_Operator_out6899_out1 <= Logical_Operator_out3803_out1 XOR Logical_Operator_out3835_out1;

  Logical_Operator_out6900_out1 <= Logical_Operator_out3804_out1 XOR Logical_Operator_out3836_out1;

  Logical_Operator_out6901_out1 <= Logical_Operator_out3805_out1 XOR Logical_Operator_out3837_out1;

  Logical_Operator_out6902_out1 <= Logical_Operator_out3806_out1 XOR Logical_Operator_out3838_out1;

  Logical_Operator_out6903_out1 <= Logical_Operator_out3807_out1 XOR Logical_Operator_out3839_out1;

  Logical_Operator_out6904_out1 <= Logical_Operator_out3808_out1 XOR Logical_Operator_out3840_out1;

  Logical_Operator_out6905_out1 <= Logical_Operator_out2781_out1 XOR Logical_Operator_out2813_out1;

  Logical_Operator_out6906_out1 <= Logical_Operator_out2782_out1 XOR Logical_Operator_out2814_out1;

  Logical_Operator_out6907_out1 <= Logical_Operator_out2783_out1 XOR Logical_Operator_out2815_out1;

  Logical_Operator_out6908_out1 <= Logical_Operator_out2784_out1 XOR Logical_Operator_out2816_out1;

  Logical_Operator_out6909_out1 <= Logical_Operator_out1759_out1 XOR Logical_Operator_out1791_out1;

  Logical_Operator_out6910_out1 <= Logical_Operator_out1760_out1 XOR Logical_Operator_out1792_out1;

  Logical_Operator_out6911_out1 <= Logical_Operator_out736_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out6912_out1 <= in1472 XOR in1536;

  Logical_Operator_out6913_out1 <= Logical_Operator_out5889_out1 XOR Logical_Operator_out5921_out1;

  Logical_Operator_out6914_out1 <= Logical_Operator_out5890_out1 XOR Logical_Operator_out5922_out1;

  Logical_Operator_out6915_out1 <= Logical_Operator_out5891_out1 XOR Logical_Operator_out5923_out1;

  Logical_Operator_out6916_out1 <= Logical_Operator_out5892_out1 XOR Logical_Operator_out5924_out1;

  Logical_Operator_out6917_out1 <= Logical_Operator_out5893_out1 XOR Logical_Operator_out5925_out1;

  Logical_Operator_out6918_out1 <= Logical_Operator_out5894_out1 XOR Logical_Operator_out5926_out1;

  Logical_Operator_out6919_out1 <= Logical_Operator_out5895_out1 XOR Logical_Operator_out5927_out1;

  Logical_Operator_out6920_out1 <= Logical_Operator_out5896_out1 XOR Logical_Operator_out5928_out1;

  Logical_Operator_out6921_out1 <= Logical_Operator_out5897_out1 XOR Logical_Operator_out5929_out1;

  Logical_Operator_out6922_out1 <= Logical_Operator_out5898_out1 XOR Logical_Operator_out5930_out1;

  Logical_Operator_out6923_out1 <= Logical_Operator_out5899_out1 XOR Logical_Operator_out5931_out1;

  Logical_Operator_out6924_out1 <= Logical_Operator_out5900_out1 XOR Logical_Operator_out5932_out1;

  Logical_Operator_out6925_out1 <= Logical_Operator_out5901_out1 XOR Logical_Operator_out5933_out1;

  Logical_Operator_out6926_out1 <= Logical_Operator_out5902_out1 XOR Logical_Operator_out5934_out1;

  Logical_Operator_out6927_out1 <= Logical_Operator_out5903_out1 XOR Logical_Operator_out5935_out1;

  Logical_Operator_out6928_out1 <= Logical_Operator_out5904_out1 XOR Logical_Operator_out5936_out1;

  Logical_Operator_out6929_out1 <= Logical_Operator_out5905_out1 XOR Logical_Operator_out5937_out1;

  Logical_Operator_out6930_out1 <= Logical_Operator_out5906_out1 XOR Logical_Operator_out5938_out1;

  Logical_Operator_out6931_out1 <= Logical_Operator_out5907_out1 XOR Logical_Operator_out5939_out1;

  Logical_Operator_out6932_out1 <= Logical_Operator_out5908_out1 XOR Logical_Operator_out5940_out1;

  Logical_Operator_out6933_out1 <= Logical_Operator_out5909_out1 XOR Logical_Operator_out5941_out1;

  Logical_Operator_out6934_out1 <= Logical_Operator_out5910_out1 XOR Logical_Operator_out5942_out1;

  Logical_Operator_out6935_out1 <= Logical_Operator_out5911_out1 XOR Logical_Operator_out5943_out1;

  Logical_Operator_out6936_out1 <= Logical_Operator_out5912_out1 XOR Logical_Operator_out5944_out1;

  Logical_Operator_out6937_out1 <= Logical_Operator_out5913_out1 XOR Logical_Operator_out5945_out1;

  Logical_Operator_out6938_out1 <= Logical_Operator_out5914_out1 XOR Logical_Operator_out5946_out1;

  Logical_Operator_out6939_out1 <= Logical_Operator_out5915_out1 XOR Logical_Operator_out5947_out1;

  Logical_Operator_out6940_out1 <= Logical_Operator_out5916_out1 XOR Logical_Operator_out5948_out1;

  Logical_Operator_out6941_out1 <= Logical_Operator_out5917_out1 XOR Logical_Operator_out5949_out1;

  Logical_Operator_out6942_out1 <= Logical_Operator_out5918_out1 XOR Logical_Operator_out5950_out1;

  Logical_Operator_out6943_out1 <= Logical_Operator_out5919_out1 XOR Logical_Operator_out5951_out1;

  Logical_Operator_out6944_out1 <= Logical_Operator_out5920_out1 XOR Logical_Operator_out5952_out1;

  Logical_Operator_out6945_out1 <= Logical_Operator_out4881_out1 XOR Logical_Operator_out4913_out1;

  Logical_Operator_out6946_out1 <= Logical_Operator_out4882_out1 XOR Logical_Operator_out4914_out1;

  Logical_Operator_out6947_out1 <= Logical_Operator_out4883_out1 XOR Logical_Operator_out4915_out1;

  Logical_Operator_out6948_out1 <= Logical_Operator_out4884_out1 XOR Logical_Operator_out4916_out1;

  Logical_Operator_out6949_out1 <= Logical_Operator_out4885_out1 XOR Logical_Operator_out4917_out1;

  Logical_Operator_out6950_out1 <= Logical_Operator_out4886_out1 XOR Logical_Operator_out4918_out1;

  Logical_Operator_out6951_out1 <= Logical_Operator_out4887_out1 XOR Logical_Operator_out4919_out1;

  Logical_Operator_out6952_out1 <= Logical_Operator_out4888_out1 XOR Logical_Operator_out4920_out1;

  Logical_Operator_out6953_out1 <= Logical_Operator_out4889_out1 XOR Logical_Operator_out4921_out1;

  Logical_Operator_out6954_out1 <= Logical_Operator_out4890_out1 XOR Logical_Operator_out4922_out1;

  Logical_Operator_out6955_out1 <= Logical_Operator_out4891_out1 XOR Logical_Operator_out4923_out1;

  Logical_Operator_out6956_out1 <= Logical_Operator_out4892_out1 XOR Logical_Operator_out4924_out1;

  Logical_Operator_out6957_out1 <= Logical_Operator_out4893_out1 XOR Logical_Operator_out4925_out1;

  Logical_Operator_out6958_out1 <= Logical_Operator_out4894_out1 XOR Logical_Operator_out4926_out1;

  Logical_Operator_out6959_out1 <= Logical_Operator_out4895_out1 XOR Logical_Operator_out4927_out1;

  Logical_Operator_out6960_out1 <= Logical_Operator_out4896_out1 XOR Logical_Operator_out4928_out1;

  Logical_Operator_out6961_out1 <= Logical_Operator_out3865_out1 XOR Logical_Operator_out3897_out1;

  Logical_Operator_out6962_out1 <= Logical_Operator_out3866_out1 XOR Logical_Operator_out3898_out1;

  Logical_Operator_out6963_out1 <= Logical_Operator_out3867_out1 XOR Logical_Operator_out3899_out1;

  Logical_Operator_out6964_out1 <= Logical_Operator_out3868_out1 XOR Logical_Operator_out3900_out1;

  Logical_Operator_out6965_out1 <= Logical_Operator_out3869_out1 XOR Logical_Operator_out3901_out1;

  Logical_Operator_out6966_out1 <= Logical_Operator_out3870_out1 XOR Logical_Operator_out3902_out1;

  Logical_Operator_out6967_out1 <= Logical_Operator_out3871_out1 XOR Logical_Operator_out3903_out1;

  Logical_Operator_out6968_out1 <= Logical_Operator_out3872_out1 XOR Logical_Operator_out3904_out1;

  Logical_Operator_out6969_out1 <= Logical_Operator_out2845_out1 XOR Logical_Operator_out2877_out1;

  Logical_Operator_out6970_out1 <= Logical_Operator_out2846_out1 XOR Logical_Operator_out2878_out1;

  Logical_Operator_out6971_out1 <= Logical_Operator_out2847_out1 XOR Logical_Operator_out2879_out1;

  Logical_Operator_out6972_out1 <= Logical_Operator_out2848_out1 XOR Logical_Operator_out2880_out1;

  Logical_Operator_out6973_out1 <= Logical_Operator_out1823_out1 XOR Logical_Operator_out1855_out1;

  Logical_Operator_out6974_out1 <= Logical_Operator_out1824_out1 XOR Logical_Operator_out1856_out1;

  Logical_Operator_out6975_out1 <= Logical_Operator_out800_out1 XOR Logical_Operator_out832_out1;

  Logical_Operator_out6976_out1 <= in1600 XOR in1664;

  Logical_Operator_out6977_out1 <= Logical_Operator_out5953_out1 XOR Logical_Operator_out5985_out1;

  Logical_Operator_out6978_out1 <= Logical_Operator_out5954_out1 XOR Logical_Operator_out5986_out1;

  Logical_Operator_out6979_out1 <= Logical_Operator_out5955_out1 XOR Logical_Operator_out5987_out1;

  Logical_Operator_out6980_out1 <= Logical_Operator_out5956_out1 XOR Logical_Operator_out5988_out1;

  Logical_Operator_out6981_out1 <= Logical_Operator_out5957_out1 XOR Logical_Operator_out5989_out1;

  Logical_Operator_out6982_out1 <= Logical_Operator_out5958_out1 XOR Logical_Operator_out5990_out1;

  Logical_Operator_out6983_out1 <= Logical_Operator_out5959_out1 XOR Logical_Operator_out5991_out1;

  Logical_Operator_out6984_out1 <= Logical_Operator_out5960_out1 XOR Logical_Operator_out5992_out1;

  Logical_Operator_out6985_out1 <= Logical_Operator_out5961_out1 XOR Logical_Operator_out5993_out1;

  Logical_Operator_out6986_out1 <= Logical_Operator_out5962_out1 XOR Logical_Operator_out5994_out1;

  Logical_Operator_out6987_out1 <= Logical_Operator_out5963_out1 XOR Logical_Operator_out5995_out1;

  Logical_Operator_out6988_out1 <= Logical_Operator_out5964_out1 XOR Logical_Operator_out5996_out1;

  Logical_Operator_out6989_out1 <= Logical_Operator_out5965_out1 XOR Logical_Operator_out5997_out1;

  Logical_Operator_out6990_out1 <= Logical_Operator_out5966_out1 XOR Logical_Operator_out5998_out1;

  Logical_Operator_out6991_out1 <= Logical_Operator_out5967_out1 XOR Logical_Operator_out5999_out1;

  Logical_Operator_out6992_out1 <= Logical_Operator_out5968_out1 XOR Logical_Operator_out6000_out1;

  Logical_Operator_out6993_out1 <= Logical_Operator_out5969_out1 XOR Logical_Operator_out6001_out1;

  Logical_Operator_out6994_out1 <= Logical_Operator_out5970_out1 XOR Logical_Operator_out6002_out1;

  Logical_Operator_out6995_out1 <= Logical_Operator_out5971_out1 XOR Logical_Operator_out6003_out1;

  Logical_Operator_out6996_out1 <= Logical_Operator_out5972_out1 XOR Logical_Operator_out6004_out1;

  Logical_Operator_out6997_out1 <= Logical_Operator_out5973_out1 XOR Logical_Operator_out6005_out1;

  Logical_Operator_out6998_out1 <= Logical_Operator_out5974_out1 XOR Logical_Operator_out6006_out1;

  Logical_Operator_out6999_out1 <= Logical_Operator_out5975_out1 XOR Logical_Operator_out6007_out1;

  Logical_Operator_out7000_out1 <= Logical_Operator_out5976_out1 XOR Logical_Operator_out6008_out1;

  Logical_Operator_out7001_out1 <= Logical_Operator_out5977_out1 XOR Logical_Operator_out6009_out1;

  Logical_Operator_out7002_out1 <= Logical_Operator_out5978_out1 XOR Logical_Operator_out6010_out1;

  Logical_Operator_out7003_out1 <= Logical_Operator_out5979_out1 XOR Logical_Operator_out6011_out1;

  Logical_Operator_out7004_out1 <= Logical_Operator_out5980_out1 XOR Logical_Operator_out6012_out1;

  Logical_Operator_out7005_out1 <= Logical_Operator_out5981_out1 XOR Logical_Operator_out6013_out1;

  Logical_Operator_out7006_out1 <= Logical_Operator_out5982_out1 XOR Logical_Operator_out6014_out1;

  Logical_Operator_out7007_out1 <= Logical_Operator_out5983_out1 XOR Logical_Operator_out6015_out1;

  Logical_Operator_out7008_out1 <= Logical_Operator_out5984_out1 XOR Logical_Operator_out6016_out1;

  Logical_Operator_out7009_out1 <= Logical_Operator_out4945_out1 XOR Logical_Operator_out4977_out1;

  Logical_Operator_out7010_out1 <= Logical_Operator_out4946_out1 XOR Logical_Operator_out4978_out1;

  Logical_Operator_out7011_out1 <= Logical_Operator_out4947_out1 XOR Logical_Operator_out4979_out1;

  Logical_Operator_out7012_out1 <= Logical_Operator_out4948_out1 XOR Logical_Operator_out4980_out1;

  Logical_Operator_out7013_out1 <= Logical_Operator_out4949_out1 XOR Logical_Operator_out4981_out1;

  Logical_Operator_out7014_out1 <= Logical_Operator_out4950_out1 XOR Logical_Operator_out4982_out1;

  Logical_Operator_out7015_out1 <= Logical_Operator_out4951_out1 XOR Logical_Operator_out4983_out1;

  Logical_Operator_out7016_out1 <= Logical_Operator_out4952_out1 XOR Logical_Operator_out4984_out1;

  Logical_Operator_out7017_out1 <= Logical_Operator_out4953_out1 XOR Logical_Operator_out4985_out1;

  Logical_Operator_out7018_out1 <= Logical_Operator_out4954_out1 XOR Logical_Operator_out4986_out1;

  Logical_Operator_out7019_out1 <= Logical_Operator_out4955_out1 XOR Logical_Operator_out4987_out1;

  Logical_Operator_out7020_out1 <= Logical_Operator_out4956_out1 XOR Logical_Operator_out4988_out1;

  Logical_Operator_out7021_out1 <= Logical_Operator_out4957_out1 XOR Logical_Operator_out4989_out1;

  Logical_Operator_out7022_out1 <= Logical_Operator_out4958_out1 XOR Logical_Operator_out4990_out1;

  Logical_Operator_out7023_out1 <= Logical_Operator_out4959_out1 XOR Logical_Operator_out4991_out1;

  Logical_Operator_out7024_out1 <= Logical_Operator_out4960_out1 XOR Logical_Operator_out4992_out1;

  Logical_Operator_out7025_out1 <= Logical_Operator_out3929_out1 XOR Logical_Operator_out3961_out1;

  Logical_Operator_out7026_out1 <= Logical_Operator_out3930_out1 XOR Logical_Operator_out3962_out1;

  Logical_Operator_out7027_out1 <= Logical_Operator_out3931_out1 XOR Logical_Operator_out3963_out1;

  Logical_Operator_out7028_out1 <= Logical_Operator_out3932_out1 XOR Logical_Operator_out3964_out1;

  Logical_Operator_out7029_out1 <= Logical_Operator_out3933_out1 XOR Logical_Operator_out3965_out1;

  Logical_Operator_out7030_out1 <= Logical_Operator_out3934_out1 XOR Logical_Operator_out3966_out1;

  Logical_Operator_out7031_out1 <= Logical_Operator_out3935_out1 XOR Logical_Operator_out3967_out1;

  Logical_Operator_out7032_out1 <= Logical_Operator_out3936_out1 XOR Logical_Operator_out3968_out1;

  Logical_Operator_out7033_out1 <= Logical_Operator_out2909_out1 XOR Logical_Operator_out2941_out1;

  Logical_Operator_out7034_out1 <= Logical_Operator_out2910_out1 XOR Logical_Operator_out2942_out1;

  Logical_Operator_out7035_out1 <= Logical_Operator_out2911_out1 XOR Logical_Operator_out2943_out1;

  Logical_Operator_out7036_out1 <= Logical_Operator_out2912_out1 XOR Logical_Operator_out2944_out1;

  Logical_Operator_out7037_out1 <= Logical_Operator_out1887_out1 XOR Logical_Operator_out1919_out1;

  Logical_Operator_out7038_out1 <= Logical_Operator_out1888_out1 XOR Logical_Operator_out1920_out1;

  Logical_Operator_out7039_out1 <= Logical_Operator_out864_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out7040_out1 <= in1728 XOR in1792;

  Logical_Operator_out7041_out1 <= Logical_Operator_out6017_out1 XOR Logical_Operator_out6049_out1;

  Logical_Operator_out7042_out1 <= Logical_Operator_out6018_out1 XOR Logical_Operator_out6050_out1;

  Logical_Operator_out7043_out1 <= Logical_Operator_out6019_out1 XOR Logical_Operator_out6051_out1;

  Logical_Operator_out7044_out1 <= Logical_Operator_out6020_out1 XOR Logical_Operator_out6052_out1;

  Logical_Operator_out7045_out1 <= Logical_Operator_out6021_out1 XOR Logical_Operator_out6053_out1;

  Logical_Operator_out7046_out1 <= Logical_Operator_out6022_out1 XOR Logical_Operator_out6054_out1;

  Logical_Operator_out7047_out1 <= Logical_Operator_out6023_out1 XOR Logical_Operator_out6055_out1;

  Logical_Operator_out7048_out1 <= Logical_Operator_out6024_out1 XOR Logical_Operator_out6056_out1;

  Logical_Operator_out7049_out1 <= Logical_Operator_out6025_out1 XOR Logical_Operator_out6057_out1;

  Logical_Operator_out7050_out1 <= Logical_Operator_out6026_out1 XOR Logical_Operator_out6058_out1;

  Logical_Operator_out7051_out1 <= Logical_Operator_out6027_out1 XOR Logical_Operator_out6059_out1;

  Logical_Operator_out7052_out1 <= Logical_Operator_out6028_out1 XOR Logical_Operator_out6060_out1;

  Logical_Operator_out7053_out1 <= Logical_Operator_out6029_out1 XOR Logical_Operator_out6061_out1;

  Logical_Operator_out7054_out1 <= Logical_Operator_out6030_out1 XOR Logical_Operator_out6062_out1;

  Logical_Operator_out7055_out1 <= Logical_Operator_out6031_out1 XOR Logical_Operator_out6063_out1;

  Logical_Operator_out7056_out1 <= Logical_Operator_out6032_out1 XOR Logical_Operator_out6064_out1;

  Logical_Operator_out7057_out1 <= Logical_Operator_out6033_out1 XOR Logical_Operator_out6065_out1;

  Logical_Operator_out7058_out1 <= Logical_Operator_out6034_out1 XOR Logical_Operator_out6066_out1;

  Logical_Operator_out7059_out1 <= Logical_Operator_out6035_out1 XOR Logical_Operator_out6067_out1;

  Logical_Operator_out7060_out1 <= Logical_Operator_out6036_out1 XOR Logical_Operator_out6068_out1;

  Logical_Operator_out7061_out1 <= Logical_Operator_out6037_out1 XOR Logical_Operator_out6069_out1;

  Logical_Operator_out7062_out1 <= Logical_Operator_out6038_out1 XOR Logical_Operator_out6070_out1;

  Logical_Operator_out7063_out1 <= Logical_Operator_out6039_out1 XOR Logical_Operator_out6071_out1;

  Logical_Operator_out7064_out1 <= Logical_Operator_out6040_out1 XOR Logical_Operator_out6072_out1;

  Logical_Operator_out7065_out1 <= Logical_Operator_out6041_out1 XOR Logical_Operator_out6073_out1;

  Logical_Operator_out7066_out1 <= Logical_Operator_out6042_out1 XOR Logical_Operator_out6074_out1;

  Logical_Operator_out7067_out1 <= Logical_Operator_out6043_out1 XOR Logical_Operator_out6075_out1;

  Logical_Operator_out7068_out1 <= Logical_Operator_out6044_out1 XOR Logical_Operator_out6076_out1;

  Logical_Operator_out7069_out1 <= Logical_Operator_out6045_out1 XOR Logical_Operator_out6077_out1;

  Logical_Operator_out7070_out1 <= Logical_Operator_out6046_out1 XOR Logical_Operator_out6078_out1;

  Logical_Operator_out7071_out1 <= Logical_Operator_out6047_out1 XOR Logical_Operator_out6079_out1;

  Logical_Operator_out7072_out1 <= Logical_Operator_out6048_out1 XOR Logical_Operator_out6080_out1;

  Logical_Operator_out7073_out1 <= Logical_Operator_out5009_out1 XOR Logical_Operator_out5041_out1;

  Logical_Operator_out7074_out1 <= Logical_Operator_out5010_out1 XOR Logical_Operator_out5042_out1;

  Logical_Operator_out7075_out1 <= Logical_Operator_out5011_out1 XOR Logical_Operator_out5043_out1;

  Logical_Operator_out7076_out1 <= Logical_Operator_out5012_out1 XOR Logical_Operator_out5044_out1;

  Logical_Operator_out7077_out1 <= Logical_Operator_out5013_out1 XOR Logical_Operator_out5045_out1;

  Logical_Operator_out7078_out1 <= Logical_Operator_out5014_out1 XOR Logical_Operator_out5046_out1;

  Logical_Operator_out7079_out1 <= Logical_Operator_out5015_out1 XOR Logical_Operator_out5047_out1;

  Logical_Operator_out7080_out1 <= Logical_Operator_out5016_out1 XOR Logical_Operator_out5048_out1;

  Logical_Operator_out7081_out1 <= Logical_Operator_out5017_out1 XOR Logical_Operator_out5049_out1;

  Logical_Operator_out7082_out1 <= Logical_Operator_out5018_out1 XOR Logical_Operator_out5050_out1;

  Logical_Operator_out7083_out1 <= Logical_Operator_out5019_out1 XOR Logical_Operator_out5051_out1;

  Logical_Operator_out7084_out1 <= Logical_Operator_out5020_out1 XOR Logical_Operator_out5052_out1;

  Logical_Operator_out7085_out1 <= Logical_Operator_out5021_out1 XOR Logical_Operator_out5053_out1;

  Logical_Operator_out7086_out1 <= Logical_Operator_out5022_out1 XOR Logical_Operator_out5054_out1;

  Logical_Operator_out7087_out1 <= Logical_Operator_out5023_out1 XOR Logical_Operator_out5055_out1;

  Logical_Operator_out7088_out1 <= Logical_Operator_out5024_out1 XOR Logical_Operator_out5056_out1;

  Logical_Operator_out7089_out1 <= Logical_Operator_out3993_out1 XOR Logical_Operator_out4025_out1;

  Logical_Operator_out7090_out1 <= Logical_Operator_out3994_out1 XOR Logical_Operator_out4026_out1;

  Logical_Operator_out7091_out1 <= Logical_Operator_out3995_out1 XOR Logical_Operator_out4027_out1;

  Logical_Operator_out7092_out1 <= Logical_Operator_out3996_out1 XOR Logical_Operator_out4028_out1;

  Logical_Operator_out7093_out1 <= Logical_Operator_out3997_out1 XOR Logical_Operator_out4029_out1;

  Logical_Operator_out7094_out1 <= Logical_Operator_out3998_out1 XOR Logical_Operator_out4030_out1;

  Logical_Operator_out7095_out1 <= Logical_Operator_out3999_out1 XOR Logical_Operator_out4031_out1;

  Logical_Operator_out7096_out1 <= Logical_Operator_out4000_out1 XOR Logical_Operator_out4032_out1;

  Logical_Operator_out7097_out1 <= Logical_Operator_out2973_out1 XOR Logical_Operator_out3005_out1;

  Logical_Operator_out7098_out1 <= Logical_Operator_out2974_out1 XOR Logical_Operator_out3006_out1;

  Logical_Operator_out7099_out1 <= Logical_Operator_out2975_out1 XOR Logical_Operator_out3007_out1;

  Logical_Operator_out7100_out1 <= Logical_Operator_out2976_out1 XOR Logical_Operator_out3008_out1;

  Logical_Operator_out7101_out1 <= Logical_Operator_out1951_out1 XOR Logical_Operator_out1983_out1;

  Logical_Operator_out7102_out1 <= Logical_Operator_out1952_out1 XOR Logical_Operator_out1984_out1;

  Logical_Operator_out7103_out1 <= Logical_Operator_out928_out1 XOR Logical_Operator_out960_out1;

  Logical_Operator_out7104_out1 <= in1856 XOR in1920;

  Logical_Operator_out7105_out1 <= Logical_Operator_out6081_out1 XOR Logical_Operator_out6113_out1;

  Logical_Operator_out7106_out1 <= Logical_Operator_out6082_out1 XOR Logical_Operator_out6114_out1;

  Logical_Operator_out7107_out1 <= Logical_Operator_out6083_out1 XOR Logical_Operator_out6115_out1;

  Logical_Operator_out7108_out1 <= Logical_Operator_out6084_out1 XOR Logical_Operator_out6116_out1;

  Logical_Operator_out7109_out1 <= Logical_Operator_out6085_out1 XOR Logical_Operator_out6117_out1;

  Logical_Operator_out7110_out1 <= Logical_Operator_out6086_out1 XOR Logical_Operator_out6118_out1;

  Logical_Operator_out7111_out1 <= Logical_Operator_out6087_out1 XOR Logical_Operator_out6119_out1;

  Logical_Operator_out7112_out1 <= Logical_Operator_out6088_out1 XOR Logical_Operator_out6120_out1;

  Logical_Operator_out7113_out1 <= Logical_Operator_out6089_out1 XOR Logical_Operator_out6121_out1;

  Logical_Operator_out7114_out1 <= Logical_Operator_out6090_out1 XOR Logical_Operator_out6122_out1;

  Logical_Operator_out7115_out1 <= Logical_Operator_out6091_out1 XOR Logical_Operator_out6123_out1;

  Logical_Operator_out7116_out1 <= Logical_Operator_out6092_out1 XOR Logical_Operator_out6124_out1;

  Logical_Operator_out7117_out1 <= Logical_Operator_out6093_out1 XOR Logical_Operator_out6125_out1;

  Logical_Operator_out7118_out1 <= Logical_Operator_out6094_out1 XOR Logical_Operator_out6126_out1;

  Logical_Operator_out7119_out1 <= Logical_Operator_out6095_out1 XOR Logical_Operator_out6127_out1;

  Logical_Operator_out7120_out1 <= Logical_Operator_out6096_out1 XOR Logical_Operator_out6128_out1;

  Logical_Operator_out7121_out1 <= Logical_Operator_out6097_out1 XOR Logical_Operator_out6129_out1;

  Logical_Operator_out7122_out1 <= Logical_Operator_out6098_out1 XOR Logical_Operator_out6130_out1;

  Logical_Operator_out7123_out1 <= Logical_Operator_out6099_out1 XOR Logical_Operator_out6131_out1;

  Logical_Operator_out7124_out1 <= Logical_Operator_out6100_out1 XOR Logical_Operator_out6132_out1;

  Logical_Operator_out7125_out1 <= Logical_Operator_out6101_out1 XOR Logical_Operator_out6133_out1;

  Logical_Operator_out7126_out1 <= Logical_Operator_out6102_out1 XOR Logical_Operator_out6134_out1;

  Logical_Operator_out7127_out1 <= Logical_Operator_out6103_out1 XOR Logical_Operator_out6135_out1;

  Logical_Operator_out7128_out1 <= Logical_Operator_out6104_out1 XOR Logical_Operator_out6136_out1;

  Logical_Operator_out7129_out1 <= Logical_Operator_out6105_out1 XOR Logical_Operator_out6137_out1;

  Logical_Operator_out7130_out1 <= Logical_Operator_out6106_out1 XOR Logical_Operator_out6138_out1;

  Logical_Operator_out7131_out1 <= Logical_Operator_out6107_out1 XOR Logical_Operator_out6139_out1;

  Logical_Operator_out7132_out1 <= Logical_Operator_out6108_out1 XOR Logical_Operator_out6140_out1;

  Logical_Operator_out7133_out1 <= Logical_Operator_out6109_out1 XOR Logical_Operator_out6141_out1;

  Logical_Operator_out7134_out1 <= Logical_Operator_out6110_out1 XOR Logical_Operator_out6142_out1;

  Logical_Operator_out7135_out1 <= Logical_Operator_out6111_out1 XOR Logical_Operator_out6143_out1;

  Logical_Operator_out7136_out1 <= Logical_Operator_out6112_out1 XOR Logical_Operator_out6144_out1;

  Logical_Operator_out7137_out1 <= Logical_Operator_out5073_out1 XOR Logical_Operator_out5105_out1;

  Logical_Operator_out7138_out1 <= Logical_Operator_out5074_out1 XOR Logical_Operator_out5106_out1;

  Logical_Operator_out7139_out1 <= Logical_Operator_out5075_out1 XOR Logical_Operator_out5107_out1;

  Logical_Operator_out7140_out1 <= Logical_Operator_out5076_out1 XOR Logical_Operator_out5108_out1;

  Logical_Operator_out7141_out1 <= Logical_Operator_out5077_out1 XOR Logical_Operator_out5109_out1;

  Logical_Operator_out7142_out1 <= Logical_Operator_out5078_out1 XOR Logical_Operator_out5110_out1;

  Logical_Operator_out7143_out1 <= Logical_Operator_out5079_out1 XOR Logical_Operator_out5111_out1;

  Logical_Operator_out7144_out1 <= Logical_Operator_out5080_out1 XOR Logical_Operator_out5112_out1;

  Logical_Operator_out7145_out1 <= Logical_Operator_out5081_out1 XOR Logical_Operator_out5113_out1;

  Logical_Operator_out7146_out1 <= Logical_Operator_out5082_out1 XOR Logical_Operator_out5114_out1;

  Logical_Operator_out7147_out1 <= Logical_Operator_out5083_out1 XOR Logical_Operator_out5115_out1;

  Logical_Operator_out7148_out1 <= Logical_Operator_out5084_out1 XOR Logical_Operator_out5116_out1;

  Logical_Operator_out7149_out1 <= Logical_Operator_out5085_out1 XOR Logical_Operator_out5117_out1;

  Logical_Operator_out7150_out1 <= Logical_Operator_out5086_out1 XOR Logical_Operator_out5118_out1;

  Logical_Operator_out7151_out1 <= Logical_Operator_out5087_out1 XOR Logical_Operator_out5119_out1;

  Logical_Operator_out7152_out1 <= Logical_Operator_out5088_out1 XOR Logical_Operator_out5120_out1;

  Logical_Operator_out7153_out1 <= Logical_Operator_out4057_out1 XOR Logical_Operator_out4089_out1;

  Logical_Operator_out7154_out1 <= Logical_Operator_out4058_out1 XOR Logical_Operator_out4090_out1;

  Logical_Operator_out7155_out1 <= Logical_Operator_out4059_out1 XOR Logical_Operator_out4091_out1;

  Logical_Operator_out7156_out1 <= Logical_Operator_out4060_out1 XOR Logical_Operator_out4092_out1;

  Logical_Operator_out7157_out1 <= Logical_Operator_out4061_out1 XOR Logical_Operator_out4093_out1;

  Logical_Operator_out7158_out1 <= Logical_Operator_out4062_out1 XOR Logical_Operator_out4094_out1;

  Logical_Operator_out7159_out1 <= Logical_Operator_out4063_out1 XOR Logical_Operator_out4095_out1;

  Logical_Operator_out7160_out1 <= Logical_Operator_out4064_out1 XOR Logical_Operator_out4096_out1;

  Logical_Operator_out7161_out1 <= Logical_Operator_out3037_out1 XOR Logical_Operator_out3069_out1;

  Logical_Operator_out7162_out1 <= Logical_Operator_out3038_out1 XOR Logical_Operator_out3070_out1;

  Logical_Operator_out7163_out1 <= Logical_Operator_out3039_out1 XOR Logical_Operator_out3071_out1;

  Logical_Operator_out7164_out1 <= Logical_Operator_out3040_out1 XOR Logical_Operator_out3072_out1;

  Logical_Operator_out7165_out1 <= Logical_Operator_out2015_out1 XOR Logical_Operator_out2047_out1;

  Logical_Operator_out7166_out1 <= Logical_Operator_out2016_out1 XOR Logical_Operator_out2048_out1;

  Logical_Operator_out7167_out1 <= Logical_Operator_out992_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out7168_out1 <= in1984 XOR in2048;

  Logical_Operator_out7169_out1 <= Logical_Operator_out6145_out1 XOR Logical_Operator_out6209_out1;

  Logical_Operator_out7170_out1 <= Logical_Operator_out6146_out1 XOR Logical_Operator_out6210_out1;

  Logical_Operator_out7171_out1 <= Logical_Operator_out6147_out1 XOR Logical_Operator_out6211_out1;

  Logical_Operator_out7172_out1 <= Logical_Operator_out6148_out1 XOR Logical_Operator_out6212_out1;

  Logical_Operator_out7173_out1 <= Logical_Operator_out6149_out1 XOR Logical_Operator_out6213_out1;

  Logical_Operator_out7174_out1 <= Logical_Operator_out6150_out1 XOR Logical_Operator_out6214_out1;

  Logical_Operator_out7175_out1 <= Logical_Operator_out6151_out1 XOR Logical_Operator_out6215_out1;

  Logical_Operator_out7176_out1 <= Logical_Operator_out6152_out1 XOR Logical_Operator_out6216_out1;

  Logical_Operator_out7177_out1 <= Logical_Operator_out6153_out1 XOR Logical_Operator_out6217_out1;

  Logical_Operator_out7178_out1 <= Logical_Operator_out6154_out1 XOR Logical_Operator_out6218_out1;

  Logical_Operator_out7179_out1 <= Logical_Operator_out6155_out1 XOR Logical_Operator_out6219_out1;

  Logical_Operator_out7180_out1 <= Logical_Operator_out6156_out1 XOR Logical_Operator_out6220_out1;

  Logical_Operator_out7181_out1 <= Logical_Operator_out6157_out1 XOR Logical_Operator_out6221_out1;

  Logical_Operator_out7182_out1 <= Logical_Operator_out6158_out1 XOR Logical_Operator_out6222_out1;

  Logical_Operator_out7183_out1 <= Logical_Operator_out6159_out1 XOR Logical_Operator_out6223_out1;

  Logical_Operator_out7184_out1 <= Logical_Operator_out6160_out1 XOR Logical_Operator_out6224_out1;

  Logical_Operator_out7185_out1 <= Logical_Operator_out6161_out1 XOR Logical_Operator_out6225_out1;

  Logical_Operator_out7186_out1 <= Logical_Operator_out6162_out1 XOR Logical_Operator_out6226_out1;

  Logical_Operator_out7187_out1 <= Logical_Operator_out6163_out1 XOR Logical_Operator_out6227_out1;

  Logical_Operator_out7188_out1 <= Logical_Operator_out6164_out1 XOR Logical_Operator_out6228_out1;

  Logical_Operator_out7189_out1 <= Logical_Operator_out6165_out1 XOR Logical_Operator_out6229_out1;

  Logical_Operator_out7190_out1 <= Logical_Operator_out6166_out1 XOR Logical_Operator_out6230_out1;

  Logical_Operator_out7191_out1 <= Logical_Operator_out6167_out1 XOR Logical_Operator_out6231_out1;

  Logical_Operator_out7192_out1 <= Logical_Operator_out6168_out1 XOR Logical_Operator_out6232_out1;

  Logical_Operator_out7193_out1 <= Logical_Operator_out6169_out1 XOR Logical_Operator_out6233_out1;

  Logical_Operator_out7194_out1 <= Logical_Operator_out6170_out1 XOR Logical_Operator_out6234_out1;

  Logical_Operator_out7195_out1 <= Logical_Operator_out6171_out1 XOR Logical_Operator_out6235_out1;

  Logical_Operator_out7196_out1 <= Logical_Operator_out6172_out1 XOR Logical_Operator_out6236_out1;

  Logical_Operator_out7197_out1 <= Logical_Operator_out6173_out1 XOR Logical_Operator_out6237_out1;

  Logical_Operator_out7198_out1 <= Logical_Operator_out6174_out1 XOR Logical_Operator_out6238_out1;

  Logical_Operator_out7199_out1 <= Logical_Operator_out6175_out1 XOR Logical_Operator_out6239_out1;

  Logical_Operator_out7200_out1 <= Logical_Operator_out6176_out1 XOR Logical_Operator_out6240_out1;

  Logical_Operator_out7201_out1 <= Logical_Operator_out6177_out1 XOR Logical_Operator_out6241_out1;

  Logical_Operator_out7202_out1 <= Logical_Operator_out6178_out1 XOR Logical_Operator_out6242_out1;

  Logical_Operator_out7203_out1 <= Logical_Operator_out6179_out1 XOR Logical_Operator_out6243_out1;

  Logical_Operator_out7204_out1 <= Logical_Operator_out6180_out1 XOR Logical_Operator_out6244_out1;

  Logical_Operator_out7205_out1 <= Logical_Operator_out6181_out1 XOR Logical_Operator_out6245_out1;

  Logical_Operator_out7206_out1 <= Logical_Operator_out6182_out1 XOR Logical_Operator_out6246_out1;

  Logical_Operator_out7207_out1 <= Logical_Operator_out6183_out1 XOR Logical_Operator_out6247_out1;

  Logical_Operator_out7208_out1 <= Logical_Operator_out6184_out1 XOR Logical_Operator_out6248_out1;

  Logical_Operator_out7209_out1 <= Logical_Operator_out6185_out1 XOR Logical_Operator_out6249_out1;

  Logical_Operator_out7210_out1 <= Logical_Operator_out6186_out1 XOR Logical_Operator_out6250_out1;

  Logical_Operator_out7211_out1 <= Logical_Operator_out6187_out1 XOR Logical_Operator_out6251_out1;

  Logical_Operator_out7212_out1 <= Logical_Operator_out6188_out1 XOR Logical_Operator_out6252_out1;

  Logical_Operator_out7213_out1 <= Logical_Operator_out6189_out1 XOR Logical_Operator_out6253_out1;

  Logical_Operator_out7214_out1 <= Logical_Operator_out6190_out1 XOR Logical_Operator_out6254_out1;

  Logical_Operator_out7215_out1 <= Logical_Operator_out6191_out1 XOR Logical_Operator_out6255_out1;

  Logical_Operator_out7216_out1 <= Logical_Operator_out6192_out1 XOR Logical_Operator_out6256_out1;

  Logical_Operator_out7217_out1 <= Logical_Operator_out6193_out1 XOR Logical_Operator_out6257_out1;

  Logical_Operator_out7218_out1 <= Logical_Operator_out6194_out1 XOR Logical_Operator_out6258_out1;

  Logical_Operator_out7219_out1 <= Logical_Operator_out6195_out1 XOR Logical_Operator_out6259_out1;

  Logical_Operator_out7220_out1 <= Logical_Operator_out6196_out1 XOR Logical_Operator_out6260_out1;

  Logical_Operator_out7221_out1 <= Logical_Operator_out6197_out1 XOR Logical_Operator_out6261_out1;

  Logical_Operator_out7222_out1 <= Logical_Operator_out6198_out1 XOR Logical_Operator_out6262_out1;

  Logical_Operator_out7223_out1 <= Logical_Operator_out6199_out1 XOR Logical_Operator_out6263_out1;

  Logical_Operator_out7224_out1 <= Logical_Operator_out6200_out1 XOR Logical_Operator_out6264_out1;

  Logical_Operator_out7225_out1 <= Logical_Operator_out6201_out1 XOR Logical_Operator_out6265_out1;

  Logical_Operator_out7226_out1 <= Logical_Operator_out6202_out1 XOR Logical_Operator_out6266_out1;

  Logical_Operator_out7227_out1 <= Logical_Operator_out6203_out1 XOR Logical_Operator_out6267_out1;

  Logical_Operator_out7228_out1 <= Logical_Operator_out6204_out1 XOR Logical_Operator_out6268_out1;

  Logical_Operator_out7229_out1 <= Logical_Operator_out6205_out1 XOR Logical_Operator_out6269_out1;

  Logical_Operator_out7230_out1 <= Logical_Operator_out6206_out1 XOR Logical_Operator_out6270_out1;

  Logical_Operator_out7231_out1 <= Logical_Operator_out6207_out1 XOR Logical_Operator_out6271_out1;

  Logical_Operator_out7232_out1 <= Logical_Operator_out6208_out1 XOR Logical_Operator_out6272_out1;

  Logical_Operator_out7233_out1 <= Logical_Operator_out5153_out1 XOR Logical_Operator_out5217_out1;

  Logical_Operator_out7234_out1 <= Logical_Operator_out5154_out1 XOR Logical_Operator_out5218_out1;

  Logical_Operator_out7235_out1 <= Logical_Operator_out5155_out1 XOR Logical_Operator_out5219_out1;

  Logical_Operator_out7236_out1 <= Logical_Operator_out5156_out1 XOR Logical_Operator_out5220_out1;

  Logical_Operator_out7237_out1 <= Logical_Operator_out5157_out1 XOR Logical_Operator_out5221_out1;

  Logical_Operator_out7238_out1 <= Logical_Operator_out5158_out1 XOR Logical_Operator_out5222_out1;

  Logical_Operator_out7239_out1 <= Logical_Operator_out5159_out1 XOR Logical_Operator_out5223_out1;

  Logical_Operator_out7240_out1 <= Logical_Operator_out5160_out1 XOR Logical_Operator_out5224_out1;

  Logical_Operator_out7241_out1 <= Logical_Operator_out5161_out1 XOR Logical_Operator_out5225_out1;

  Logical_Operator_out7242_out1 <= Logical_Operator_out5162_out1 XOR Logical_Operator_out5226_out1;

  Logical_Operator_out7243_out1 <= Logical_Operator_out5163_out1 XOR Logical_Operator_out5227_out1;

  Logical_Operator_out7244_out1 <= Logical_Operator_out5164_out1 XOR Logical_Operator_out5228_out1;

  Logical_Operator_out7245_out1 <= Logical_Operator_out5165_out1 XOR Logical_Operator_out5229_out1;

  Logical_Operator_out7246_out1 <= Logical_Operator_out5166_out1 XOR Logical_Operator_out5230_out1;

  Logical_Operator_out7247_out1 <= Logical_Operator_out5167_out1 XOR Logical_Operator_out5231_out1;

  Logical_Operator_out7248_out1 <= Logical_Operator_out5168_out1 XOR Logical_Operator_out5232_out1;

  Logical_Operator_out7249_out1 <= Logical_Operator_out5169_out1 XOR Logical_Operator_out5233_out1;

  Logical_Operator_out7250_out1 <= Logical_Operator_out5170_out1 XOR Logical_Operator_out5234_out1;

  Logical_Operator_out7251_out1 <= Logical_Operator_out5171_out1 XOR Logical_Operator_out5235_out1;

  Logical_Operator_out7252_out1 <= Logical_Operator_out5172_out1 XOR Logical_Operator_out5236_out1;

  Logical_Operator_out7253_out1 <= Logical_Operator_out5173_out1 XOR Logical_Operator_out5237_out1;

  Logical_Operator_out7254_out1 <= Logical_Operator_out5174_out1 XOR Logical_Operator_out5238_out1;

  Logical_Operator_out7255_out1 <= Logical_Operator_out5175_out1 XOR Logical_Operator_out5239_out1;

  Logical_Operator_out7256_out1 <= Logical_Operator_out5176_out1 XOR Logical_Operator_out5240_out1;

  Logical_Operator_out7257_out1 <= Logical_Operator_out5177_out1 XOR Logical_Operator_out5241_out1;

  Logical_Operator_out7258_out1 <= Logical_Operator_out5178_out1 XOR Logical_Operator_out5242_out1;

  Logical_Operator_out7259_out1 <= Logical_Operator_out5179_out1 XOR Logical_Operator_out5243_out1;

  Logical_Operator_out7260_out1 <= Logical_Operator_out5180_out1 XOR Logical_Operator_out5244_out1;

  Logical_Operator_out7261_out1 <= Logical_Operator_out5181_out1 XOR Logical_Operator_out5245_out1;

  Logical_Operator_out7262_out1 <= Logical_Operator_out5182_out1 XOR Logical_Operator_out5246_out1;

  Logical_Operator_out7263_out1 <= Logical_Operator_out5183_out1 XOR Logical_Operator_out5247_out1;

  Logical_Operator_out7264_out1 <= Logical_Operator_out5184_out1 XOR Logical_Operator_out5248_out1;

  Logical_Operator_out7265_out1 <= Logical_Operator_out4145_out1 XOR Logical_Operator_out4209_out1;

  Logical_Operator_out7266_out1 <= Logical_Operator_out4146_out1 XOR Logical_Operator_out4210_out1;

  Logical_Operator_out7267_out1 <= Logical_Operator_out4147_out1 XOR Logical_Operator_out4211_out1;

  Logical_Operator_out7268_out1 <= Logical_Operator_out4148_out1 XOR Logical_Operator_out4212_out1;

  Logical_Operator_out7269_out1 <= Logical_Operator_out4149_out1 XOR Logical_Operator_out4213_out1;

  Logical_Operator_out7270_out1 <= Logical_Operator_out4150_out1 XOR Logical_Operator_out4214_out1;

  Logical_Operator_out7271_out1 <= Logical_Operator_out4151_out1 XOR Logical_Operator_out4215_out1;

  Logical_Operator_out7272_out1 <= Logical_Operator_out4152_out1 XOR Logical_Operator_out4216_out1;

  Logical_Operator_out7273_out1 <= Logical_Operator_out4153_out1 XOR Logical_Operator_out4217_out1;

  Logical_Operator_out7274_out1 <= Logical_Operator_out4154_out1 XOR Logical_Operator_out4218_out1;

  Logical_Operator_out7275_out1 <= Logical_Operator_out4155_out1 XOR Logical_Operator_out4219_out1;

  Logical_Operator_out7276_out1 <= Logical_Operator_out4156_out1 XOR Logical_Operator_out4220_out1;

  Logical_Operator_out7277_out1 <= Logical_Operator_out4157_out1 XOR Logical_Operator_out4221_out1;

  Logical_Operator_out7278_out1 <= Logical_Operator_out4158_out1 XOR Logical_Operator_out4222_out1;

  Logical_Operator_out7279_out1 <= Logical_Operator_out4159_out1 XOR Logical_Operator_out4223_out1;

  Logical_Operator_out7280_out1 <= Logical_Operator_out4160_out1 XOR Logical_Operator_out4224_out1;

  Logical_Operator_out7281_out1 <= Logical_Operator_out3129_out1 XOR Logical_Operator_out3193_out1;

  Logical_Operator_out7282_out1 <= Logical_Operator_out3130_out1 XOR Logical_Operator_out3194_out1;

  Logical_Operator_out7283_out1 <= Logical_Operator_out3131_out1 XOR Logical_Operator_out3195_out1;

  Logical_Operator_out7284_out1 <= Logical_Operator_out3132_out1 XOR Logical_Operator_out3196_out1;

  Logical_Operator_out7285_out1 <= Logical_Operator_out3133_out1 XOR Logical_Operator_out3197_out1;

  Logical_Operator_out7286_out1 <= Logical_Operator_out3134_out1 XOR Logical_Operator_out3198_out1;

  Logical_Operator_out7287_out1 <= Logical_Operator_out3135_out1 XOR Logical_Operator_out3199_out1;

  Logical_Operator_out7288_out1 <= Logical_Operator_out3136_out1 XOR Logical_Operator_out3200_out1;

  Logical_Operator_out7289_out1 <= Logical_Operator_out2109_out1 XOR Logical_Operator_out2173_out1;

  Logical_Operator_out7290_out1 <= Logical_Operator_out2110_out1 XOR Logical_Operator_out2174_out1;

  Logical_Operator_out7291_out1 <= Logical_Operator_out2111_out1 XOR Logical_Operator_out2175_out1;

  Logical_Operator_out7292_out1 <= Logical_Operator_out2112_out1 XOR Logical_Operator_out2176_out1;

  Logical_Operator_out7293_out1 <= Logical_Operator_out1087_out1 XOR Logical_Operator_out1151_out1;

  Logical_Operator_out7294_out1 <= Logical_Operator_out1088_out1 XOR Logical_Operator_out1152_out1;

  Logical_Operator_out7295_out1 <= Logical_Operator_out64_out1 XOR Logical_Operator_out128_out1;

  Logical_Operator_out7296_out1 <= in128 XOR in256;

  Logical_Operator_out7297_out1 <= Logical_Operator_out6273_out1 XOR Logical_Operator_out6337_out1;

  Logical_Operator_out7298_out1 <= Logical_Operator_out6274_out1 XOR Logical_Operator_out6338_out1;

  Logical_Operator_out7299_out1 <= Logical_Operator_out6275_out1 XOR Logical_Operator_out6339_out1;

  Logical_Operator_out7300_out1 <= Logical_Operator_out6276_out1 XOR Logical_Operator_out6340_out1;

  Logical_Operator_out7301_out1 <= Logical_Operator_out6277_out1 XOR Logical_Operator_out6341_out1;

  Logical_Operator_out7302_out1 <= Logical_Operator_out6278_out1 XOR Logical_Operator_out6342_out1;

  Logical_Operator_out7303_out1 <= Logical_Operator_out6279_out1 XOR Logical_Operator_out6343_out1;

  Logical_Operator_out7304_out1 <= Logical_Operator_out6280_out1 XOR Logical_Operator_out6344_out1;

  Logical_Operator_out7305_out1 <= Logical_Operator_out6281_out1 XOR Logical_Operator_out6345_out1;

  Logical_Operator_out7306_out1 <= Logical_Operator_out6282_out1 XOR Logical_Operator_out6346_out1;

  Logical_Operator_out7307_out1 <= Logical_Operator_out6283_out1 XOR Logical_Operator_out6347_out1;

  Logical_Operator_out7308_out1 <= Logical_Operator_out6284_out1 XOR Logical_Operator_out6348_out1;

  Logical_Operator_out7309_out1 <= Logical_Operator_out6285_out1 XOR Logical_Operator_out6349_out1;

  Logical_Operator_out7310_out1 <= Logical_Operator_out6286_out1 XOR Logical_Operator_out6350_out1;

  Logical_Operator_out7311_out1 <= Logical_Operator_out6287_out1 XOR Logical_Operator_out6351_out1;

  Logical_Operator_out7312_out1 <= Logical_Operator_out6288_out1 XOR Logical_Operator_out6352_out1;

  Logical_Operator_out7313_out1 <= Logical_Operator_out6289_out1 XOR Logical_Operator_out6353_out1;

  Logical_Operator_out7314_out1 <= Logical_Operator_out6290_out1 XOR Logical_Operator_out6354_out1;

  Logical_Operator_out7315_out1 <= Logical_Operator_out6291_out1 XOR Logical_Operator_out6355_out1;

  Logical_Operator_out7316_out1 <= Logical_Operator_out6292_out1 XOR Logical_Operator_out6356_out1;

  Logical_Operator_out7317_out1 <= Logical_Operator_out6293_out1 XOR Logical_Operator_out6357_out1;

  Logical_Operator_out7318_out1 <= Logical_Operator_out6294_out1 XOR Logical_Operator_out6358_out1;

  Logical_Operator_out7319_out1 <= Logical_Operator_out6295_out1 XOR Logical_Operator_out6359_out1;

  Logical_Operator_out7320_out1 <= Logical_Operator_out6296_out1 XOR Logical_Operator_out6360_out1;

  Logical_Operator_out7321_out1 <= Logical_Operator_out6297_out1 XOR Logical_Operator_out6361_out1;

  Logical_Operator_out7322_out1 <= Logical_Operator_out6298_out1 XOR Logical_Operator_out6362_out1;

  Logical_Operator_out7323_out1 <= Logical_Operator_out6299_out1 XOR Logical_Operator_out6363_out1;

  Logical_Operator_out7324_out1 <= Logical_Operator_out6300_out1 XOR Logical_Operator_out6364_out1;

  Logical_Operator_out7325_out1 <= Logical_Operator_out6301_out1 XOR Logical_Operator_out6365_out1;

  Logical_Operator_out7326_out1 <= Logical_Operator_out6302_out1 XOR Logical_Operator_out6366_out1;

  Logical_Operator_out7327_out1 <= Logical_Operator_out6303_out1 XOR Logical_Operator_out6367_out1;

  Logical_Operator_out7328_out1 <= Logical_Operator_out6304_out1 XOR Logical_Operator_out6368_out1;

  Logical_Operator_out7329_out1 <= Logical_Operator_out6305_out1 XOR Logical_Operator_out6369_out1;

  Logical_Operator_out7330_out1 <= Logical_Operator_out6306_out1 XOR Logical_Operator_out6370_out1;

  Logical_Operator_out7331_out1 <= Logical_Operator_out6307_out1 XOR Logical_Operator_out6371_out1;

  Logical_Operator_out7332_out1 <= Logical_Operator_out6308_out1 XOR Logical_Operator_out6372_out1;

  Logical_Operator_out7333_out1 <= Logical_Operator_out6309_out1 XOR Logical_Operator_out6373_out1;

  Logical_Operator_out7334_out1 <= Logical_Operator_out6310_out1 XOR Logical_Operator_out6374_out1;

  Logical_Operator_out7335_out1 <= Logical_Operator_out6311_out1 XOR Logical_Operator_out6375_out1;

  Logical_Operator_out7336_out1 <= Logical_Operator_out6312_out1 XOR Logical_Operator_out6376_out1;

  Logical_Operator_out7337_out1 <= Logical_Operator_out6313_out1 XOR Logical_Operator_out6377_out1;

  Logical_Operator_out7338_out1 <= Logical_Operator_out6314_out1 XOR Logical_Operator_out6378_out1;

  Logical_Operator_out7339_out1 <= Logical_Operator_out6315_out1 XOR Logical_Operator_out6379_out1;

  Logical_Operator_out7340_out1 <= Logical_Operator_out6316_out1 XOR Logical_Operator_out6380_out1;

  Logical_Operator_out7341_out1 <= Logical_Operator_out6317_out1 XOR Logical_Operator_out6381_out1;

  Logical_Operator_out7342_out1 <= Logical_Operator_out6318_out1 XOR Logical_Operator_out6382_out1;

  Logical_Operator_out7343_out1 <= Logical_Operator_out6319_out1 XOR Logical_Operator_out6383_out1;

  Logical_Operator_out7344_out1 <= Logical_Operator_out6320_out1 XOR Logical_Operator_out6384_out1;

  Logical_Operator_out7345_out1 <= Logical_Operator_out6321_out1 XOR Logical_Operator_out6385_out1;

  Logical_Operator_out7346_out1 <= Logical_Operator_out6322_out1 XOR Logical_Operator_out6386_out1;

  Logical_Operator_out7347_out1 <= Logical_Operator_out6323_out1 XOR Logical_Operator_out6387_out1;

  Logical_Operator_out7348_out1 <= Logical_Operator_out6324_out1 XOR Logical_Operator_out6388_out1;

  Logical_Operator_out7349_out1 <= Logical_Operator_out6325_out1 XOR Logical_Operator_out6389_out1;

  Logical_Operator_out7350_out1 <= Logical_Operator_out6326_out1 XOR Logical_Operator_out6390_out1;

  Logical_Operator_out7351_out1 <= Logical_Operator_out6327_out1 XOR Logical_Operator_out6391_out1;

  Logical_Operator_out7352_out1 <= Logical_Operator_out6328_out1 XOR Logical_Operator_out6392_out1;

  Logical_Operator_out7353_out1 <= Logical_Operator_out6329_out1 XOR Logical_Operator_out6393_out1;

  Logical_Operator_out7354_out1 <= Logical_Operator_out6330_out1 XOR Logical_Operator_out6394_out1;

  Logical_Operator_out7355_out1 <= Logical_Operator_out6331_out1 XOR Logical_Operator_out6395_out1;

  Logical_Operator_out7356_out1 <= Logical_Operator_out6332_out1 XOR Logical_Operator_out6396_out1;

  Logical_Operator_out7357_out1 <= Logical_Operator_out6333_out1 XOR Logical_Operator_out6397_out1;

  Logical_Operator_out7358_out1 <= Logical_Operator_out6334_out1 XOR Logical_Operator_out6398_out1;

  Logical_Operator_out7359_out1 <= Logical_Operator_out6335_out1 XOR Logical_Operator_out6399_out1;

  Logical_Operator_out7360_out1 <= Logical_Operator_out6336_out1 XOR Logical_Operator_out6400_out1;

  Logical_Operator_out7361_out1 <= Logical_Operator_out5281_out1 XOR Logical_Operator_out5345_out1;

  Logical_Operator_out7362_out1 <= Logical_Operator_out5282_out1 XOR Logical_Operator_out5346_out1;

  Logical_Operator_out7363_out1 <= Logical_Operator_out5283_out1 XOR Logical_Operator_out5347_out1;

  Logical_Operator_out7364_out1 <= Logical_Operator_out5284_out1 XOR Logical_Operator_out5348_out1;

  Logical_Operator_out7365_out1 <= Logical_Operator_out5285_out1 XOR Logical_Operator_out5349_out1;

  Logical_Operator_out7366_out1 <= Logical_Operator_out5286_out1 XOR Logical_Operator_out5350_out1;

  Logical_Operator_out7367_out1 <= Logical_Operator_out5287_out1 XOR Logical_Operator_out5351_out1;

  Logical_Operator_out7368_out1 <= Logical_Operator_out5288_out1 XOR Logical_Operator_out5352_out1;

  Logical_Operator_out7369_out1 <= Logical_Operator_out5289_out1 XOR Logical_Operator_out5353_out1;

  Logical_Operator_out7370_out1 <= Logical_Operator_out5290_out1 XOR Logical_Operator_out5354_out1;

  Logical_Operator_out7371_out1 <= Logical_Operator_out5291_out1 XOR Logical_Operator_out5355_out1;

  Logical_Operator_out7372_out1 <= Logical_Operator_out5292_out1 XOR Logical_Operator_out5356_out1;

  Logical_Operator_out7373_out1 <= Logical_Operator_out5293_out1 XOR Logical_Operator_out5357_out1;

  Logical_Operator_out7374_out1 <= Logical_Operator_out5294_out1 XOR Logical_Operator_out5358_out1;

  Logical_Operator_out7375_out1 <= Logical_Operator_out5295_out1 XOR Logical_Operator_out5359_out1;

  Logical_Operator_out7376_out1 <= Logical_Operator_out5296_out1 XOR Logical_Operator_out5360_out1;

  Logical_Operator_out7377_out1 <= Logical_Operator_out5297_out1 XOR Logical_Operator_out5361_out1;

  Logical_Operator_out7378_out1 <= Logical_Operator_out5298_out1 XOR Logical_Operator_out5362_out1;

  Logical_Operator_out7379_out1 <= Logical_Operator_out5299_out1 XOR Logical_Operator_out5363_out1;

  Logical_Operator_out7380_out1 <= Logical_Operator_out5300_out1 XOR Logical_Operator_out5364_out1;

  Logical_Operator_out7381_out1 <= Logical_Operator_out5301_out1 XOR Logical_Operator_out5365_out1;

  Logical_Operator_out7382_out1 <= Logical_Operator_out5302_out1 XOR Logical_Operator_out5366_out1;

  Logical_Operator_out7383_out1 <= Logical_Operator_out5303_out1 XOR Logical_Operator_out5367_out1;

  Logical_Operator_out7384_out1 <= Logical_Operator_out5304_out1 XOR Logical_Operator_out5368_out1;

  Logical_Operator_out7385_out1 <= Logical_Operator_out5305_out1 XOR Logical_Operator_out5369_out1;

  Logical_Operator_out7386_out1 <= Logical_Operator_out5306_out1 XOR Logical_Operator_out5370_out1;

  Logical_Operator_out7387_out1 <= Logical_Operator_out5307_out1 XOR Logical_Operator_out5371_out1;

  Logical_Operator_out7388_out1 <= Logical_Operator_out5308_out1 XOR Logical_Operator_out5372_out1;

  Logical_Operator_out7389_out1 <= Logical_Operator_out5309_out1 XOR Logical_Operator_out5373_out1;

  Logical_Operator_out7390_out1 <= Logical_Operator_out5310_out1 XOR Logical_Operator_out5374_out1;

  Logical_Operator_out7391_out1 <= Logical_Operator_out5311_out1 XOR Logical_Operator_out5375_out1;

  Logical_Operator_out7392_out1 <= Logical_Operator_out5312_out1 XOR Logical_Operator_out5376_out1;

  Logical_Operator_out7393_out1 <= Logical_Operator_out4273_out1 XOR Logical_Operator_out4337_out1;

  Logical_Operator_out7394_out1 <= Logical_Operator_out4274_out1 XOR Logical_Operator_out4338_out1;

  Logical_Operator_out7395_out1 <= Logical_Operator_out4275_out1 XOR Logical_Operator_out4339_out1;

  Logical_Operator_out7396_out1 <= Logical_Operator_out4276_out1 XOR Logical_Operator_out4340_out1;

  Logical_Operator_out7397_out1 <= Logical_Operator_out4277_out1 XOR Logical_Operator_out4341_out1;

  Logical_Operator_out7398_out1 <= Logical_Operator_out4278_out1 XOR Logical_Operator_out4342_out1;

  Logical_Operator_out7399_out1 <= Logical_Operator_out4279_out1 XOR Logical_Operator_out4343_out1;

  Logical_Operator_out7400_out1 <= Logical_Operator_out4280_out1 XOR Logical_Operator_out4344_out1;

  Logical_Operator_out7401_out1 <= Logical_Operator_out4281_out1 XOR Logical_Operator_out4345_out1;

  Logical_Operator_out7402_out1 <= Logical_Operator_out4282_out1 XOR Logical_Operator_out4346_out1;

  Logical_Operator_out7403_out1 <= Logical_Operator_out4283_out1 XOR Logical_Operator_out4347_out1;

  Logical_Operator_out7404_out1 <= Logical_Operator_out4284_out1 XOR Logical_Operator_out4348_out1;

  Logical_Operator_out7405_out1 <= Logical_Operator_out4285_out1 XOR Logical_Operator_out4349_out1;

  Logical_Operator_out7406_out1 <= Logical_Operator_out4286_out1 XOR Logical_Operator_out4350_out1;

  Logical_Operator_out7407_out1 <= Logical_Operator_out4287_out1 XOR Logical_Operator_out4351_out1;

  Logical_Operator_out7408_out1 <= Logical_Operator_out4288_out1 XOR Logical_Operator_out4352_out1;

  Logical_Operator_out7409_out1 <= Logical_Operator_out3257_out1 XOR Logical_Operator_out3321_out1;

  Logical_Operator_out7410_out1 <= Logical_Operator_out3258_out1 XOR Logical_Operator_out3322_out1;

  Logical_Operator_out7411_out1 <= Logical_Operator_out3259_out1 XOR Logical_Operator_out3323_out1;

  Logical_Operator_out7412_out1 <= Logical_Operator_out3260_out1 XOR Logical_Operator_out3324_out1;

  Logical_Operator_out7413_out1 <= Logical_Operator_out3261_out1 XOR Logical_Operator_out3325_out1;

  Logical_Operator_out7414_out1 <= Logical_Operator_out3262_out1 XOR Logical_Operator_out3326_out1;

  Logical_Operator_out7415_out1 <= Logical_Operator_out3263_out1 XOR Logical_Operator_out3327_out1;

  Logical_Operator_out7416_out1 <= Logical_Operator_out3264_out1 XOR Logical_Operator_out3328_out1;

  Logical_Operator_out7417_out1 <= Logical_Operator_out2237_out1 XOR Logical_Operator_out2301_out1;

  Logical_Operator_out7418_out1 <= Logical_Operator_out2238_out1 XOR Logical_Operator_out2302_out1;

  Logical_Operator_out7419_out1 <= Logical_Operator_out2239_out1 XOR Logical_Operator_out2303_out1;

  Logical_Operator_out7420_out1 <= Logical_Operator_out2240_out1 XOR Logical_Operator_out2304_out1;

  Logical_Operator_out7421_out1 <= Logical_Operator_out1215_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out7422_out1 <= Logical_Operator_out1216_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out7423_out1 <= Logical_Operator_out192_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out7424_out1 <= in384 XOR in512;

  Logical_Operator_out7425_out1 <= Logical_Operator_out6401_out1 XOR Logical_Operator_out6465_out1;

  Logical_Operator_out7426_out1 <= Logical_Operator_out6402_out1 XOR Logical_Operator_out6466_out1;

  Logical_Operator_out7427_out1 <= Logical_Operator_out6403_out1 XOR Logical_Operator_out6467_out1;

  Logical_Operator_out7428_out1 <= Logical_Operator_out6404_out1 XOR Logical_Operator_out6468_out1;

  Logical_Operator_out7429_out1 <= Logical_Operator_out6405_out1 XOR Logical_Operator_out6469_out1;

  Logical_Operator_out7430_out1 <= Logical_Operator_out6406_out1 XOR Logical_Operator_out6470_out1;

  Logical_Operator_out7431_out1 <= Logical_Operator_out6407_out1 XOR Logical_Operator_out6471_out1;

  Logical_Operator_out7432_out1 <= Logical_Operator_out6408_out1 XOR Logical_Operator_out6472_out1;

  Logical_Operator_out7433_out1 <= Logical_Operator_out6409_out1 XOR Logical_Operator_out6473_out1;

  Logical_Operator_out7434_out1 <= Logical_Operator_out6410_out1 XOR Logical_Operator_out6474_out1;

  Logical_Operator_out7435_out1 <= Logical_Operator_out6411_out1 XOR Logical_Operator_out6475_out1;

  Logical_Operator_out7436_out1 <= Logical_Operator_out6412_out1 XOR Logical_Operator_out6476_out1;

  Logical_Operator_out7437_out1 <= Logical_Operator_out6413_out1 XOR Logical_Operator_out6477_out1;

  Logical_Operator_out7438_out1 <= Logical_Operator_out6414_out1 XOR Logical_Operator_out6478_out1;

  Logical_Operator_out7439_out1 <= Logical_Operator_out6415_out1 XOR Logical_Operator_out6479_out1;

  Logical_Operator_out7440_out1 <= Logical_Operator_out6416_out1 XOR Logical_Operator_out6480_out1;

  Logical_Operator_out7441_out1 <= Logical_Operator_out6417_out1 XOR Logical_Operator_out6481_out1;

  Logical_Operator_out7442_out1 <= Logical_Operator_out6418_out1 XOR Logical_Operator_out6482_out1;

  Logical_Operator_out7443_out1 <= Logical_Operator_out6419_out1 XOR Logical_Operator_out6483_out1;

  Logical_Operator_out7444_out1 <= Logical_Operator_out6420_out1 XOR Logical_Operator_out6484_out1;

  Logical_Operator_out7445_out1 <= Logical_Operator_out6421_out1 XOR Logical_Operator_out6485_out1;

  Logical_Operator_out7446_out1 <= Logical_Operator_out6422_out1 XOR Logical_Operator_out6486_out1;

  Logical_Operator_out7447_out1 <= Logical_Operator_out6423_out1 XOR Logical_Operator_out6487_out1;

  Logical_Operator_out7448_out1 <= Logical_Operator_out6424_out1 XOR Logical_Operator_out6488_out1;

  Logical_Operator_out7449_out1 <= Logical_Operator_out6425_out1 XOR Logical_Operator_out6489_out1;

  Logical_Operator_out7450_out1 <= Logical_Operator_out6426_out1 XOR Logical_Operator_out6490_out1;

  Logical_Operator_out7451_out1 <= Logical_Operator_out6427_out1 XOR Logical_Operator_out6491_out1;

  Logical_Operator_out7452_out1 <= Logical_Operator_out6428_out1 XOR Logical_Operator_out6492_out1;

  Logical_Operator_out7453_out1 <= Logical_Operator_out6429_out1 XOR Logical_Operator_out6493_out1;

  Logical_Operator_out7454_out1 <= Logical_Operator_out6430_out1 XOR Logical_Operator_out6494_out1;

  Logical_Operator_out7455_out1 <= Logical_Operator_out6431_out1 XOR Logical_Operator_out6495_out1;

  Logical_Operator_out7456_out1 <= Logical_Operator_out6432_out1 XOR Logical_Operator_out6496_out1;

  Logical_Operator_out7457_out1 <= Logical_Operator_out6433_out1 XOR Logical_Operator_out6497_out1;

  Logical_Operator_out7458_out1 <= Logical_Operator_out6434_out1 XOR Logical_Operator_out6498_out1;

  Logical_Operator_out7459_out1 <= Logical_Operator_out6435_out1 XOR Logical_Operator_out6499_out1;

  Logical_Operator_out7460_out1 <= Logical_Operator_out6436_out1 XOR Logical_Operator_out6500_out1;

  Logical_Operator_out7461_out1 <= Logical_Operator_out6437_out1 XOR Logical_Operator_out6501_out1;

  Logical_Operator_out7462_out1 <= Logical_Operator_out6438_out1 XOR Logical_Operator_out6502_out1;

  Logical_Operator_out7463_out1 <= Logical_Operator_out6439_out1 XOR Logical_Operator_out6503_out1;

  Logical_Operator_out7464_out1 <= Logical_Operator_out6440_out1 XOR Logical_Operator_out6504_out1;

  Logical_Operator_out7465_out1 <= Logical_Operator_out6441_out1 XOR Logical_Operator_out6505_out1;

  Logical_Operator_out7466_out1 <= Logical_Operator_out6442_out1 XOR Logical_Operator_out6506_out1;

  Logical_Operator_out7467_out1 <= Logical_Operator_out6443_out1 XOR Logical_Operator_out6507_out1;

  Logical_Operator_out7468_out1 <= Logical_Operator_out6444_out1 XOR Logical_Operator_out6508_out1;

  Logical_Operator_out7469_out1 <= Logical_Operator_out6445_out1 XOR Logical_Operator_out6509_out1;

  Logical_Operator_out7470_out1 <= Logical_Operator_out6446_out1 XOR Logical_Operator_out6510_out1;

  Logical_Operator_out7471_out1 <= Logical_Operator_out6447_out1 XOR Logical_Operator_out6511_out1;

  Logical_Operator_out7472_out1 <= Logical_Operator_out6448_out1 XOR Logical_Operator_out6512_out1;

  Logical_Operator_out7473_out1 <= Logical_Operator_out6449_out1 XOR Logical_Operator_out6513_out1;

  Logical_Operator_out7474_out1 <= Logical_Operator_out6450_out1 XOR Logical_Operator_out6514_out1;

  Logical_Operator_out7475_out1 <= Logical_Operator_out6451_out1 XOR Logical_Operator_out6515_out1;

  Logical_Operator_out7476_out1 <= Logical_Operator_out6452_out1 XOR Logical_Operator_out6516_out1;

  Logical_Operator_out7477_out1 <= Logical_Operator_out6453_out1 XOR Logical_Operator_out6517_out1;

  Logical_Operator_out7478_out1 <= Logical_Operator_out6454_out1 XOR Logical_Operator_out6518_out1;

  Logical_Operator_out7479_out1 <= Logical_Operator_out6455_out1 XOR Logical_Operator_out6519_out1;

  Logical_Operator_out7480_out1 <= Logical_Operator_out6456_out1 XOR Logical_Operator_out6520_out1;

  Logical_Operator_out7481_out1 <= Logical_Operator_out6457_out1 XOR Logical_Operator_out6521_out1;

  Logical_Operator_out7482_out1 <= Logical_Operator_out6458_out1 XOR Logical_Operator_out6522_out1;

  Logical_Operator_out7483_out1 <= Logical_Operator_out6459_out1 XOR Logical_Operator_out6523_out1;

  Logical_Operator_out7484_out1 <= Logical_Operator_out6460_out1 XOR Logical_Operator_out6524_out1;

  Logical_Operator_out7485_out1 <= Logical_Operator_out6461_out1 XOR Logical_Operator_out6525_out1;

  Logical_Operator_out7486_out1 <= Logical_Operator_out6462_out1 XOR Logical_Operator_out6526_out1;

  Logical_Operator_out7487_out1 <= Logical_Operator_out6463_out1 XOR Logical_Operator_out6527_out1;

  Logical_Operator_out7488_out1 <= Logical_Operator_out6464_out1 XOR Logical_Operator_out6528_out1;

  Logical_Operator_out7489_out1 <= Logical_Operator_out5409_out1 XOR Logical_Operator_out5473_out1;

  Logical_Operator_out7490_out1 <= Logical_Operator_out5410_out1 XOR Logical_Operator_out5474_out1;

  Logical_Operator_out7491_out1 <= Logical_Operator_out5411_out1 XOR Logical_Operator_out5475_out1;

  Logical_Operator_out7492_out1 <= Logical_Operator_out5412_out1 XOR Logical_Operator_out5476_out1;

  Logical_Operator_out7493_out1 <= Logical_Operator_out5413_out1 XOR Logical_Operator_out5477_out1;

  Logical_Operator_out7494_out1 <= Logical_Operator_out5414_out1 XOR Logical_Operator_out5478_out1;

  Logical_Operator_out7495_out1 <= Logical_Operator_out5415_out1 XOR Logical_Operator_out5479_out1;

  Logical_Operator_out7496_out1 <= Logical_Operator_out5416_out1 XOR Logical_Operator_out5480_out1;

  Logical_Operator_out7497_out1 <= Logical_Operator_out5417_out1 XOR Logical_Operator_out5481_out1;

  Logical_Operator_out7498_out1 <= Logical_Operator_out5418_out1 XOR Logical_Operator_out5482_out1;

  Logical_Operator_out7499_out1 <= Logical_Operator_out5419_out1 XOR Logical_Operator_out5483_out1;

  Logical_Operator_out7500_out1 <= Logical_Operator_out5420_out1 XOR Logical_Operator_out5484_out1;

  Logical_Operator_out7501_out1 <= Logical_Operator_out5421_out1 XOR Logical_Operator_out5485_out1;

  Logical_Operator_out7502_out1 <= Logical_Operator_out5422_out1 XOR Logical_Operator_out5486_out1;

  Logical_Operator_out7503_out1 <= Logical_Operator_out5423_out1 XOR Logical_Operator_out5487_out1;

  Logical_Operator_out7504_out1 <= Logical_Operator_out5424_out1 XOR Logical_Operator_out5488_out1;

  Logical_Operator_out7505_out1 <= Logical_Operator_out5425_out1 XOR Logical_Operator_out5489_out1;

  Logical_Operator_out7506_out1 <= Logical_Operator_out5426_out1 XOR Logical_Operator_out5490_out1;

  Logical_Operator_out7507_out1 <= Logical_Operator_out5427_out1 XOR Logical_Operator_out5491_out1;

  Logical_Operator_out7508_out1 <= Logical_Operator_out5428_out1 XOR Logical_Operator_out5492_out1;

  Logical_Operator_out7509_out1 <= Logical_Operator_out5429_out1 XOR Logical_Operator_out5493_out1;

  Logical_Operator_out7510_out1 <= Logical_Operator_out5430_out1 XOR Logical_Operator_out5494_out1;

  Logical_Operator_out7511_out1 <= Logical_Operator_out5431_out1 XOR Logical_Operator_out5495_out1;

  Logical_Operator_out7512_out1 <= Logical_Operator_out5432_out1 XOR Logical_Operator_out5496_out1;

  Logical_Operator_out7513_out1 <= Logical_Operator_out5433_out1 XOR Logical_Operator_out5497_out1;

  Logical_Operator_out7514_out1 <= Logical_Operator_out5434_out1 XOR Logical_Operator_out5498_out1;

  Logical_Operator_out7515_out1 <= Logical_Operator_out5435_out1 XOR Logical_Operator_out5499_out1;

  Logical_Operator_out7516_out1 <= Logical_Operator_out5436_out1 XOR Logical_Operator_out5500_out1;

  Logical_Operator_out7517_out1 <= Logical_Operator_out5437_out1 XOR Logical_Operator_out5501_out1;

  Logical_Operator_out7518_out1 <= Logical_Operator_out5438_out1 XOR Logical_Operator_out5502_out1;

  Logical_Operator_out7519_out1 <= Logical_Operator_out5439_out1 XOR Logical_Operator_out5503_out1;

  Logical_Operator_out7520_out1 <= Logical_Operator_out5440_out1 XOR Logical_Operator_out5504_out1;

  Logical_Operator_out7521_out1 <= Logical_Operator_out4401_out1 XOR Logical_Operator_out4465_out1;

  Logical_Operator_out7522_out1 <= Logical_Operator_out4402_out1 XOR Logical_Operator_out4466_out1;

  Logical_Operator_out7523_out1 <= Logical_Operator_out4403_out1 XOR Logical_Operator_out4467_out1;

  Logical_Operator_out7524_out1 <= Logical_Operator_out4404_out1 XOR Logical_Operator_out4468_out1;

  Logical_Operator_out7525_out1 <= Logical_Operator_out4405_out1 XOR Logical_Operator_out4469_out1;

  Logical_Operator_out7526_out1 <= Logical_Operator_out4406_out1 XOR Logical_Operator_out4470_out1;

  Logical_Operator_out7527_out1 <= Logical_Operator_out4407_out1 XOR Logical_Operator_out4471_out1;

  Logical_Operator_out7528_out1 <= Logical_Operator_out4408_out1 XOR Logical_Operator_out4472_out1;

  Logical_Operator_out7529_out1 <= Logical_Operator_out4409_out1 XOR Logical_Operator_out4473_out1;

  Logical_Operator_out7530_out1 <= Logical_Operator_out4410_out1 XOR Logical_Operator_out4474_out1;

  Logical_Operator_out7531_out1 <= Logical_Operator_out4411_out1 XOR Logical_Operator_out4475_out1;

  Logical_Operator_out7532_out1 <= Logical_Operator_out4412_out1 XOR Logical_Operator_out4476_out1;

  Logical_Operator_out7533_out1 <= Logical_Operator_out4413_out1 XOR Logical_Operator_out4477_out1;

  Logical_Operator_out7534_out1 <= Logical_Operator_out4414_out1 XOR Logical_Operator_out4478_out1;

  Logical_Operator_out7535_out1 <= Logical_Operator_out4415_out1 XOR Logical_Operator_out4479_out1;

  Logical_Operator_out7536_out1 <= Logical_Operator_out4416_out1 XOR Logical_Operator_out4480_out1;

  Logical_Operator_out7537_out1 <= Logical_Operator_out3385_out1 XOR Logical_Operator_out3449_out1;

  Logical_Operator_out7538_out1 <= Logical_Operator_out3386_out1 XOR Logical_Operator_out3450_out1;

  Logical_Operator_out7539_out1 <= Logical_Operator_out3387_out1 XOR Logical_Operator_out3451_out1;

  Logical_Operator_out7540_out1 <= Logical_Operator_out3388_out1 XOR Logical_Operator_out3452_out1;

  Logical_Operator_out7541_out1 <= Logical_Operator_out3389_out1 XOR Logical_Operator_out3453_out1;

  Logical_Operator_out7542_out1 <= Logical_Operator_out3390_out1 XOR Logical_Operator_out3454_out1;

  Logical_Operator_out7543_out1 <= Logical_Operator_out3391_out1 XOR Logical_Operator_out3455_out1;

  Logical_Operator_out7544_out1 <= Logical_Operator_out3392_out1 XOR Logical_Operator_out3456_out1;

  Logical_Operator_out7545_out1 <= Logical_Operator_out2365_out1 XOR Logical_Operator_out2429_out1;

  Logical_Operator_out7546_out1 <= Logical_Operator_out2366_out1 XOR Logical_Operator_out2430_out1;

  Logical_Operator_out7547_out1 <= Logical_Operator_out2367_out1 XOR Logical_Operator_out2431_out1;

  Logical_Operator_out7548_out1 <= Logical_Operator_out2368_out1 XOR Logical_Operator_out2432_out1;

  Logical_Operator_out7549_out1 <= Logical_Operator_out1343_out1 XOR Logical_Operator_out1407_out1;

  Logical_Operator_out7550_out1 <= Logical_Operator_out1344_out1 XOR Logical_Operator_out1408_out1;

  Logical_Operator_out7551_out1 <= Logical_Operator_out320_out1 XOR Logical_Operator_out384_out1;

  Logical_Operator_out7552_out1 <= in640 XOR in768;

  Logical_Operator_out7553_out1 <= Logical_Operator_out6529_out1 XOR Logical_Operator_out6593_out1;

  Logical_Operator_out7554_out1 <= Logical_Operator_out6530_out1 XOR Logical_Operator_out6594_out1;

  Logical_Operator_out7555_out1 <= Logical_Operator_out6531_out1 XOR Logical_Operator_out6595_out1;

  Logical_Operator_out7556_out1 <= Logical_Operator_out6532_out1 XOR Logical_Operator_out6596_out1;

  Logical_Operator_out7557_out1 <= Logical_Operator_out6533_out1 XOR Logical_Operator_out6597_out1;

  Logical_Operator_out7558_out1 <= Logical_Operator_out6534_out1 XOR Logical_Operator_out6598_out1;

  Logical_Operator_out7559_out1 <= Logical_Operator_out6535_out1 XOR Logical_Operator_out6599_out1;

  Logical_Operator_out7560_out1 <= Logical_Operator_out6536_out1 XOR Logical_Operator_out6600_out1;

  Logical_Operator_out7561_out1 <= Logical_Operator_out6537_out1 XOR Logical_Operator_out6601_out1;

  Logical_Operator_out7562_out1 <= Logical_Operator_out6538_out1 XOR Logical_Operator_out6602_out1;

  Logical_Operator_out7563_out1 <= Logical_Operator_out6539_out1 XOR Logical_Operator_out6603_out1;

  Logical_Operator_out7564_out1 <= Logical_Operator_out6540_out1 XOR Logical_Operator_out6604_out1;

  Logical_Operator_out7565_out1 <= Logical_Operator_out6541_out1 XOR Logical_Operator_out6605_out1;

  Logical_Operator_out7566_out1 <= Logical_Operator_out6542_out1 XOR Logical_Operator_out6606_out1;

  Logical_Operator_out7567_out1 <= Logical_Operator_out6543_out1 XOR Logical_Operator_out6607_out1;

  Logical_Operator_out7568_out1 <= Logical_Operator_out6544_out1 XOR Logical_Operator_out6608_out1;

  Logical_Operator_out7569_out1 <= Logical_Operator_out6545_out1 XOR Logical_Operator_out6609_out1;

  Logical_Operator_out7570_out1 <= Logical_Operator_out6546_out1 XOR Logical_Operator_out6610_out1;

  Logical_Operator_out7571_out1 <= Logical_Operator_out6547_out1 XOR Logical_Operator_out6611_out1;

  Logical_Operator_out7572_out1 <= Logical_Operator_out6548_out1 XOR Logical_Operator_out6612_out1;

  Logical_Operator_out7573_out1 <= Logical_Operator_out6549_out1 XOR Logical_Operator_out6613_out1;

  Logical_Operator_out7574_out1 <= Logical_Operator_out6550_out1 XOR Logical_Operator_out6614_out1;

  Logical_Operator_out7575_out1 <= Logical_Operator_out6551_out1 XOR Logical_Operator_out6615_out1;

  Logical_Operator_out7576_out1 <= Logical_Operator_out6552_out1 XOR Logical_Operator_out6616_out1;

  Logical_Operator_out7577_out1 <= Logical_Operator_out6553_out1 XOR Logical_Operator_out6617_out1;

  Logical_Operator_out7578_out1 <= Logical_Operator_out6554_out1 XOR Logical_Operator_out6618_out1;

  Logical_Operator_out7579_out1 <= Logical_Operator_out6555_out1 XOR Logical_Operator_out6619_out1;

  Logical_Operator_out7580_out1 <= Logical_Operator_out6556_out1 XOR Logical_Operator_out6620_out1;

  Logical_Operator_out7581_out1 <= Logical_Operator_out6557_out1 XOR Logical_Operator_out6621_out1;

  Logical_Operator_out7582_out1 <= Logical_Operator_out6558_out1 XOR Logical_Operator_out6622_out1;

  Logical_Operator_out7583_out1 <= Logical_Operator_out6559_out1 XOR Logical_Operator_out6623_out1;

  Logical_Operator_out7584_out1 <= Logical_Operator_out6560_out1 XOR Logical_Operator_out6624_out1;

  Logical_Operator_out7585_out1 <= Logical_Operator_out6561_out1 XOR Logical_Operator_out6625_out1;

  Logical_Operator_out7586_out1 <= Logical_Operator_out6562_out1 XOR Logical_Operator_out6626_out1;

  Logical_Operator_out7587_out1 <= Logical_Operator_out6563_out1 XOR Logical_Operator_out6627_out1;

  Logical_Operator_out7588_out1 <= Logical_Operator_out6564_out1 XOR Logical_Operator_out6628_out1;

  Logical_Operator_out7589_out1 <= Logical_Operator_out6565_out1 XOR Logical_Operator_out6629_out1;

  Logical_Operator_out7590_out1 <= Logical_Operator_out6566_out1 XOR Logical_Operator_out6630_out1;

  Logical_Operator_out7591_out1 <= Logical_Operator_out6567_out1 XOR Logical_Operator_out6631_out1;

  Logical_Operator_out7592_out1 <= Logical_Operator_out6568_out1 XOR Logical_Operator_out6632_out1;

  Logical_Operator_out7593_out1 <= Logical_Operator_out6569_out1 XOR Logical_Operator_out6633_out1;

  Logical_Operator_out7594_out1 <= Logical_Operator_out6570_out1 XOR Logical_Operator_out6634_out1;

  Logical_Operator_out7595_out1 <= Logical_Operator_out6571_out1 XOR Logical_Operator_out6635_out1;

  Logical_Operator_out7596_out1 <= Logical_Operator_out6572_out1 XOR Logical_Operator_out6636_out1;

  Logical_Operator_out7597_out1 <= Logical_Operator_out6573_out1 XOR Logical_Operator_out6637_out1;

  Logical_Operator_out7598_out1 <= Logical_Operator_out6574_out1 XOR Logical_Operator_out6638_out1;

  Logical_Operator_out7599_out1 <= Logical_Operator_out6575_out1 XOR Logical_Operator_out6639_out1;

  Logical_Operator_out7600_out1 <= Logical_Operator_out6576_out1 XOR Logical_Operator_out6640_out1;

  Logical_Operator_out7601_out1 <= Logical_Operator_out6577_out1 XOR Logical_Operator_out6641_out1;

  Logical_Operator_out7602_out1 <= Logical_Operator_out6578_out1 XOR Logical_Operator_out6642_out1;

  Logical_Operator_out7603_out1 <= Logical_Operator_out6579_out1 XOR Logical_Operator_out6643_out1;

  Logical_Operator_out7604_out1 <= Logical_Operator_out6580_out1 XOR Logical_Operator_out6644_out1;

  Logical_Operator_out7605_out1 <= Logical_Operator_out6581_out1 XOR Logical_Operator_out6645_out1;

  Logical_Operator_out7606_out1 <= Logical_Operator_out6582_out1 XOR Logical_Operator_out6646_out1;

  Logical_Operator_out7607_out1 <= Logical_Operator_out6583_out1 XOR Logical_Operator_out6647_out1;

  Logical_Operator_out7608_out1 <= Logical_Operator_out6584_out1 XOR Logical_Operator_out6648_out1;

  Logical_Operator_out7609_out1 <= Logical_Operator_out6585_out1 XOR Logical_Operator_out6649_out1;

  Logical_Operator_out7610_out1 <= Logical_Operator_out6586_out1 XOR Logical_Operator_out6650_out1;

  Logical_Operator_out7611_out1 <= Logical_Operator_out6587_out1 XOR Logical_Operator_out6651_out1;

  Logical_Operator_out7612_out1 <= Logical_Operator_out6588_out1 XOR Logical_Operator_out6652_out1;

  Logical_Operator_out7613_out1 <= Logical_Operator_out6589_out1 XOR Logical_Operator_out6653_out1;

  Logical_Operator_out7614_out1 <= Logical_Operator_out6590_out1 XOR Logical_Operator_out6654_out1;

  Logical_Operator_out7615_out1 <= Logical_Operator_out6591_out1 XOR Logical_Operator_out6655_out1;

  Logical_Operator_out7616_out1 <= Logical_Operator_out6592_out1 XOR Logical_Operator_out6656_out1;

  Logical_Operator_out7617_out1 <= Logical_Operator_out5537_out1 XOR Logical_Operator_out5601_out1;

  Logical_Operator_out7618_out1 <= Logical_Operator_out5538_out1 XOR Logical_Operator_out5602_out1;

  Logical_Operator_out7619_out1 <= Logical_Operator_out5539_out1 XOR Logical_Operator_out5603_out1;

  Logical_Operator_out7620_out1 <= Logical_Operator_out5540_out1 XOR Logical_Operator_out5604_out1;

  Logical_Operator_out7621_out1 <= Logical_Operator_out5541_out1 XOR Logical_Operator_out5605_out1;

  Logical_Operator_out7622_out1 <= Logical_Operator_out5542_out1 XOR Logical_Operator_out5606_out1;

  Logical_Operator_out7623_out1 <= Logical_Operator_out5543_out1 XOR Logical_Operator_out5607_out1;

  Logical_Operator_out7624_out1 <= Logical_Operator_out5544_out1 XOR Logical_Operator_out5608_out1;

  Logical_Operator_out7625_out1 <= Logical_Operator_out5545_out1 XOR Logical_Operator_out5609_out1;

  Logical_Operator_out7626_out1 <= Logical_Operator_out5546_out1 XOR Logical_Operator_out5610_out1;

  Logical_Operator_out7627_out1 <= Logical_Operator_out5547_out1 XOR Logical_Operator_out5611_out1;

  Logical_Operator_out7628_out1 <= Logical_Operator_out5548_out1 XOR Logical_Operator_out5612_out1;

  Logical_Operator_out7629_out1 <= Logical_Operator_out5549_out1 XOR Logical_Operator_out5613_out1;

  Logical_Operator_out7630_out1 <= Logical_Operator_out5550_out1 XOR Logical_Operator_out5614_out1;

  Logical_Operator_out7631_out1 <= Logical_Operator_out5551_out1 XOR Logical_Operator_out5615_out1;

  Logical_Operator_out7632_out1 <= Logical_Operator_out5552_out1 XOR Logical_Operator_out5616_out1;

  Logical_Operator_out7633_out1 <= Logical_Operator_out5553_out1 XOR Logical_Operator_out5617_out1;

  Logical_Operator_out7634_out1 <= Logical_Operator_out5554_out1 XOR Logical_Operator_out5618_out1;

  Logical_Operator_out7635_out1 <= Logical_Operator_out5555_out1 XOR Logical_Operator_out5619_out1;

  Logical_Operator_out7636_out1 <= Logical_Operator_out5556_out1 XOR Logical_Operator_out5620_out1;

  Logical_Operator_out7637_out1 <= Logical_Operator_out5557_out1 XOR Logical_Operator_out5621_out1;

  Logical_Operator_out7638_out1 <= Logical_Operator_out5558_out1 XOR Logical_Operator_out5622_out1;

  Logical_Operator_out7639_out1 <= Logical_Operator_out5559_out1 XOR Logical_Operator_out5623_out1;

  Logical_Operator_out7640_out1 <= Logical_Operator_out5560_out1 XOR Logical_Operator_out5624_out1;

  Logical_Operator_out7641_out1 <= Logical_Operator_out5561_out1 XOR Logical_Operator_out5625_out1;

  Logical_Operator_out7642_out1 <= Logical_Operator_out5562_out1 XOR Logical_Operator_out5626_out1;

  Logical_Operator_out7643_out1 <= Logical_Operator_out5563_out1 XOR Logical_Operator_out5627_out1;

  Logical_Operator_out7644_out1 <= Logical_Operator_out5564_out1 XOR Logical_Operator_out5628_out1;

  Logical_Operator_out7645_out1 <= Logical_Operator_out5565_out1 XOR Logical_Operator_out5629_out1;

  Logical_Operator_out7646_out1 <= Logical_Operator_out5566_out1 XOR Logical_Operator_out5630_out1;

  Logical_Operator_out7647_out1 <= Logical_Operator_out5567_out1 XOR Logical_Operator_out5631_out1;

  Logical_Operator_out7648_out1 <= Logical_Operator_out5568_out1 XOR Logical_Operator_out5632_out1;

  Logical_Operator_out7649_out1 <= Logical_Operator_out4529_out1 XOR Logical_Operator_out4593_out1;

  Logical_Operator_out7650_out1 <= Logical_Operator_out4530_out1 XOR Logical_Operator_out4594_out1;

  Logical_Operator_out7651_out1 <= Logical_Operator_out4531_out1 XOR Logical_Operator_out4595_out1;

  Logical_Operator_out7652_out1 <= Logical_Operator_out4532_out1 XOR Logical_Operator_out4596_out1;

  Logical_Operator_out7653_out1 <= Logical_Operator_out4533_out1 XOR Logical_Operator_out4597_out1;

  Logical_Operator_out7654_out1 <= Logical_Operator_out4534_out1 XOR Logical_Operator_out4598_out1;

  Logical_Operator_out7655_out1 <= Logical_Operator_out4535_out1 XOR Logical_Operator_out4599_out1;

  Logical_Operator_out7656_out1 <= Logical_Operator_out4536_out1 XOR Logical_Operator_out4600_out1;

  Logical_Operator_out7657_out1 <= Logical_Operator_out4537_out1 XOR Logical_Operator_out4601_out1;

  Logical_Operator_out7658_out1 <= Logical_Operator_out4538_out1 XOR Logical_Operator_out4602_out1;

  Logical_Operator_out7659_out1 <= Logical_Operator_out4539_out1 XOR Logical_Operator_out4603_out1;

  Logical_Operator_out7660_out1 <= Logical_Operator_out4540_out1 XOR Logical_Operator_out4604_out1;

  Logical_Operator_out7661_out1 <= Logical_Operator_out4541_out1 XOR Logical_Operator_out4605_out1;

  Logical_Operator_out7662_out1 <= Logical_Operator_out4542_out1 XOR Logical_Operator_out4606_out1;

  Logical_Operator_out7663_out1 <= Logical_Operator_out4543_out1 XOR Logical_Operator_out4607_out1;

  Logical_Operator_out7664_out1 <= Logical_Operator_out4544_out1 XOR Logical_Operator_out4608_out1;

  Logical_Operator_out7665_out1 <= Logical_Operator_out3513_out1 XOR Logical_Operator_out3577_out1;

  Logical_Operator_out7666_out1 <= Logical_Operator_out3514_out1 XOR Logical_Operator_out3578_out1;

  Logical_Operator_out7667_out1 <= Logical_Operator_out3515_out1 XOR Logical_Operator_out3579_out1;

  Logical_Operator_out7668_out1 <= Logical_Operator_out3516_out1 XOR Logical_Operator_out3580_out1;

  Logical_Operator_out7669_out1 <= Logical_Operator_out3517_out1 XOR Logical_Operator_out3581_out1;

  Logical_Operator_out7670_out1 <= Logical_Operator_out3518_out1 XOR Logical_Operator_out3582_out1;

  Logical_Operator_out7671_out1 <= Logical_Operator_out3519_out1 XOR Logical_Operator_out3583_out1;

  Logical_Operator_out7672_out1 <= Logical_Operator_out3520_out1 XOR Logical_Operator_out3584_out1;

  Logical_Operator_out7673_out1 <= Logical_Operator_out2493_out1 XOR Logical_Operator_out2557_out1;

  Logical_Operator_out7674_out1 <= Logical_Operator_out2494_out1 XOR Logical_Operator_out2558_out1;

  Logical_Operator_out7675_out1 <= Logical_Operator_out2495_out1 XOR Logical_Operator_out2559_out1;

  Logical_Operator_out7676_out1 <= Logical_Operator_out2496_out1 XOR Logical_Operator_out2560_out1;

  Logical_Operator_out7677_out1 <= Logical_Operator_out1471_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out7678_out1 <= Logical_Operator_out1472_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out7679_out1 <= Logical_Operator_out448_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out7680_out1 <= in896 XOR in1024;

  Logical_Operator_out7681_out1 <= Logical_Operator_out6657_out1 XOR Logical_Operator_out6721_out1;

  Logical_Operator_out7682_out1 <= Logical_Operator_out6658_out1 XOR Logical_Operator_out6722_out1;

  Logical_Operator_out7683_out1 <= Logical_Operator_out6659_out1 XOR Logical_Operator_out6723_out1;

  Logical_Operator_out7684_out1 <= Logical_Operator_out6660_out1 XOR Logical_Operator_out6724_out1;

  Logical_Operator_out7685_out1 <= Logical_Operator_out6661_out1 XOR Logical_Operator_out6725_out1;

  Logical_Operator_out7686_out1 <= Logical_Operator_out6662_out1 XOR Logical_Operator_out6726_out1;

  Logical_Operator_out7687_out1 <= Logical_Operator_out6663_out1 XOR Logical_Operator_out6727_out1;

  Logical_Operator_out7688_out1 <= Logical_Operator_out6664_out1 XOR Logical_Operator_out6728_out1;

  Logical_Operator_out7689_out1 <= Logical_Operator_out6665_out1 XOR Logical_Operator_out6729_out1;

  Logical_Operator_out7690_out1 <= Logical_Operator_out6666_out1 XOR Logical_Operator_out6730_out1;

  Logical_Operator_out7691_out1 <= Logical_Operator_out6667_out1 XOR Logical_Operator_out6731_out1;

  Logical_Operator_out7692_out1 <= Logical_Operator_out6668_out1 XOR Logical_Operator_out6732_out1;

  Logical_Operator_out7693_out1 <= Logical_Operator_out6669_out1 XOR Logical_Operator_out6733_out1;

  Logical_Operator_out7694_out1 <= Logical_Operator_out6670_out1 XOR Logical_Operator_out6734_out1;

  Logical_Operator_out7695_out1 <= Logical_Operator_out6671_out1 XOR Logical_Operator_out6735_out1;

  Logical_Operator_out7696_out1 <= Logical_Operator_out6672_out1 XOR Logical_Operator_out6736_out1;

  Logical_Operator_out7697_out1 <= Logical_Operator_out6673_out1 XOR Logical_Operator_out6737_out1;

  Logical_Operator_out7698_out1 <= Logical_Operator_out6674_out1 XOR Logical_Operator_out6738_out1;

  Logical_Operator_out7699_out1 <= Logical_Operator_out6675_out1 XOR Logical_Operator_out6739_out1;

  Logical_Operator_out7700_out1 <= Logical_Operator_out6676_out1 XOR Logical_Operator_out6740_out1;

  Logical_Operator_out7701_out1 <= Logical_Operator_out6677_out1 XOR Logical_Operator_out6741_out1;

  Logical_Operator_out7702_out1 <= Logical_Operator_out6678_out1 XOR Logical_Operator_out6742_out1;

  Logical_Operator_out7703_out1 <= Logical_Operator_out6679_out1 XOR Logical_Operator_out6743_out1;

  Logical_Operator_out7704_out1 <= Logical_Operator_out6680_out1 XOR Logical_Operator_out6744_out1;

  Logical_Operator_out7705_out1 <= Logical_Operator_out6681_out1 XOR Logical_Operator_out6745_out1;

  Logical_Operator_out7706_out1 <= Logical_Operator_out6682_out1 XOR Logical_Operator_out6746_out1;

  Logical_Operator_out7707_out1 <= Logical_Operator_out6683_out1 XOR Logical_Operator_out6747_out1;

  Logical_Operator_out7708_out1 <= Logical_Operator_out6684_out1 XOR Logical_Operator_out6748_out1;

  Logical_Operator_out7709_out1 <= Logical_Operator_out6685_out1 XOR Logical_Operator_out6749_out1;

  Logical_Operator_out7710_out1 <= Logical_Operator_out6686_out1 XOR Logical_Operator_out6750_out1;

  Logical_Operator_out7711_out1 <= Logical_Operator_out6687_out1 XOR Logical_Operator_out6751_out1;

  Logical_Operator_out7712_out1 <= Logical_Operator_out6688_out1 XOR Logical_Operator_out6752_out1;

  Logical_Operator_out7713_out1 <= Logical_Operator_out6689_out1 XOR Logical_Operator_out6753_out1;

  Logical_Operator_out7714_out1 <= Logical_Operator_out6690_out1 XOR Logical_Operator_out6754_out1;

  Logical_Operator_out7715_out1 <= Logical_Operator_out6691_out1 XOR Logical_Operator_out6755_out1;

  Logical_Operator_out7716_out1 <= Logical_Operator_out6692_out1 XOR Logical_Operator_out6756_out1;

  Logical_Operator_out7717_out1 <= Logical_Operator_out6693_out1 XOR Logical_Operator_out6757_out1;

  Logical_Operator_out7718_out1 <= Logical_Operator_out6694_out1 XOR Logical_Operator_out6758_out1;

  Logical_Operator_out7719_out1 <= Logical_Operator_out6695_out1 XOR Logical_Operator_out6759_out1;

  Logical_Operator_out7720_out1 <= Logical_Operator_out6696_out1 XOR Logical_Operator_out6760_out1;

  Logical_Operator_out7721_out1 <= Logical_Operator_out6697_out1 XOR Logical_Operator_out6761_out1;

  Logical_Operator_out7722_out1 <= Logical_Operator_out6698_out1 XOR Logical_Operator_out6762_out1;

  Logical_Operator_out7723_out1 <= Logical_Operator_out6699_out1 XOR Logical_Operator_out6763_out1;

  Logical_Operator_out7724_out1 <= Logical_Operator_out6700_out1 XOR Logical_Operator_out6764_out1;

  Logical_Operator_out7725_out1 <= Logical_Operator_out6701_out1 XOR Logical_Operator_out6765_out1;

  Logical_Operator_out7726_out1 <= Logical_Operator_out6702_out1 XOR Logical_Operator_out6766_out1;

  Logical_Operator_out7727_out1 <= Logical_Operator_out6703_out1 XOR Logical_Operator_out6767_out1;

  Logical_Operator_out7728_out1 <= Logical_Operator_out6704_out1 XOR Logical_Operator_out6768_out1;

  Logical_Operator_out7729_out1 <= Logical_Operator_out6705_out1 XOR Logical_Operator_out6769_out1;

  Logical_Operator_out7730_out1 <= Logical_Operator_out6706_out1 XOR Logical_Operator_out6770_out1;

  Logical_Operator_out7731_out1 <= Logical_Operator_out6707_out1 XOR Logical_Operator_out6771_out1;

  Logical_Operator_out7732_out1 <= Logical_Operator_out6708_out1 XOR Logical_Operator_out6772_out1;

  Logical_Operator_out7733_out1 <= Logical_Operator_out6709_out1 XOR Logical_Operator_out6773_out1;

  Logical_Operator_out7734_out1 <= Logical_Operator_out6710_out1 XOR Logical_Operator_out6774_out1;

  Logical_Operator_out7735_out1 <= Logical_Operator_out6711_out1 XOR Logical_Operator_out6775_out1;

  Logical_Operator_out7736_out1 <= Logical_Operator_out6712_out1 XOR Logical_Operator_out6776_out1;

  Logical_Operator_out7737_out1 <= Logical_Operator_out6713_out1 XOR Logical_Operator_out6777_out1;

  Logical_Operator_out7738_out1 <= Logical_Operator_out6714_out1 XOR Logical_Operator_out6778_out1;

  Logical_Operator_out7739_out1 <= Logical_Operator_out6715_out1 XOR Logical_Operator_out6779_out1;

  Logical_Operator_out7740_out1 <= Logical_Operator_out6716_out1 XOR Logical_Operator_out6780_out1;

  Logical_Operator_out7741_out1 <= Logical_Operator_out6717_out1 XOR Logical_Operator_out6781_out1;

  Logical_Operator_out7742_out1 <= Logical_Operator_out6718_out1 XOR Logical_Operator_out6782_out1;

  Logical_Operator_out7743_out1 <= Logical_Operator_out6719_out1 XOR Logical_Operator_out6783_out1;

  Logical_Operator_out7744_out1 <= Logical_Operator_out6720_out1 XOR Logical_Operator_out6784_out1;

  Logical_Operator_out7745_out1 <= Logical_Operator_out5665_out1 XOR Logical_Operator_out5729_out1;

  Logical_Operator_out7746_out1 <= Logical_Operator_out5666_out1 XOR Logical_Operator_out5730_out1;

  Logical_Operator_out7747_out1 <= Logical_Operator_out5667_out1 XOR Logical_Operator_out5731_out1;

  Logical_Operator_out7748_out1 <= Logical_Operator_out5668_out1 XOR Logical_Operator_out5732_out1;

  Logical_Operator_out7749_out1 <= Logical_Operator_out5669_out1 XOR Logical_Operator_out5733_out1;

  Logical_Operator_out7750_out1 <= Logical_Operator_out5670_out1 XOR Logical_Operator_out5734_out1;

  Logical_Operator_out7751_out1 <= Logical_Operator_out5671_out1 XOR Logical_Operator_out5735_out1;

  Logical_Operator_out7752_out1 <= Logical_Operator_out5672_out1 XOR Logical_Operator_out5736_out1;

  Logical_Operator_out7753_out1 <= Logical_Operator_out5673_out1 XOR Logical_Operator_out5737_out1;

  Logical_Operator_out7754_out1 <= Logical_Operator_out5674_out1 XOR Logical_Operator_out5738_out1;

  Logical_Operator_out7755_out1 <= Logical_Operator_out5675_out1 XOR Logical_Operator_out5739_out1;

  Logical_Operator_out7756_out1 <= Logical_Operator_out5676_out1 XOR Logical_Operator_out5740_out1;

  Logical_Operator_out7757_out1 <= Logical_Operator_out5677_out1 XOR Logical_Operator_out5741_out1;

  Logical_Operator_out7758_out1 <= Logical_Operator_out5678_out1 XOR Logical_Operator_out5742_out1;

  Logical_Operator_out7759_out1 <= Logical_Operator_out5679_out1 XOR Logical_Operator_out5743_out1;

  Logical_Operator_out7760_out1 <= Logical_Operator_out5680_out1 XOR Logical_Operator_out5744_out1;

  Logical_Operator_out7761_out1 <= Logical_Operator_out5681_out1 XOR Logical_Operator_out5745_out1;

  Logical_Operator_out7762_out1 <= Logical_Operator_out5682_out1 XOR Logical_Operator_out5746_out1;

  Logical_Operator_out7763_out1 <= Logical_Operator_out5683_out1 XOR Logical_Operator_out5747_out1;

  Logical_Operator_out7764_out1 <= Logical_Operator_out5684_out1 XOR Logical_Operator_out5748_out1;

  Logical_Operator_out7765_out1 <= Logical_Operator_out5685_out1 XOR Logical_Operator_out5749_out1;

  Logical_Operator_out7766_out1 <= Logical_Operator_out5686_out1 XOR Logical_Operator_out5750_out1;

  Logical_Operator_out7767_out1 <= Logical_Operator_out5687_out1 XOR Logical_Operator_out5751_out1;

  Logical_Operator_out7768_out1 <= Logical_Operator_out5688_out1 XOR Logical_Operator_out5752_out1;

  Logical_Operator_out7769_out1 <= Logical_Operator_out5689_out1 XOR Logical_Operator_out5753_out1;

  Logical_Operator_out7770_out1 <= Logical_Operator_out5690_out1 XOR Logical_Operator_out5754_out1;

  Logical_Operator_out7771_out1 <= Logical_Operator_out5691_out1 XOR Logical_Operator_out5755_out1;

  Logical_Operator_out7772_out1 <= Logical_Operator_out5692_out1 XOR Logical_Operator_out5756_out1;

  Logical_Operator_out7773_out1 <= Logical_Operator_out5693_out1 XOR Logical_Operator_out5757_out1;

  Logical_Operator_out7774_out1 <= Logical_Operator_out5694_out1 XOR Logical_Operator_out5758_out1;

  Logical_Operator_out7775_out1 <= Logical_Operator_out5695_out1 XOR Logical_Operator_out5759_out1;

  Logical_Operator_out7776_out1 <= Logical_Operator_out5696_out1 XOR Logical_Operator_out5760_out1;

  Logical_Operator_out7777_out1 <= Logical_Operator_out4657_out1 XOR Logical_Operator_out4721_out1;

  Logical_Operator_out7778_out1 <= Logical_Operator_out4658_out1 XOR Logical_Operator_out4722_out1;

  Logical_Operator_out7779_out1 <= Logical_Operator_out4659_out1 XOR Logical_Operator_out4723_out1;

  Logical_Operator_out7780_out1 <= Logical_Operator_out4660_out1 XOR Logical_Operator_out4724_out1;

  Logical_Operator_out7781_out1 <= Logical_Operator_out4661_out1 XOR Logical_Operator_out4725_out1;

  Logical_Operator_out7782_out1 <= Logical_Operator_out4662_out1 XOR Logical_Operator_out4726_out1;

  Logical_Operator_out7783_out1 <= Logical_Operator_out4663_out1 XOR Logical_Operator_out4727_out1;

  Logical_Operator_out7784_out1 <= Logical_Operator_out4664_out1 XOR Logical_Operator_out4728_out1;

  Logical_Operator_out7785_out1 <= Logical_Operator_out4665_out1 XOR Logical_Operator_out4729_out1;

  Logical_Operator_out7786_out1 <= Logical_Operator_out4666_out1 XOR Logical_Operator_out4730_out1;

  Logical_Operator_out7787_out1 <= Logical_Operator_out4667_out1 XOR Logical_Operator_out4731_out1;

  Logical_Operator_out7788_out1 <= Logical_Operator_out4668_out1 XOR Logical_Operator_out4732_out1;

  Logical_Operator_out7789_out1 <= Logical_Operator_out4669_out1 XOR Logical_Operator_out4733_out1;

  Logical_Operator_out7790_out1 <= Logical_Operator_out4670_out1 XOR Logical_Operator_out4734_out1;

  Logical_Operator_out7791_out1 <= Logical_Operator_out4671_out1 XOR Logical_Operator_out4735_out1;

  Logical_Operator_out7792_out1 <= Logical_Operator_out4672_out1 XOR Logical_Operator_out4736_out1;

  Logical_Operator_out7793_out1 <= Logical_Operator_out3641_out1 XOR Logical_Operator_out3705_out1;

  Logical_Operator_out7794_out1 <= Logical_Operator_out3642_out1 XOR Logical_Operator_out3706_out1;

  Logical_Operator_out7795_out1 <= Logical_Operator_out3643_out1 XOR Logical_Operator_out3707_out1;

  Logical_Operator_out7796_out1 <= Logical_Operator_out3644_out1 XOR Logical_Operator_out3708_out1;

  Logical_Operator_out7797_out1 <= Logical_Operator_out3645_out1 XOR Logical_Operator_out3709_out1;

  Logical_Operator_out7798_out1 <= Logical_Operator_out3646_out1 XOR Logical_Operator_out3710_out1;

  Logical_Operator_out7799_out1 <= Logical_Operator_out3647_out1 XOR Logical_Operator_out3711_out1;

  Logical_Operator_out7800_out1 <= Logical_Operator_out3648_out1 XOR Logical_Operator_out3712_out1;

  Logical_Operator_out7801_out1 <= Logical_Operator_out2621_out1 XOR Logical_Operator_out2685_out1;

  Logical_Operator_out7802_out1 <= Logical_Operator_out2622_out1 XOR Logical_Operator_out2686_out1;

  Logical_Operator_out7803_out1 <= Logical_Operator_out2623_out1 XOR Logical_Operator_out2687_out1;

  Logical_Operator_out7804_out1 <= Logical_Operator_out2624_out1 XOR Logical_Operator_out2688_out1;

  Logical_Operator_out7805_out1 <= Logical_Operator_out1599_out1 XOR Logical_Operator_out1663_out1;

  Logical_Operator_out7806_out1 <= Logical_Operator_out1600_out1 XOR Logical_Operator_out1664_out1;

  Logical_Operator_out7807_out1 <= Logical_Operator_out576_out1 XOR Logical_Operator_out640_out1;

  Logical_Operator_out7808_out1 <= in1152 XOR in1280;

  Logical_Operator_out7809_out1 <= Logical_Operator_out6785_out1 XOR Logical_Operator_out6849_out1;

  Logical_Operator_out7810_out1 <= Logical_Operator_out6786_out1 XOR Logical_Operator_out6850_out1;

  Logical_Operator_out7811_out1 <= Logical_Operator_out6787_out1 XOR Logical_Operator_out6851_out1;

  Logical_Operator_out7812_out1 <= Logical_Operator_out6788_out1 XOR Logical_Operator_out6852_out1;

  Logical_Operator_out7813_out1 <= Logical_Operator_out6789_out1 XOR Logical_Operator_out6853_out1;

  Logical_Operator_out7814_out1 <= Logical_Operator_out6790_out1 XOR Logical_Operator_out6854_out1;

  Logical_Operator_out7815_out1 <= Logical_Operator_out6791_out1 XOR Logical_Operator_out6855_out1;

  Logical_Operator_out7816_out1 <= Logical_Operator_out6792_out1 XOR Logical_Operator_out6856_out1;

  Logical_Operator_out7817_out1 <= Logical_Operator_out6793_out1 XOR Logical_Operator_out6857_out1;

  Logical_Operator_out7818_out1 <= Logical_Operator_out6794_out1 XOR Logical_Operator_out6858_out1;

  Logical_Operator_out7819_out1 <= Logical_Operator_out6795_out1 XOR Logical_Operator_out6859_out1;

  Logical_Operator_out7820_out1 <= Logical_Operator_out6796_out1 XOR Logical_Operator_out6860_out1;

  Logical_Operator_out7821_out1 <= Logical_Operator_out6797_out1 XOR Logical_Operator_out6861_out1;

  Logical_Operator_out7822_out1 <= Logical_Operator_out6798_out1 XOR Logical_Operator_out6862_out1;

  Logical_Operator_out7823_out1 <= Logical_Operator_out6799_out1 XOR Logical_Operator_out6863_out1;

  Logical_Operator_out7824_out1 <= Logical_Operator_out6800_out1 XOR Logical_Operator_out6864_out1;

  Logical_Operator_out7825_out1 <= Logical_Operator_out6801_out1 XOR Logical_Operator_out6865_out1;

  Logical_Operator_out7826_out1 <= Logical_Operator_out6802_out1 XOR Logical_Operator_out6866_out1;

  Logical_Operator_out7827_out1 <= Logical_Operator_out6803_out1 XOR Logical_Operator_out6867_out1;

  Logical_Operator_out7828_out1 <= Logical_Operator_out6804_out1 XOR Logical_Operator_out6868_out1;

  Logical_Operator_out7829_out1 <= Logical_Operator_out6805_out1 XOR Logical_Operator_out6869_out1;

  Logical_Operator_out7830_out1 <= Logical_Operator_out6806_out1 XOR Logical_Operator_out6870_out1;

  Logical_Operator_out7831_out1 <= Logical_Operator_out6807_out1 XOR Logical_Operator_out6871_out1;

  Logical_Operator_out7832_out1 <= Logical_Operator_out6808_out1 XOR Logical_Operator_out6872_out1;

  Logical_Operator_out7833_out1 <= Logical_Operator_out6809_out1 XOR Logical_Operator_out6873_out1;

  Logical_Operator_out7834_out1 <= Logical_Operator_out6810_out1 XOR Logical_Operator_out6874_out1;

  Logical_Operator_out7835_out1 <= Logical_Operator_out6811_out1 XOR Logical_Operator_out6875_out1;

  Logical_Operator_out7836_out1 <= Logical_Operator_out6812_out1 XOR Logical_Operator_out6876_out1;

  Logical_Operator_out7837_out1 <= Logical_Operator_out6813_out1 XOR Logical_Operator_out6877_out1;

  Logical_Operator_out7838_out1 <= Logical_Operator_out6814_out1 XOR Logical_Operator_out6878_out1;

  Logical_Operator_out7839_out1 <= Logical_Operator_out6815_out1 XOR Logical_Operator_out6879_out1;

  Logical_Operator_out7840_out1 <= Logical_Operator_out6816_out1 XOR Logical_Operator_out6880_out1;

  Logical_Operator_out7841_out1 <= Logical_Operator_out6817_out1 XOR Logical_Operator_out6881_out1;

  Logical_Operator_out7842_out1 <= Logical_Operator_out6818_out1 XOR Logical_Operator_out6882_out1;

  Logical_Operator_out7843_out1 <= Logical_Operator_out6819_out1 XOR Logical_Operator_out6883_out1;

  Logical_Operator_out7844_out1 <= Logical_Operator_out6820_out1 XOR Logical_Operator_out6884_out1;

  Logical_Operator_out7845_out1 <= Logical_Operator_out6821_out1 XOR Logical_Operator_out6885_out1;

  Logical_Operator_out7846_out1 <= Logical_Operator_out6822_out1 XOR Logical_Operator_out6886_out1;

  Logical_Operator_out7847_out1 <= Logical_Operator_out6823_out1 XOR Logical_Operator_out6887_out1;

  Logical_Operator_out7848_out1 <= Logical_Operator_out6824_out1 XOR Logical_Operator_out6888_out1;

  Logical_Operator_out7849_out1 <= Logical_Operator_out6825_out1 XOR Logical_Operator_out6889_out1;

  Logical_Operator_out7850_out1 <= Logical_Operator_out6826_out1 XOR Logical_Operator_out6890_out1;

  Logical_Operator_out7851_out1 <= Logical_Operator_out6827_out1 XOR Logical_Operator_out6891_out1;

  Logical_Operator_out7852_out1 <= Logical_Operator_out6828_out1 XOR Logical_Operator_out6892_out1;

  Logical_Operator_out7853_out1 <= Logical_Operator_out6829_out1 XOR Logical_Operator_out6893_out1;

  Logical_Operator_out7854_out1 <= Logical_Operator_out6830_out1 XOR Logical_Operator_out6894_out1;

  Logical_Operator_out7855_out1 <= Logical_Operator_out6831_out1 XOR Logical_Operator_out6895_out1;

  Logical_Operator_out7856_out1 <= Logical_Operator_out6832_out1 XOR Logical_Operator_out6896_out1;

  Logical_Operator_out7857_out1 <= Logical_Operator_out6833_out1 XOR Logical_Operator_out6897_out1;

  Logical_Operator_out7858_out1 <= Logical_Operator_out6834_out1 XOR Logical_Operator_out6898_out1;

  Logical_Operator_out7859_out1 <= Logical_Operator_out6835_out1 XOR Logical_Operator_out6899_out1;

  Logical_Operator_out7860_out1 <= Logical_Operator_out6836_out1 XOR Logical_Operator_out6900_out1;

  Logical_Operator_out7861_out1 <= Logical_Operator_out6837_out1 XOR Logical_Operator_out6901_out1;

  Logical_Operator_out7862_out1 <= Logical_Operator_out6838_out1 XOR Logical_Operator_out6902_out1;

  Logical_Operator_out7863_out1 <= Logical_Operator_out6839_out1 XOR Logical_Operator_out6903_out1;

  Logical_Operator_out7864_out1 <= Logical_Operator_out6840_out1 XOR Logical_Operator_out6904_out1;

  Logical_Operator_out7865_out1 <= Logical_Operator_out6841_out1 XOR Logical_Operator_out6905_out1;

  Logical_Operator_out7866_out1 <= Logical_Operator_out6842_out1 XOR Logical_Operator_out6906_out1;

  Logical_Operator_out7867_out1 <= Logical_Operator_out6843_out1 XOR Logical_Operator_out6907_out1;

  Logical_Operator_out7868_out1 <= Logical_Operator_out6844_out1 XOR Logical_Operator_out6908_out1;

  Logical_Operator_out7869_out1 <= Logical_Operator_out6845_out1 XOR Logical_Operator_out6909_out1;

  Logical_Operator_out7870_out1 <= Logical_Operator_out6846_out1 XOR Logical_Operator_out6910_out1;

  Logical_Operator_out7871_out1 <= Logical_Operator_out6847_out1 XOR Logical_Operator_out6911_out1;

  Logical_Operator_out7872_out1 <= Logical_Operator_out6848_out1 XOR Logical_Operator_out6912_out1;

  Logical_Operator_out7873_out1 <= Logical_Operator_out5793_out1 XOR Logical_Operator_out5857_out1;

  Logical_Operator_out7874_out1 <= Logical_Operator_out5794_out1 XOR Logical_Operator_out5858_out1;

  Logical_Operator_out7875_out1 <= Logical_Operator_out5795_out1 XOR Logical_Operator_out5859_out1;

  Logical_Operator_out7876_out1 <= Logical_Operator_out5796_out1 XOR Logical_Operator_out5860_out1;

  Logical_Operator_out7877_out1 <= Logical_Operator_out5797_out1 XOR Logical_Operator_out5861_out1;

  Logical_Operator_out7878_out1 <= Logical_Operator_out5798_out1 XOR Logical_Operator_out5862_out1;

  Logical_Operator_out7879_out1 <= Logical_Operator_out5799_out1 XOR Logical_Operator_out5863_out1;

  Logical_Operator_out7880_out1 <= Logical_Operator_out5800_out1 XOR Logical_Operator_out5864_out1;

  Logical_Operator_out7881_out1 <= Logical_Operator_out5801_out1 XOR Logical_Operator_out5865_out1;

  Logical_Operator_out7882_out1 <= Logical_Operator_out5802_out1 XOR Logical_Operator_out5866_out1;

  Logical_Operator_out7883_out1 <= Logical_Operator_out5803_out1 XOR Logical_Operator_out5867_out1;

  Logical_Operator_out7884_out1 <= Logical_Operator_out5804_out1 XOR Logical_Operator_out5868_out1;

  Logical_Operator_out7885_out1 <= Logical_Operator_out5805_out1 XOR Logical_Operator_out5869_out1;

  Logical_Operator_out7886_out1 <= Logical_Operator_out5806_out1 XOR Logical_Operator_out5870_out1;

  Logical_Operator_out7887_out1 <= Logical_Operator_out5807_out1 XOR Logical_Operator_out5871_out1;

  Logical_Operator_out7888_out1 <= Logical_Operator_out5808_out1 XOR Logical_Operator_out5872_out1;

  Logical_Operator_out7889_out1 <= Logical_Operator_out5809_out1 XOR Logical_Operator_out5873_out1;

  Logical_Operator_out7890_out1 <= Logical_Operator_out5810_out1 XOR Logical_Operator_out5874_out1;

  Logical_Operator_out7891_out1 <= Logical_Operator_out5811_out1 XOR Logical_Operator_out5875_out1;

  Logical_Operator_out7892_out1 <= Logical_Operator_out5812_out1 XOR Logical_Operator_out5876_out1;

  Logical_Operator_out7893_out1 <= Logical_Operator_out5813_out1 XOR Logical_Operator_out5877_out1;

  Logical_Operator_out7894_out1 <= Logical_Operator_out5814_out1 XOR Logical_Operator_out5878_out1;

  Logical_Operator_out7895_out1 <= Logical_Operator_out5815_out1 XOR Logical_Operator_out5879_out1;

  Logical_Operator_out7896_out1 <= Logical_Operator_out5816_out1 XOR Logical_Operator_out5880_out1;

  Logical_Operator_out7897_out1 <= Logical_Operator_out5817_out1 XOR Logical_Operator_out5881_out1;

  Logical_Operator_out7898_out1 <= Logical_Operator_out5818_out1 XOR Logical_Operator_out5882_out1;

  Logical_Operator_out7899_out1 <= Logical_Operator_out5819_out1 XOR Logical_Operator_out5883_out1;

  Logical_Operator_out7900_out1 <= Logical_Operator_out5820_out1 XOR Logical_Operator_out5884_out1;

  Logical_Operator_out7901_out1 <= Logical_Operator_out5821_out1 XOR Logical_Operator_out5885_out1;

  Logical_Operator_out7902_out1 <= Logical_Operator_out5822_out1 XOR Logical_Operator_out5886_out1;

  Logical_Operator_out7903_out1 <= Logical_Operator_out5823_out1 XOR Logical_Operator_out5887_out1;

  Logical_Operator_out7904_out1 <= Logical_Operator_out5824_out1 XOR Logical_Operator_out5888_out1;

  Logical_Operator_out7905_out1 <= Logical_Operator_out4785_out1 XOR Logical_Operator_out4849_out1;

  Logical_Operator_out7906_out1 <= Logical_Operator_out4786_out1 XOR Logical_Operator_out4850_out1;

  Logical_Operator_out7907_out1 <= Logical_Operator_out4787_out1 XOR Logical_Operator_out4851_out1;

  Logical_Operator_out7908_out1 <= Logical_Operator_out4788_out1 XOR Logical_Operator_out4852_out1;

  Logical_Operator_out7909_out1 <= Logical_Operator_out4789_out1 XOR Logical_Operator_out4853_out1;

  Logical_Operator_out7910_out1 <= Logical_Operator_out4790_out1 XOR Logical_Operator_out4854_out1;

  Logical_Operator_out7911_out1 <= Logical_Operator_out4791_out1 XOR Logical_Operator_out4855_out1;

  Logical_Operator_out7912_out1 <= Logical_Operator_out4792_out1 XOR Logical_Operator_out4856_out1;

  Logical_Operator_out7913_out1 <= Logical_Operator_out4793_out1 XOR Logical_Operator_out4857_out1;

  Logical_Operator_out7914_out1 <= Logical_Operator_out4794_out1 XOR Logical_Operator_out4858_out1;

  Logical_Operator_out7915_out1 <= Logical_Operator_out4795_out1 XOR Logical_Operator_out4859_out1;

  Logical_Operator_out7916_out1 <= Logical_Operator_out4796_out1 XOR Logical_Operator_out4860_out1;

  Logical_Operator_out7917_out1 <= Logical_Operator_out4797_out1 XOR Logical_Operator_out4861_out1;

  Logical_Operator_out7918_out1 <= Logical_Operator_out4798_out1 XOR Logical_Operator_out4862_out1;

  Logical_Operator_out7919_out1 <= Logical_Operator_out4799_out1 XOR Logical_Operator_out4863_out1;

  Logical_Operator_out7920_out1 <= Logical_Operator_out4800_out1 XOR Logical_Operator_out4864_out1;

  Logical_Operator_out7921_out1 <= Logical_Operator_out3769_out1 XOR Logical_Operator_out3833_out1;

  Logical_Operator_out7922_out1 <= Logical_Operator_out3770_out1 XOR Logical_Operator_out3834_out1;

  Logical_Operator_out7923_out1 <= Logical_Operator_out3771_out1 XOR Logical_Operator_out3835_out1;

  Logical_Operator_out7924_out1 <= Logical_Operator_out3772_out1 XOR Logical_Operator_out3836_out1;

  Logical_Operator_out7925_out1 <= Logical_Operator_out3773_out1 XOR Logical_Operator_out3837_out1;

  Logical_Operator_out7926_out1 <= Logical_Operator_out3774_out1 XOR Logical_Operator_out3838_out1;

  Logical_Operator_out7927_out1 <= Logical_Operator_out3775_out1 XOR Logical_Operator_out3839_out1;

  Logical_Operator_out7928_out1 <= Logical_Operator_out3776_out1 XOR Logical_Operator_out3840_out1;

  Logical_Operator_out7929_out1 <= Logical_Operator_out2749_out1 XOR Logical_Operator_out2813_out1;

  Logical_Operator_out7930_out1 <= Logical_Operator_out2750_out1 XOR Logical_Operator_out2814_out1;

  Logical_Operator_out7931_out1 <= Logical_Operator_out2751_out1 XOR Logical_Operator_out2815_out1;

  Logical_Operator_out7932_out1 <= Logical_Operator_out2752_out1 XOR Logical_Operator_out2816_out1;

  Logical_Operator_out7933_out1 <= Logical_Operator_out1727_out1 XOR Logical_Operator_out1791_out1;

  Logical_Operator_out7934_out1 <= Logical_Operator_out1728_out1 XOR Logical_Operator_out1792_out1;

  Logical_Operator_out7935_out1 <= Logical_Operator_out704_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out7936_out1 <= in1408 XOR in1536;

  Logical_Operator_out7937_out1 <= Logical_Operator_out6913_out1 XOR Logical_Operator_out6977_out1;

  Logical_Operator_out7938_out1 <= Logical_Operator_out6914_out1 XOR Logical_Operator_out6978_out1;

  Logical_Operator_out7939_out1 <= Logical_Operator_out6915_out1 XOR Logical_Operator_out6979_out1;

  Logical_Operator_out7940_out1 <= Logical_Operator_out6916_out1 XOR Logical_Operator_out6980_out1;

  Logical_Operator_out7941_out1 <= Logical_Operator_out6917_out1 XOR Logical_Operator_out6981_out1;

  Logical_Operator_out7942_out1 <= Logical_Operator_out6918_out1 XOR Logical_Operator_out6982_out1;

  Logical_Operator_out7943_out1 <= Logical_Operator_out6919_out1 XOR Logical_Operator_out6983_out1;

  Logical_Operator_out7944_out1 <= Logical_Operator_out6920_out1 XOR Logical_Operator_out6984_out1;

  Logical_Operator_out7945_out1 <= Logical_Operator_out6921_out1 XOR Logical_Operator_out6985_out1;

  Logical_Operator_out7946_out1 <= Logical_Operator_out6922_out1 XOR Logical_Operator_out6986_out1;

  Logical_Operator_out7947_out1 <= Logical_Operator_out6923_out1 XOR Logical_Operator_out6987_out1;

  Logical_Operator_out7948_out1 <= Logical_Operator_out6924_out1 XOR Logical_Operator_out6988_out1;

  Logical_Operator_out7949_out1 <= Logical_Operator_out6925_out1 XOR Logical_Operator_out6989_out1;

  Logical_Operator_out7950_out1 <= Logical_Operator_out6926_out1 XOR Logical_Operator_out6990_out1;

  Logical_Operator_out7951_out1 <= Logical_Operator_out6927_out1 XOR Logical_Operator_out6991_out1;

  Logical_Operator_out7952_out1 <= Logical_Operator_out6928_out1 XOR Logical_Operator_out6992_out1;

  Logical_Operator_out7953_out1 <= Logical_Operator_out6929_out1 XOR Logical_Operator_out6993_out1;

  Logical_Operator_out7954_out1 <= Logical_Operator_out6930_out1 XOR Logical_Operator_out6994_out1;

  Logical_Operator_out7955_out1 <= Logical_Operator_out6931_out1 XOR Logical_Operator_out6995_out1;

  Logical_Operator_out7956_out1 <= Logical_Operator_out6932_out1 XOR Logical_Operator_out6996_out1;

  Logical_Operator_out7957_out1 <= Logical_Operator_out6933_out1 XOR Logical_Operator_out6997_out1;

  Logical_Operator_out7958_out1 <= Logical_Operator_out6934_out1 XOR Logical_Operator_out6998_out1;

  Logical_Operator_out7959_out1 <= Logical_Operator_out6935_out1 XOR Logical_Operator_out6999_out1;

  Logical_Operator_out7960_out1 <= Logical_Operator_out6936_out1 XOR Logical_Operator_out7000_out1;

  Logical_Operator_out7961_out1 <= Logical_Operator_out6937_out1 XOR Logical_Operator_out7001_out1;

  Logical_Operator_out7962_out1 <= Logical_Operator_out6938_out1 XOR Logical_Operator_out7002_out1;

  Logical_Operator_out7963_out1 <= Logical_Operator_out6939_out1 XOR Logical_Operator_out7003_out1;

  Logical_Operator_out7964_out1 <= Logical_Operator_out6940_out1 XOR Logical_Operator_out7004_out1;

  Logical_Operator_out7965_out1 <= Logical_Operator_out6941_out1 XOR Logical_Operator_out7005_out1;

  Logical_Operator_out7966_out1 <= Logical_Operator_out6942_out1 XOR Logical_Operator_out7006_out1;

  Logical_Operator_out7967_out1 <= Logical_Operator_out6943_out1 XOR Logical_Operator_out7007_out1;

  Logical_Operator_out7968_out1 <= Logical_Operator_out6944_out1 XOR Logical_Operator_out7008_out1;

  Logical_Operator_out7969_out1 <= Logical_Operator_out6945_out1 XOR Logical_Operator_out7009_out1;

  Logical_Operator_out7970_out1 <= Logical_Operator_out6946_out1 XOR Logical_Operator_out7010_out1;

  Logical_Operator_out7971_out1 <= Logical_Operator_out6947_out1 XOR Logical_Operator_out7011_out1;

  Logical_Operator_out7972_out1 <= Logical_Operator_out6948_out1 XOR Logical_Operator_out7012_out1;

  Logical_Operator_out7973_out1 <= Logical_Operator_out6949_out1 XOR Logical_Operator_out7013_out1;

  Logical_Operator_out7974_out1 <= Logical_Operator_out6950_out1 XOR Logical_Operator_out7014_out1;

  Logical_Operator_out7975_out1 <= Logical_Operator_out6951_out1 XOR Logical_Operator_out7015_out1;

  Logical_Operator_out7976_out1 <= Logical_Operator_out6952_out1 XOR Logical_Operator_out7016_out1;

  Logical_Operator_out7977_out1 <= Logical_Operator_out6953_out1 XOR Logical_Operator_out7017_out1;

  Logical_Operator_out7978_out1 <= Logical_Operator_out6954_out1 XOR Logical_Operator_out7018_out1;

  Logical_Operator_out7979_out1 <= Logical_Operator_out6955_out1 XOR Logical_Operator_out7019_out1;

  Logical_Operator_out7980_out1 <= Logical_Operator_out6956_out1 XOR Logical_Operator_out7020_out1;

  Logical_Operator_out7981_out1 <= Logical_Operator_out6957_out1 XOR Logical_Operator_out7021_out1;

  Logical_Operator_out7982_out1 <= Logical_Operator_out6958_out1 XOR Logical_Operator_out7022_out1;

  Logical_Operator_out7983_out1 <= Logical_Operator_out6959_out1 XOR Logical_Operator_out7023_out1;

  Logical_Operator_out7984_out1 <= Logical_Operator_out6960_out1 XOR Logical_Operator_out7024_out1;

  Logical_Operator_out7985_out1 <= Logical_Operator_out6961_out1 XOR Logical_Operator_out7025_out1;

  Logical_Operator_out7986_out1 <= Logical_Operator_out6962_out1 XOR Logical_Operator_out7026_out1;

  Logical_Operator_out7987_out1 <= Logical_Operator_out6963_out1 XOR Logical_Operator_out7027_out1;

  Logical_Operator_out7988_out1 <= Logical_Operator_out6964_out1 XOR Logical_Operator_out7028_out1;

  Logical_Operator_out7989_out1 <= Logical_Operator_out6965_out1 XOR Logical_Operator_out7029_out1;

  Logical_Operator_out7990_out1 <= Logical_Operator_out6966_out1 XOR Logical_Operator_out7030_out1;

  Logical_Operator_out7991_out1 <= Logical_Operator_out6967_out1 XOR Logical_Operator_out7031_out1;

  Logical_Operator_out7992_out1 <= Logical_Operator_out6968_out1 XOR Logical_Operator_out7032_out1;

  Logical_Operator_out7993_out1 <= Logical_Operator_out6969_out1 XOR Logical_Operator_out7033_out1;

  Logical_Operator_out7994_out1 <= Logical_Operator_out6970_out1 XOR Logical_Operator_out7034_out1;

  Logical_Operator_out7995_out1 <= Logical_Operator_out6971_out1 XOR Logical_Operator_out7035_out1;

  Logical_Operator_out7996_out1 <= Logical_Operator_out6972_out1 XOR Logical_Operator_out7036_out1;

  Logical_Operator_out7997_out1 <= Logical_Operator_out6973_out1 XOR Logical_Operator_out7037_out1;

  Logical_Operator_out7998_out1 <= Logical_Operator_out6974_out1 XOR Logical_Operator_out7038_out1;

  Logical_Operator_out7999_out1 <= Logical_Operator_out6975_out1 XOR Logical_Operator_out7039_out1;

  Logical_Operator_out8000_out1 <= Logical_Operator_out6976_out1 XOR Logical_Operator_out7040_out1;

  Logical_Operator_out8001_out1 <= Logical_Operator_out5921_out1 XOR Logical_Operator_out5985_out1;

  Logical_Operator_out8002_out1 <= Logical_Operator_out5922_out1 XOR Logical_Operator_out5986_out1;

  Logical_Operator_out8003_out1 <= Logical_Operator_out5923_out1 XOR Logical_Operator_out5987_out1;

  Logical_Operator_out8004_out1 <= Logical_Operator_out5924_out1 XOR Logical_Operator_out5988_out1;

  Logical_Operator_out8005_out1 <= Logical_Operator_out5925_out1 XOR Logical_Operator_out5989_out1;

  Logical_Operator_out8006_out1 <= Logical_Operator_out5926_out1 XOR Logical_Operator_out5990_out1;

  Logical_Operator_out8007_out1 <= Logical_Operator_out5927_out1 XOR Logical_Operator_out5991_out1;

  Logical_Operator_out8008_out1 <= Logical_Operator_out5928_out1 XOR Logical_Operator_out5992_out1;

  Logical_Operator_out8009_out1 <= Logical_Operator_out5929_out1 XOR Logical_Operator_out5993_out1;

  Logical_Operator_out8010_out1 <= Logical_Operator_out5930_out1 XOR Logical_Operator_out5994_out1;

  Logical_Operator_out8011_out1 <= Logical_Operator_out5931_out1 XOR Logical_Operator_out5995_out1;

  Logical_Operator_out8012_out1 <= Logical_Operator_out5932_out1 XOR Logical_Operator_out5996_out1;

  Logical_Operator_out8013_out1 <= Logical_Operator_out5933_out1 XOR Logical_Operator_out5997_out1;

  Logical_Operator_out8014_out1 <= Logical_Operator_out5934_out1 XOR Logical_Operator_out5998_out1;

  Logical_Operator_out8015_out1 <= Logical_Operator_out5935_out1 XOR Logical_Operator_out5999_out1;

  Logical_Operator_out8016_out1 <= Logical_Operator_out5936_out1 XOR Logical_Operator_out6000_out1;

  Logical_Operator_out8017_out1 <= Logical_Operator_out5937_out1 XOR Logical_Operator_out6001_out1;

  Logical_Operator_out8018_out1 <= Logical_Operator_out5938_out1 XOR Logical_Operator_out6002_out1;

  Logical_Operator_out8019_out1 <= Logical_Operator_out5939_out1 XOR Logical_Operator_out6003_out1;

  Logical_Operator_out8020_out1 <= Logical_Operator_out5940_out1 XOR Logical_Operator_out6004_out1;

  Logical_Operator_out8021_out1 <= Logical_Operator_out5941_out1 XOR Logical_Operator_out6005_out1;

  Logical_Operator_out8022_out1 <= Logical_Operator_out5942_out1 XOR Logical_Operator_out6006_out1;

  Logical_Operator_out8023_out1 <= Logical_Operator_out5943_out1 XOR Logical_Operator_out6007_out1;

  Logical_Operator_out8024_out1 <= Logical_Operator_out5944_out1 XOR Logical_Operator_out6008_out1;

  Logical_Operator_out8025_out1 <= Logical_Operator_out5945_out1 XOR Logical_Operator_out6009_out1;

  Logical_Operator_out8026_out1 <= Logical_Operator_out5946_out1 XOR Logical_Operator_out6010_out1;

  Logical_Operator_out8027_out1 <= Logical_Operator_out5947_out1 XOR Logical_Operator_out6011_out1;

  Logical_Operator_out8028_out1 <= Logical_Operator_out5948_out1 XOR Logical_Operator_out6012_out1;

  Logical_Operator_out8029_out1 <= Logical_Operator_out5949_out1 XOR Logical_Operator_out6013_out1;

  Logical_Operator_out8030_out1 <= Logical_Operator_out5950_out1 XOR Logical_Operator_out6014_out1;

  Logical_Operator_out8031_out1 <= Logical_Operator_out5951_out1 XOR Logical_Operator_out6015_out1;

  Logical_Operator_out8032_out1 <= Logical_Operator_out5952_out1 XOR Logical_Operator_out6016_out1;

  Logical_Operator_out8033_out1 <= Logical_Operator_out4913_out1 XOR Logical_Operator_out4977_out1;

  Logical_Operator_out8034_out1 <= Logical_Operator_out4914_out1 XOR Logical_Operator_out4978_out1;

  Logical_Operator_out8035_out1 <= Logical_Operator_out4915_out1 XOR Logical_Operator_out4979_out1;

  Logical_Operator_out8036_out1 <= Logical_Operator_out4916_out1 XOR Logical_Operator_out4980_out1;

  Logical_Operator_out8037_out1 <= Logical_Operator_out4917_out1 XOR Logical_Operator_out4981_out1;

  Logical_Operator_out8038_out1 <= Logical_Operator_out4918_out1 XOR Logical_Operator_out4982_out1;

  Logical_Operator_out8039_out1 <= Logical_Operator_out4919_out1 XOR Logical_Operator_out4983_out1;

  Logical_Operator_out8040_out1 <= Logical_Operator_out4920_out1 XOR Logical_Operator_out4984_out1;

  Logical_Operator_out8041_out1 <= Logical_Operator_out4921_out1 XOR Logical_Operator_out4985_out1;

  Logical_Operator_out8042_out1 <= Logical_Operator_out4922_out1 XOR Logical_Operator_out4986_out1;

  Logical_Operator_out8043_out1 <= Logical_Operator_out4923_out1 XOR Logical_Operator_out4987_out1;

  Logical_Operator_out8044_out1 <= Logical_Operator_out4924_out1 XOR Logical_Operator_out4988_out1;

  Logical_Operator_out8045_out1 <= Logical_Operator_out4925_out1 XOR Logical_Operator_out4989_out1;

  Logical_Operator_out8046_out1 <= Logical_Operator_out4926_out1 XOR Logical_Operator_out4990_out1;

  Logical_Operator_out8047_out1 <= Logical_Operator_out4927_out1 XOR Logical_Operator_out4991_out1;

  Logical_Operator_out8048_out1 <= Logical_Operator_out4928_out1 XOR Logical_Operator_out4992_out1;

  Logical_Operator_out8049_out1 <= Logical_Operator_out3897_out1 XOR Logical_Operator_out3961_out1;

  Logical_Operator_out8050_out1 <= Logical_Operator_out3898_out1 XOR Logical_Operator_out3962_out1;

  Logical_Operator_out8051_out1 <= Logical_Operator_out3899_out1 XOR Logical_Operator_out3963_out1;

  Logical_Operator_out8052_out1 <= Logical_Operator_out3900_out1 XOR Logical_Operator_out3964_out1;

  Logical_Operator_out8053_out1 <= Logical_Operator_out3901_out1 XOR Logical_Operator_out3965_out1;

  Logical_Operator_out8054_out1 <= Logical_Operator_out3902_out1 XOR Logical_Operator_out3966_out1;

  Logical_Operator_out8055_out1 <= Logical_Operator_out3903_out1 XOR Logical_Operator_out3967_out1;

  Logical_Operator_out8056_out1 <= Logical_Operator_out3904_out1 XOR Logical_Operator_out3968_out1;

  Logical_Operator_out8057_out1 <= Logical_Operator_out2877_out1 XOR Logical_Operator_out2941_out1;

  Logical_Operator_out8058_out1 <= Logical_Operator_out2878_out1 XOR Logical_Operator_out2942_out1;

  Logical_Operator_out8059_out1 <= Logical_Operator_out2879_out1 XOR Logical_Operator_out2943_out1;

  Logical_Operator_out8060_out1 <= Logical_Operator_out2880_out1 XOR Logical_Operator_out2944_out1;

  Logical_Operator_out8061_out1 <= Logical_Operator_out1855_out1 XOR Logical_Operator_out1919_out1;

  Logical_Operator_out8062_out1 <= Logical_Operator_out1856_out1 XOR Logical_Operator_out1920_out1;

  Logical_Operator_out8063_out1 <= Logical_Operator_out832_out1 XOR Logical_Operator_out896_out1;

  Logical_Operator_out8064_out1 <= in1664 XOR in1792;

  Logical_Operator_out8065_out1 <= Logical_Operator_out7041_out1 XOR Logical_Operator_out7105_out1;

  Logical_Operator_out8066_out1 <= Logical_Operator_out7042_out1 XOR Logical_Operator_out7106_out1;

  Logical_Operator_out8067_out1 <= Logical_Operator_out7043_out1 XOR Logical_Operator_out7107_out1;

  Logical_Operator_out8068_out1 <= Logical_Operator_out7044_out1 XOR Logical_Operator_out7108_out1;

  Logical_Operator_out8069_out1 <= Logical_Operator_out7045_out1 XOR Logical_Operator_out7109_out1;

  Logical_Operator_out8070_out1 <= Logical_Operator_out7046_out1 XOR Logical_Operator_out7110_out1;

  Logical_Operator_out8071_out1 <= Logical_Operator_out7047_out1 XOR Logical_Operator_out7111_out1;

  Logical_Operator_out8072_out1 <= Logical_Operator_out7048_out1 XOR Logical_Operator_out7112_out1;

  Logical_Operator_out8073_out1 <= Logical_Operator_out7049_out1 XOR Logical_Operator_out7113_out1;

  Logical_Operator_out8074_out1 <= Logical_Operator_out7050_out1 XOR Logical_Operator_out7114_out1;

  Logical_Operator_out8075_out1 <= Logical_Operator_out7051_out1 XOR Logical_Operator_out7115_out1;

  Logical_Operator_out8076_out1 <= Logical_Operator_out7052_out1 XOR Logical_Operator_out7116_out1;

  Logical_Operator_out8077_out1 <= Logical_Operator_out7053_out1 XOR Logical_Operator_out7117_out1;

  Logical_Operator_out8078_out1 <= Logical_Operator_out7054_out1 XOR Logical_Operator_out7118_out1;

  Logical_Operator_out8079_out1 <= Logical_Operator_out7055_out1 XOR Logical_Operator_out7119_out1;

  Logical_Operator_out8080_out1 <= Logical_Operator_out7056_out1 XOR Logical_Operator_out7120_out1;

  Logical_Operator_out8081_out1 <= Logical_Operator_out7057_out1 XOR Logical_Operator_out7121_out1;

  Logical_Operator_out8082_out1 <= Logical_Operator_out7058_out1 XOR Logical_Operator_out7122_out1;

  Logical_Operator_out8083_out1 <= Logical_Operator_out7059_out1 XOR Logical_Operator_out7123_out1;

  Logical_Operator_out8084_out1 <= Logical_Operator_out7060_out1 XOR Logical_Operator_out7124_out1;

  Logical_Operator_out8085_out1 <= Logical_Operator_out7061_out1 XOR Logical_Operator_out7125_out1;

  Logical_Operator_out8086_out1 <= Logical_Operator_out7062_out1 XOR Logical_Operator_out7126_out1;

  Logical_Operator_out8087_out1 <= Logical_Operator_out7063_out1 XOR Logical_Operator_out7127_out1;

  Logical_Operator_out8088_out1 <= Logical_Operator_out7064_out1 XOR Logical_Operator_out7128_out1;

  Logical_Operator_out8089_out1 <= Logical_Operator_out7065_out1 XOR Logical_Operator_out7129_out1;

  Logical_Operator_out8090_out1 <= Logical_Operator_out7066_out1 XOR Logical_Operator_out7130_out1;

  Logical_Operator_out8091_out1 <= Logical_Operator_out7067_out1 XOR Logical_Operator_out7131_out1;

  Logical_Operator_out8092_out1 <= Logical_Operator_out7068_out1 XOR Logical_Operator_out7132_out1;

  Logical_Operator_out8093_out1 <= Logical_Operator_out7069_out1 XOR Logical_Operator_out7133_out1;

  Logical_Operator_out8094_out1 <= Logical_Operator_out7070_out1 XOR Logical_Operator_out7134_out1;

  Logical_Operator_out8095_out1 <= Logical_Operator_out7071_out1 XOR Logical_Operator_out7135_out1;

  Logical_Operator_out8096_out1 <= Logical_Operator_out7072_out1 XOR Logical_Operator_out7136_out1;

  Logical_Operator_out8097_out1 <= Logical_Operator_out7073_out1 XOR Logical_Operator_out7137_out1;

  Logical_Operator_out8098_out1 <= Logical_Operator_out7074_out1 XOR Logical_Operator_out7138_out1;

  Logical_Operator_out8099_out1 <= Logical_Operator_out7075_out1 XOR Logical_Operator_out7139_out1;

  Logical_Operator_out8100_out1 <= Logical_Operator_out7076_out1 XOR Logical_Operator_out7140_out1;

  Logical_Operator_out8101_out1 <= Logical_Operator_out7077_out1 XOR Logical_Operator_out7141_out1;

  Logical_Operator_out8102_out1 <= Logical_Operator_out7078_out1 XOR Logical_Operator_out7142_out1;

  Logical_Operator_out8103_out1 <= Logical_Operator_out7079_out1 XOR Logical_Operator_out7143_out1;

  Logical_Operator_out8104_out1 <= Logical_Operator_out7080_out1 XOR Logical_Operator_out7144_out1;

  Logical_Operator_out8105_out1 <= Logical_Operator_out7081_out1 XOR Logical_Operator_out7145_out1;

  Logical_Operator_out8106_out1 <= Logical_Operator_out7082_out1 XOR Logical_Operator_out7146_out1;

  Logical_Operator_out8107_out1 <= Logical_Operator_out7083_out1 XOR Logical_Operator_out7147_out1;

  Logical_Operator_out8108_out1 <= Logical_Operator_out7084_out1 XOR Logical_Operator_out7148_out1;

  Logical_Operator_out8109_out1 <= Logical_Operator_out7085_out1 XOR Logical_Operator_out7149_out1;

  Logical_Operator_out8110_out1 <= Logical_Operator_out7086_out1 XOR Logical_Operator_out7150_out1;

  Logical_Operator_out8111_out1 <= Logical_Operator_out7087_out1 XOR Logical_Operator_out7151_out1;

  Logical_Operator_out8112_out1 <= Logical_Operator_out7088_out1 XOR Logical_Operator_out7152_out1;

  Logical_Operator_out8113_out1 <= Logical_Operator_out7089_out1 XOR Logical_Operator_out7153_out1;

  Logical_Operator_out8114_out1 <= Logical_Operator_out7090_out1 XOR Logical_Operator_out7154_out1;

  Logical_Operator_out8115_out1 <= Logical_Operator_out7091_out1 XOR Logical_Operator_out7155_out1;

  Logical_Operator_out8116_out1 <= Logical_Operator_out7092_out1 XOR Logical_Operator_out7156_out1;

  Logical_Operator_out8117_out1 <= Logical_Operator_out7093_out1 XOR Logical_Operator_out7157_out1;

  Logical_Operator_out8118_out1 <= Logical_Operator_out7094_out1 XOR Logical_Operator_out7158_out1;

  Logical_Operator_out8119_out1 <= Logical_Operator_out7095_out1 XOR Logical_Operator_out7159_out1;

  Logical_Operator_out8120_out1 <= Logical_Operator_out7096_out1 XOR Logical_Operator_out7160_out1;

  Logical_Operator_out8121_out1 <= Logical_Operator_out7097_out1 XOR Logical_Operator_out7161_out1;

  Logical_Operator_out8122_out1 <= Logical_Operator_out7098_out1 XOR Logical_Operator_out7162_out1;

  Logical_Operator_out8123_out1 <= Logical_Operator_out7099_out1 XOR Logical_Operator_out7163_out1;

  Logical_Operator_out8124_out1 <= Logical_Operator_out7100_out1 XOR Logical_Operator_out7164_out1;

  Logical_Operator_out8125_out1 <= Logical_Operator_out7101_out1 XOR Logical_Operator_out7165_out1;

  Logical_Operator_out8126_out1 <= Logical_Operator_out7102_out1 XOR Logical_Operator_out7166_out1;

  Logical_Operator_out8127_out1 <= Logical_Operator_out7103_out1 XOR Logical_Operator_out7167_out1;

  Logical_Operator_out8128_out1 <= Logical_Operator_out7104_out1 XOR Logical_Operator_out7168_out1;

  Logical_Operator_out8129_out1 <= Logical_Operator_out6049_out1 XOR Logical_Operator_out6113_out1;

  Logical_Operator_out8130_out1 <= Logical_Operator_out6050_out1 XOR Logical_Operator_out6114_out1;

  Logical_Operator_out8131_out1 <= Logical_Operator_out6051_out1 XOR Logical_Operator_out6115_out1;

  Logical_Operator_out8132_out1 <= Logical_Operator_out6052_out1 XOR Logical_Operator_out6116_out1;

  Logical_Operator_out8133_out1 <= Logical_Operator_out6053_out1 XOR Logical_Operator_out6117_out1;

  Logical_Operator_out8134_out1 <= Logical_Operator_out6054_out1 XOR Logical_Operator_out6118_out1;

  Logical_Operator_out8135_out1 <= Logical_Operator_out6055_out1 XOR Logical_Operator_out6119_out1;

  Logical_Operator_out8136_out1 <= Logical_Operator_out6056_out1 XOR Logical_Operator_out6120_out1;

  Logical_Operator_out8137_out1 <= Logical_Operator_out6057_out1 XOR Logical_Operator_out6121_out1;

  Logical_Operator_out8138_out1 <= Logical_Operator_out6058_out1 XOR Logical_Operator_out6122_out1;

  Logical_Operator_out8139_out1 <= Logical_Operator_out6059_out1 XOR Logical_Operator_out6123_out1;

  Logical_Operator_out8140_out1 <= Logical_Operator_out6060_out1 XOR Logical_Operator_out6124_out1;

  Logical_Operator_out8141_out1 <= Logical_Operator_out6061_out1 XOR Logical_Operator_out6125_out1;

  Logical_Operator_out8142_out1 <= Logical_Operator_out6062_out1 XOR Logical_Operator_out6126_out1;

  Logical_Operator_out8143_out1 <= Logical_Operator_out6063_out1 XOR Logical_Operator_out6127_out1;

  Logical_Operator_out8144_out1 <= Logical_Operator_out6064_out1 XOR Logical_Operator_out6128_out1;

  Logical_Operator_out8145_out1 <= Logical_Operator_out6065_out1 XOR Logical_Operator_out6129_out1;

  Logical_Operator_out8146_out1 <= Logical_Operator_out6066_out1 XOR Logical_Operator_out6130_out1;

  Logical_Operator_out8147_out1 <= Logical_Operator_out6067_out1 XOR Logical_Operator_out6131_out1;

  Logical_Operator_out8148_out1 <= Logical_Operator_out6068_out1 XOR Logical_Operator_out6132_out1;

  Logical_Operator_out8149_out1 <= Logical_Operator_out6069_out1 XOR Logical_Operator_out6133_out1;

  Logical_Operator_out8150_out1 <= Logical_Operator_out6070_out1 XOR Logical_Operator_out6134_out1;

  Logical_Operator_out8151_out1 <= Logical_Operator_out6071_out1 XOR Logical_Operator_out6135_out1;

  Logical_Operator_out8152_out1 <= Logical_Operator_out6072_out1 XOR Logical_Operator_out6136_out1;

  Logical_Operator_out8153_out1 <= Logical_Operator_out6073_out1 XOR Logical_Operator_out6137_out1;

  Logical_Operator_out8154_out1 <= Logical_Operator_out6074_out1 XOR Logical_Operator_out6138_out1;

  Logical_Operator_out8155_out1 <= Logical_Operator_out6075_out1 XOR Logical_Operator_out6139_out1;

  Logical_Operator_out8156_out1 <= Logical_Operator_out6076_out1 XOR Logical_Operator_out6140_out1;

  Logical_Operator_out8157_out1 <= Logical_Operator_out6077_out1 XOR Logical_Operator_out6141_out1;

  Logical_Operator_out8158_out1 <= Logical_Operator_out6078_out1 XOR Logical_Operator_out6142_out1;

  Logical_Operator_out8159_out1 <= Logical_Operator_out6079_out1 XOR Logical_Operator_out6143_out1;

  Logical_Operator_out8160_out1 <= Logical_Operator_out6080_out1 XOR Logical_Operator_out6144_out1;

  Logical_Operator_out8161_out1 <= Logical_Operator_out5041_out1 XOR Logical_Operator_out5105_out1;

  Logical_Operator_out8162_out1 <= Logical_Operator_out5042_out1 XOR Logical_Operator_out5106_out1;

  Logical_Operator_out8163_out1 <= Logical_Operator_out5043_out1 XOR Logical_Operator_out5107_out1;

  Logical_Operator_out8164_out1 <= Logical_Operator_out5044_out1 XOR Logical_Operator_out5108_out1;

  Logical_Operator_out8165_out1 <= Logical_Operator_out5045_out1 XOR Logical_Operator_out5109_out1;

  Logical_Operator_out8166_out1 <= Logical_Operator_out5046_out1 XOR Logical_Operator_out5110_out1;

  Logical_Operator_out8167_out1 <= Logical_Operator_out5047_out1 XOR Logical_Operator_out5111_out1;

  Logical_Operator_out8168_out1 <= Logical_Operator_out5048_out1 XOR Logical_Operator_out5112_out1;

  Logical_Operator_out8169_out1 <= Logical_Operator_out5049_out1 XOR Logical_Operator_out5113_out1;

  Logical_Operator_out8170_out1 <= Logical_Operator_out5050_out1 XOR Logical_Operator_out5114_out1;

  Logical_Operator_out8171_out1 <= Logical_Operator_out5051_out1 XOR Logical_Operator_out5115_out1;

  Logical_Operator_out8172_out1 <= Logical_Operator_out5052_out1 XOR Logical_Operator_out5116_out1;

  Logical_Operator_out8173_out1 <= Logical_Operator_out5053_out1 XOR Logical_Operator_out5117_out1;

  Logical_Operator_out8174_out1 <= Logical_Operator_out5054_out1 XOR Logical_Operator_out5118_out1;

  Logical_Operator_out8175_out1 <= Logical_Operator_out5055_out1 XOR Logical_Operator_out5119_out1;

  Logical_Operator_out8176_out1 <= Logical_Operator_out5056_out1 XOR Logical_Operator_out5120_out1;

  Logical_Operator_out8177_out1 <= Logical_Operator_out4025_out1 XOR Logical_Operator_out4089_out1;

  Logical_Operator_out8178_out1 <= Logical_Operator_out4026_out1 XOR Logical_Operator_out4090_out1;

  Logical_Operator_out8179_out1 <= Logical_Operator_out4027_out1 XOR Logical_Operator_out4091_out1;

  Logical_Operator_out8180_out1 <= Logical_Operator_out4028_out1 XOR Logical_Operator_out4092_out1;

  Logical_Operator_out8181_out1 <= Logical_Operator_out4029_out1 XOR Logical_Operator_out4093_out1;

  Logical_Operator_out8182_out1 <= Logical_Operator_out4030_out1 XOR Logical_Operator_out4094_out1;

  Logical_Operator_out8183_out1 <= Logical_Operator_out4031_out1 XOR Logical_Operator_out4095_out1;

  Logical_Operator_out8184_out1 <= Logical_Operator_out4032_out1 XOR Logical_Operator_out4096_out1;

  Logical_Operator_out8185_out1 <= Logical_Operator_out3005_out1 XOR Logical_Operator_out3069_out1;

  Logical_Operator_out8186_out1 <= Logical_Operator_out3006_out1 XOR Logical_Operator_out3070_out1;

  Logical_Operator_out8187_out1 <= Logical_Operator_out3007_out1 XOR Logical_Operator_out3071_out1;

  Logical_Operator_out8188_out1 <= Logical_Operator_out3008_out1 XOR Logical_Operator_out3072_out1;

  Logical_Operator_out8189_out1 <= Logical_Operator_out1983_out1 XOR Logical_Operator_out2047_out1;

  Logical_Operator_out8190_out1 <= Logical_Operator_out1984_out1 XOR Logical_Operator_out2048_out1;

  Logical_Operator_out8191_out1 <= Logical_Operator_out960_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out8192_out1 <= in1920 XOR in2048;

  Logical_Operator_out8193_out1 <= Logical_Operator_out7169_out1 XOR Logical_Operator_out7297_out1;

  Logical_Operator_out8194_out1 <= Logical_Operator_out7170_out1 XOR Logical_Operator_out7298_out1;

  Logical_Operator_out8195_out1 <= Logical_Operator_out7171_out1 XOR Logical_Operator_out7299_out1;

  Logical_Operator_out8196_out1 <= Logical_Operator_out7172_out1 XOR Logical_Operator_out7300_out1;

  Logical_Operator_out8197_out1 <= Logical_Operator_out7173_out1 XOR Logical_Operator_out7301_out1;

  Logical_Operator_out8198_out1 <= Logical_Operator_out7174_out1 XOR Logical_Operator_out7302_out1;

  Logical_Operator_out8199_out1 <= Logical_Operator_out7175_out1 XOR Logical_Operator_out7303_out1;

  Logical_Operator_out8200_out1 <= Logical_Operator_out7176_out1 XOR Logical_Operator_out7304_out1;

  Logical_Operator_out8201_out1 <= Logical_Operator_out7177_out1 XOR Logical_Operator_out7305_out1;

  Logical_Operator_out8202_out1 <= Logical_Operator_out7178_out1 XOR Logical_Operator_out7306_out1;

  Logical_Operator_out8203_out1 <= Logical_Operator_out7179_out1 XOR Logical_Operator_out7307_out1;

  Logical_Operator_out8204_out1 <= Logical_Operator_out7180_out1 XOR Logical_Operator_out7308_out1;

  Logical_Operator_out8205_out1 <= Logical_Operator_out7181_out1 XOR Logical_Operator_out7309_out1;

  Logical_Operator_out8206_out1 <= Logical_Operator_out7182_out1 XOR Logical_Operator_out7310_out1;

  Logical_Operator_out8207_out1 <= Logical_Operator_out7183_out1 XOR Logical_Operator_out7311_out1;

  Logical_Operator_out8208_out1 <= Logical_Operator_out7184_out1 XOR Logical_Operator_out7312_out1;

  Logical_Operator_out8209_out1 <= Logical_Operator_out7185_out1 XOR Logical_Operator_out7313_out1;

  Logical_Operator_out8210_out1 <= Logical_Operator_out7186_out1 XOR Logical_Operator_out7314_out1;

  Logical_Operator_out8211_out1 <= Logical_Operator_out7187_out1 XOR Logical_Operator_out7315_out1;

  Logical_Operator_out8212_out1 <= Logical_Operator_out7188_out1 XOR Logical_Operator_out7316_out1;

  Logical_Operator_out8213_out1 <= Logical_Operator_out7189_out1 XOR Logical_Operator_out7317_out1;

  Logical_Operator_out8214_out1 <= Logical_Operator_out7190_out1 XOR Logical_Operator_out7318_out1;

  Logical_Operator_out8215_out1 <= Logical_Operator_out7191_out1 XOR Logical_Operator_out7319_out1;

  Logical_Operator_out8216_out1 <= Logical_Operator_out7192_out1 XOR Logical_Operator_out7320_out1;

  Logical_Operator_out8217_out1 <= Logical_Operator_out7193_out1 XOR Logical_Operator_out7321_out1;

  Logical_Operator_out8218_out1 <= Logical_Operator_out7194_out1 XOR Logical_Operator_out7322_out1;

  Logical_Operator_out8219_out1 <= Logical_Operator_out7195_out1 XOR Logical_Operator_out7323_out1;

  Logical_Operator_out8220_out1 <= Logical_Operator_out7196_out1 XOR Logical_Operator_out7324_out1;

  Logical_Operator_out8221_out1 <= Logical_Operator_out7197_out1 XOR Logical_Operator_out7325_out1;

  Logical_Operator_out8222_out1 <= Logical_Operator_out7198_out1 XOR Logical_Operator_out7326_out1;

  Logical_Operator_out8223_out1 <= Logical_Operator_out7199_out1 XOR Logical_Operator_out7327_out1;

  Logical_Operator_out8224_out1 <= Logical_Operator_out7200_out1 XOR Logical_Operator_out7328_out1;

  Logical_Operator_out8225_out1 <= Logical_Operator_out7201_out1 XOR Logical_Operator_out7329_out1;

  Logical_Operator_out8226_out1 <= Logical_Operator_out7202_out1 XOR Logical_Operator_out7330_out1;

  Logical_Operator_out8227_out1 <= Logical_Operator_out7203_out1 XOR Logical_Operator_out7331_out1;

  Logical_Operator_out8228_out1 <= Logical_Operator_out7204_out1 XOR Logical_Operator_out7332_out1;

  Logical_Operator_out8229_out1 <= Logical_Operator_out7205_out1 XOR Logical_Operator_out7333_out1;

  Logical_Operator_out8230_out1 <= Logical_Operator_out7206_out1 XOR Logical_Operator_out7334_out1;

  Logical_Operator_out8231_out1 <= Logical_Operator_out7207_out1 XOR Logical_Operator_out7335_out1;

  Logical_Operator_out8232_out1 <= Logical_Operator_out7208_out1 XOR Logical_Operator_out7336_out1;

  Logical_Operator_out8233_out1 <= Logical_Operator_out7209_out1 XOR Logical_Operator_out7337_out1;

  Logical_Operator_out8234_out1 <= Logical_Operator_out7210_out1 XOR Logical_Operator_out7338_out1;

  Logical_Operator_out8235_out1 <= Logical_Operator_out7211_out1 XOR Logical_Operator_out7339_out1;

  Logical_Operator_out8236_out1 <= Logical_Operator_out7212_out1 XOR Logical_Operator_out7340_out1;

  Logical_Operator_out8237_out1 <= Logical_Operator_out7213_out1 XOR Logical_Operator_out7341_out1;

  Logical_Operator_out8238_out1 <= Logical_Operator_out7214_out1 XOR Logical_Operator_out7342_out1;

  Logical_Operator_out8239_out1 <= Logical_Operator_out7215_out1 XOR Logical_Operator_out7343_out1;

  Logical_Operator_out8240_out1 <= Logical_Operator_out7216_out1 XOR Logical_Operator_out7344_out1;

  Logical_Operator_out8241_out1 <= Logical_Operator_out7217_out1 XOR Logical_Operator_out7345_out1;

  Logical_Operator_out8242_out1 <= Logical_Operator_out7218_out1 XOR Logical_Operator_out7346_out1;

  Logical_Operator_out8243_out1 <= Logical_Operator_out7219_out1 XOR Logical_Operator_out7347_out1;

  Logical_Operator_out8244_out1 <= Logical_Operator_out7220_out1 XOR Logical_Operator_out7348_out1;

  Logical_Operator_out8245_out1 <= Logical_Operator_out7221_out1 XOR Logical_Operator_out7349_out1;

  Logical_Operator_out8246_out1 <= Logical_Operator_out7222_out1 XOR Logical_Operator_out7350_out1;

  Logical_Operator_out8247_out1 <= Logical_Operator_out7223_out1 XOR Logical_Operator_out7351_out1;

  Logical_Operator_out8248_out1 <= Logical_Operator_out7224_out1 XOR Logical_Operator_out7352_out1;

  Logical_Operator_out8249_out1 <= Logical_Operator_out7225_out1 XOR Logical_Operator_out7353_out1;

  Logical_Operator_out8250_out1 <= Logical_Operator_out7226_out1 XOR Logical_Operator_out7354_out1;

  Logical_Operator_out8251_out1 <= Logical_Operator_out7227_out1 XOR Logical_Operator_out7355_out1;

  Logical_Operator_out8252_out1 <= Logical_Operator_out7228_out1 XOR Logical_Operator_out7356_out1;

  Logical_Operator_out8253_out1 <= Logical_Operator_out7229_out1 XOR Logical_Operator_out7357_out1;

  Logical_Operator_out8254_out1 <= Logical_Operator_out7230_out1 XOR Logical_Operator_out7358_out1;

  Logical_Operator_out8255_out1 <= Logical_Operator_out7231_out1 XOR Logical_Operator_out7359_out1;

  Logical_Operator_out8256_out1 <= Logical_Operator_out7232_out1 XOR Logical_Operator_out7360_out1;

  Logical_Operator_out8257_out1 <= Logical_Operator_out7233_out1 XOR Logical_Operator_out7361_out1;

  Logical_Operator_out8258_out1 <= Logical_Operator_out7234_out1 XOR Logical_Operator_out7362_out1;

  Logical_Operator_out8259_out1 <= Logical_Operator_out7235_out1 XOR Logical_Operator_out7363_out1;

  Logical_Operator_out8260_out1 <= Logical_Operator_out7236_out1 XOR Logical_Operator_out7364_out1;

  Logical_Operator_out8261_out1 <= Logical_Operator_out7237_out1 XOR Logical_Operator_out7365_out1;

  Logical_Operator_out8262_out1 <= Logical_Operator_out7238_out1 XOR Logical_Operator_out7366_out1;

  Logical_Operator_out8263_out1 <= Logical_Operator_out7239_out1 XOR Logical_Operator_out7367_out1;

  Logical_Operator_out8264_out1 <= Logical_Operator_out7240_out1 XOR Logical_Operator_out7368_out1;

  Logical_Operator_out8265_out1 <= Logical_Operator_out7241_out1 XOR Logical_Operator_out7369_out1;

  Logical_Operator_out8266_out1 <= Logical_Operator_out7242_out1 XOR Logical_Operator_out7370_out1;

  Logical_Operator_out8267_out1 <= Logical_Operator_out7243_out1 XOR Logical_Operator_out7371_out1;

  Logical_Operator_out8268_out1 <= Logical_Operator_out7244_out1 XOR Logical_Operator_out7372_out1;

  Logical_Operator_out8269_out1 <= Logical_Operator_out7245_out1 XOR Logical_Operator_out7373_out1;

  Logical_Operator_out8270_out1 <= Logical_Operator_out7246_out1 XOR Logical_Operator_out7374_out1;

  Logical_Operator_out8271_out1 <= Logical_Operator_out7247_out1 XOR Logical_Operator_out7375_out1;

  Logical_Operator_out8272_out1 <= Logical_Operator_out7248_out1 XOR Logical_Operator_out7376_out1;

  Logical_Operator_out8273_out1 <= Logical_Operator_out7249_out1 XOR Logical_Operator_out7377_out1;

  Logical_Operator_out8274_out1 <= Logical_Operator_out7250_out1 XOR Logical_Operator_out7378_out1;

  Logical_Operator_out8275_out1 <= Logical_Operator_out7251_out1 XOR Logical_Operator_out7379_out1;

  Logical_Operator_out8276_out1 <= Logical_Operator_out7252_out1 XOR Logical_Operator_out7380_out1;

  Logical_Operator_out8277_out1 <= Logical_Operator_out7253_out1 XOR Logical_Operator_out7381_out1;

  Logical_Operator_out8278_out1 <= Logical_Operator_out7254_out1 XOR Logical_Operator_out7382_out1;

  Logical_Operator_out8279_out1 <= Logical_Operator_out7255_out1 XOR Logical_Operator_out7383_out1;

  Logical_Operator_out8280_out1 <= Logical_Operator_out7256_out1 XOR Logical_Operator_out7384_out1;

  Logical_Operator_out8281_out1 <= Logical_Operator_out7257_out1 XOR Logical_Operator_out7385_out1;

  Logical_Operator_out8282_out1 <= Logical_Operator_out7258_out1 XOR Logical_Operator_out7386_out1;

  Logical_Operator_out8283_out1 <= Logical_Operator_out7259_out1 XOR Logical_Operator_out7387_out1;

  Logical_Operator_out8284_out1 <= Logical_Operator_out7260_out1 XOR Logical_Operator_out7388_out1;

  Logical_Operator_out8285_out1 <= Logical_Operator_out7261_out1 XOR Logical_Operator_out7389_out1;

  Logical_Operator_out8286_out1 <= Logical_Operator_out7262_out1 XOR Logical_Operator_out7390_out1;

  Logical_Operator_out8287_out1 <= Logical_Operator_out7263_out1 XOR Logical_Operator_out7391_out1;

  Logical_Operator_out8288_out1 <= Logical_Operator_out7264_out1 XOR Logical_Operator_out7392_out1;

  Logical_Operator_out8289_out1 <= Logical_Operator_out7265_out1 XOR Logical_Operator_out7393_out1;

  Logical_Operator_out8290_out1 <= Logical_Operator_out7266_out1 XOR Logical_Operator_out7394_out1;

  Logical_Operator_out8291_out1 <= Logical_Operator_out7267_out1 XOR Logical_Operator_out7395_out1;

  Logical_Operator_out8292_out1 <= Logical_Operator_out7268_out1 XOR Logical_Operator_out7396_out1;

  Logical_Operator_out8293_out1 <= Logical_Operator_out7269_out1 XOR Logical_Operator_out7397_out1;

  Logical_Operator_out8294_out1 <= Logical_Operator_out7270_out1 XOR Logical_Operator_out7398_out1;

  Logical_Operator_out8295_out1 <= Logical_Operator_out7271_out1 XOR Logical_Operator_out7399_out1;

  Logical_Operator_out8296_out1 <= Logical_Operator_out7272_out1 XOR Logical_Operator_out7400_out1;

  Logical_Operator_out8297_out1 <= Logical_Operator_out7273_out1 XOR Logical_Operator_out7401_out1;

  Logical_Operator_out8298_out1 <= Logical_Operator_out7274_out1 XOR Logical_Operator_out7402_out1;

  Logical_Operator_out8299_out1 <= Logical_Operator_out7275_out1 XOR Logical_Operator_out7403_out1;

  Logical_Operator_out8300_out1 <= Logical_Operator_out7276_out1 XOR Logical_Operator_out7404_out1;

  Logical_Operator_out8301_out1 <= Logical_Operator_out7277_out1 XOR Logical_Operator_out7405_out1;

  Logical_Operator_out8302_out1 <= Logical_Operator_out7278_out1 XOR Logical_Operator_out7406_out1;

  Logical_Operator_out8303_out1 <= Logical_Operator_out7279_out1 XOR Logical_Operator_out7407_out1;

  Logical_Operator_out8304_out1 <= Logical_Operator_out7280_out1 XOR Logical_Operator_out7408_out1;

  Logical_Operator_out8305_out1 <= Logical_Operator_out7281_out1 XOR Logical_Operator_out7409_out1;

  Logical_Operator_out8306_out1 <= Logical_Operator_out7282_out1 XOR Logical_Operator_out7410_out1;

  Logical_Operator_out8307_out1 <= Logical_Operator_out7283_out1 XOR Logical_Operator_out7411_out1;

  Logical_Operator_out8308_out1 <= Logical_Operator_out7284_out1 XOR Logical_Operator_out7412_out1;

  Logical_Operator_out8309_out1 <= Logical_Operator_out7285_out1 XOR Logical_Operator_out7413_out1;

  Logical_Operator_out8310_out1 <= Logical_Operator_out7286_out1 XOR Logical_Operator_out7414_out1;

  Logical_Operator_out8311_out1 <= Logical_Operator_out7287_out1 XOR Logical_Operator_out7415_out1;

  Logical_Operator_out8312_out1 <= Logical_Operator_out7288_out1 XOR Logical_Operator_out7416_out1;

  Logical_Operator_out8313_out1 <= Logical_Operator_out7289_out1 XOR Logical_Operator_out7417_out1;

  Logical_Operator_out8314_out1 <= Logical_Operator_out7290_out1 XOR Logical_Operator_out7418_out1;

  Logical_Operator_out8315_out1 <= Logical_Operator_out7291_out1 XOR Logical_Operator_out7419_out1;

  Logical_Operator_out8316_out1 <= Logical_Operator_out7292_out1 XOR Logical_Operator_out7420_out1;

  Logical_Operator_out8317_out1 <= Logical_Operator_out7293_out1 XOR Logical_Operator_out7421_out1;

  Logical_Operator_out8318_out1 <= Logical_Operator_out7294_out1 XOR Logical_Operator_out7422_out1;

  Logical_Operator_out8319_out1 <= Logical_Operator_out7295_out1 XOR Logical_Operator_out7423_out1;

  Logical_Operator_out8320_out1 <= Logical_Operator_out7296_out1 XOR Logical_Operator_out7424_out1;

  Logical_Operator_out8321_out1 <= Logical_Operator_out6209_out1 XOR Logical_Operator_out6337_out1;

  Logical_Operator_out8322_out1 <= Logical_Operator_out6210_out1 XOR Logical_Operator_out6338_out1;

  Logical_Operator_out8323_out1 <= Logical_Operator_out6211_out1 XOR Logical_Operator_out6339_out1;

  Logical_Operator_out8324_out1 <= Logical_Operator_out6212_out1 XOR Logical_Operator_out6340_out1;

  Logical_Operator_out8325_out1 <= Logical_Operator_out6213_out1 XOR Logical_Operator_out6341_out1;

  Logical_Operator_out8326_out1 <= Logical_Operator_out6214_out1 XOR Logical_Operator_out6342_out1;

  Logical_Operator_out8327_out1 <= Logical_Operator_out6215_out1 XOR Logical_Operator_out6343_out1;

  Logical_Operator_out8328_out1 <= Logical_Operator_out6216_out1 XOR Logical_Operator_out6344_out1;

  Logical_Operator_out8329_out1 <= Logical_Operator_out6217_out1 XOR Logical_Operator_out6345_out1;

  Logical_Operator_out8330_out1 <= Logical_Operator_out6218_out1 XOR Logical_Operator_out6346_out1;

  Logical_Operator_out8331_out1 <= Logical_Operator_out6219_out1 XOR Logical_Operator_out6347_out1;

  Logical_Operator_out8332_out1 <= Logical_Operator_out6220_out1 XOR Logical_Operator_out6348_out1;

  Logical_Operator_out8333_out1 <= Logical_Operator_out6221_out1 XOR Logical_Operator_out6349_out1;

  Logical_Operator_out8334_out1 <= Logical_Operator_out6222_out1 XOR Logical_Operator_out6350_out1;

  Logical_Operator_out8335_out1 <= Logical_Operator_out6223_out1 XOR Logical_Operator_out6351_out1;

  Logical_Operator_out8336_out1 <= Logical_Operator_out6224_out1 XOR Logical_Operator_out6352_out1;

  Logical_Operator_out8337_out1 <= Logical_Operator_out6225_out1 XOR Logical_Operator_out6353_out1;

  Logical_Operator_out8338_out1 <= Logical_Operator_out6226_out1 XOR Logical_Operator_out6354_out1;

  Logical_Operator_out8339_out1 <= Logical_Operator_out6227_out1 XOR Logical_Operator_out6355_out1;

  Logical_Operator_out8340_out1 <= Logical_Operator_out6228_out1 XOR Logical_Operator_out6356_out1;

  Logical_Operator_out8341_out1 <= Logical_Operator_out6229_out1 XOR Logical_Operator_out6357_out1;

  Logical_Operator_out8342_out1 <= Logical_Operator_out6230_out1 XOR Logical_Operator_out6358_out1;

  Logical_Operator_out8343_out1 <= Logical_Operator_out6231_out1 XOR Logical_Operator_out6359_out1;

  Logical_Operator_out8344_out1 <= Logical_Operator_out6232_out1 XOR Logical_Operator_out6360_out1;

  Logical_Operator_out8345_out1 <= Logical_Operator_out6233_out1 XOR Logical_Operator_out6361_out1;

  Logical_Operator_out8346_out1 <= Logical_Operator_out6234_out1 XOR Logical_Operator_out6362_out1;

  Logical_Operator_out8347_out1 <= Logical_Operator_out6235_out1 XOR Logical_Operator_out6363_out1;

  Logical_Operator_out8348_out1 <= Logical_Operator_out6236_out1 XOR Logical_Operator_out6364_out1;

  Logical_Operator_out8349_out1 <= Logical_Operator_out6237_out1 XOR Logical_Operator_out6365_out1;

  Logical_Operator_out8350_out1 <= Logical_Operator_out6238_out1 XOR Logical_Operator_out6366_out1;

  Logical_Operator_out8351_out1 <= Logical_Operator_out6239_out1 XOR Logical_Operator_out6367_out1;

  Logical_Operator_out8352_out1 <= Logical_Operator_out6240_out1 XOR Logical_Operator_out6368_out1;

  Logical_Operator_out8353_out1 <= Logical_Operator_out6241_out1 XOR Logical_Operator_out6369_out1;

  Logical_Operator_out8354_out1 <= Logical_Operator_out6242_out1 XOR Logical_Operator_out6370_out1;

  Logical_Operator_out8355_out1 <= Logical_Operator_out6243_out1 XOR Logical_Operator_out6371_out1;

  Logical_Operator_out8356_out1 <= Logical_Operator_out6244_out1 XOR Logical_Operator_out6372_out1;

  Logical_Operator_out8357_out1 <= Logical_Operator_out6245_out1 XOR Logical_Operator_out6373_out1;

  Logical_Operator_out8358_out1 <= Logical_Operator_out6246_out1 XOR Logical_Operator_out6374_out1;

  Logical_Operator_out8359_out1 <= Logical_Operator_out6247_out1 XOR Logical_Operator_out6375_out1;

  Logical_Operator_out8360_out1 <= Logical_Operator_out6248_out1 XOR Logical_Operator_out6376_out1;

  Logical_Operator_out8361_out1 <= Logical_Operator_out6249_out1 XOR Logical_Operator_out6377_out1;

  Logical_Operator_out8362_out1 <= Logical_Operator_out6250_out1 XOR Logical_Operator_out6378_out1;

  Logical_Operator_out8363_out1 <= Logical_Operator_out6251_out1 XOR Logical_Operator_out6379_out1;

  Logical_Operator_out8364_out1 <= Logical_Operator_out6252_out1 XOR Logical_Operator_out6380_out1;

  Logical_Operator_out8365_out1 <= Logical_Operator_out6253_out1 XOR Logical_Operator_out6381_out1;

  Logical_Operator_out8366_out1 <= Logical_Operator_out6254_out1 XOR Logical_Operator_out6382_out1;

  Logical_Operator_out8367_out1 <= Logical_Operator_out6255_out1 XOR Logical_Operator_out6383_out1;

  Logical_Operator_out8368_out1 <= Logical_Operator_out6256_out1 XOR Logical_Operator_out6384_out1;

  Logical_Operator_out8369_out1 <= Logical_Operator_out6257_out1 XOR Logical_Operator_out6385_out1;

  Logical_Operator_out8370_out1 <= Logical_Operator_out6258_out1 XOR Logical_Operator_out6386_out1;

  Logical_Operator_out8371_out1 <= Logical_Operator_out6259_out1 XOR Logical_Operator_out6387_out1;

  Logical_Operator_out8372_out1 <= Logical_Operator_out6260_out1 XOR Logical_Operator_out6388_out1;

  Logical_Operator_out8373_out1 <= Logical_Operator_out6261_out1 XOR Logical_Operator_out6389_out1;

  Logical_Operator_out8374_out1 <= Logical_Operator_out6262_out1 XOR Logical_Operator_out6390_out1;

  Logical_Operator_out8375_out1 <= Logical_Operator_out6263_out1 XOR Logical_Operator_out6391_out1;

  Logical_Operator_out8376_out1 <= Logical_Operator_out6264_out1 XOR Logical_Operator_out6392_out1;

  Logical_Operator_out8377_out1 <= Logical_Operator_out6265_out1 XOR Logical_Operator_out6393_out1;

  Logical_Operator_out8378_out1 <= Logical_Operator_out6266_out1 XOR Logical_Operator_out6394_out1;

  Logical_Operator_out8379_out1 <= Logical_Operator_out6267_out1 XOR Logical_Operator_out6395_out1;

  Logical_Operator_out8380_out1 <= Logical_Operator_out6268_out1 XOR Logical_Operator_out6396_out1;

  Logical_Operator_out8381_out1 <= Logical_Operator_out6269_out1 XOR Logical_Operator_out6397_out1;

  Logical_Operator_out8382_out1 <= Logical_Operator_out6270_out1 XOR Logical_Operator_out6398_out1;

  Logical_Operator_out8383_out1 <= Logical_Operator_out6271_out1 XOR Logical_Operator_out6399_out1;

  Logical_Operator_out8384_out1 <= Logical_Operator_out6272_out1 XOR Logical_Operator_out6400_out1;

  Logical_Operator_out8385_out1 <= Logical_Operator_out5217_out1 XOR Logical_Operator_out5345_out1;

  Logical_Operator_out8386_out1 <= Logical_Operator_out5218_out1 XOR Logical_Operator_out5346_out1;

  Logical_Operator_out8387_out1 <= Logical_Operator_out5219_out1 XOR Logical_Operator_out5347_out1;

  Logical_Operator_out8388_out1 <= Logical_Operator_out5220_out1 XOR Logical_Operator_out5348_out1;

  Logical_Operator_out8389_out1 <= Logical_Operator_out5221_out1 XOR Logical_Operator_out5349_out1;

  Logical_Operator_out8390_out1 <= Logical_Operator_out5222_out1 XOR Logical_Operator_out5350_out1;

  Logical_Operator_out8391_out1 <= Logical_Operator_out5223_out1 XOR Logical_Operator_out5351_out1;

  Logical_Operator_out8392_out1 <= Logical_Operator_out5224_out1 XOR Logical_Operator_out5352_out1;

  Logical_Operator_out8393_out1 <= Logical_Operator_out5225_out1 XOR Logical_Operator_out5353_out1;

  Logical_Operator_out8394_out1 <= Logical_Operator_out5226_out1 XOR Logical_Operator_out5354_out1;

  Logical_Operator_out8395_out1 <= Logical_Operator_out5227_out1 XOR Logical_Operator_out5355_out1;

  Logical_Operator_out8396_out1 <= Logical_Operator_out5228_out1 XOR Logical_Operator_out5356_out1;

  Logical_Operator_out8397_out1 <= Logical_Operator_out5229_out1 XOR Logical_Operator_out5357_out1;

  Logical_Operator_out8398_out1 <= Logical_Operator_out5230_out1 XOR Logical_Operator_out5358_out1;

  Logical_Operator_out8399_out1 <= Logical_Operator_out5231_out1 XOR Logical_Operator_out5359_out1;

  Logical_Operator_out8400_out1 <= Logical_Operator_out5232_out1 XOR Logical_Operator_out5360_out1;

  Logical_Operator_out8401_out1 <= Logical_Operator_out5233_out1 XOR Logical_Operator_out5361_out1;

  Logical_Operator_out8402_out1 <= Logical_Operator_out5234_out1 XOR Logical_Operator_out5362_out1;

  Logical_Operator_out8403_out1 <= Logical_Operator_out5235_out1 XOR Logical_Operator_out5363_out1;

  Logical_Operator_out8404_out1 <= Logical_Operator_out5236_out1 XOR Logical_Operator_out5364_out1;

  Logical_Operator_out8405_out1 <= Logical_Operator_out5237_out1 XOR Logical_Operator_out5365_out1;

  Logical_Operator_out8406_out1 <= Logical_Operator_out5238_out1 XOR Logical_Operator_out5366_out1;

  Logical_Operator_out8407_out1 <= Logical_Operator_out5239_out1 XOR Logical_Operator_out5367_out1;

  Logical_Operator_out8408_out1 <= Logical_Operator_out5240_out1 XOR Logical_Operator_out5368_out1;

  Logical_Operator_out8409_out1 <= Logical_Operator_out5241_out1 XOR Logical_Operator_out5369_out1;

  Logical_Operator_out8410_out1 <= Logical_Operator_out5242_out1 XOR Logical_Operator_out5370_out1;

  Logical_Operator_out8411_out1 <= Logical_Operator_out5243_out1 XOR Logical_Operator_out5371_out1;

  Logical_Operator_out8412_out1 <= Logical_Operator_out5244_out1 XOR Logical_Operator_out5372_out1;

  Logical_Operator_out8413_out1 <= Logical_Operator_out5245_out1 XOR Logical_Operator_out5373_out1;

  Logical_Operator_out8414_out1 <= Logical_Operator_out5246_out1 XOR Logical_Operator_out5374_out1;

  Logical_Operator_out8415_out1 <= Logical_Operator_out5247_out1 XOR Logical_Operator_out5375_out1;

  Logical_Operator_out8416_out1 <= Logical_Operator_out5248_out1 XOR Logical_Operator_out5376_out1;

  Logical_Operator_out8417_out1 <= Logical_Operator_out4209_out1 XOR Logical_Operator_out4337_out1;

  Logical_Operator_out8418_out1 <= Logical_Operator_out4210_out1 XOR Logical_Operator_out4338_out1;

  Logical_Operator_out8419_out1 <= Logical_Operator_out4211_out1 XOR Logical_Operator_out4339_out1;

  Logical_Operator_out8420_out1 <= Logical_Operator_out4212_out1 XOR Logical_Operator_out4340_out1;

  Logical_Operator_out8421_out1 <= Logical_Operator_out4213_out1 XOR Logical_Operator_out4341_out1;

  Logical_Operator_out8422_out1 <= Logical_Operator_out4214_out1 XOR Logical_Operator_out4342_out1;

  Logical_Operator_out8423_out1 <= Logical_Operator_out4215_out1 XOR Logical_Operator_out4343_out1;

  Logical_Operator_out8424_out1 <= Logical_Operator_out4216_out1 XOR Logical_Operator_out4344_out1;

  Logical_Operator_out8425_out1 <= Logical_Operator_out4217_out1 XOR Logical_Operator_out4345_out1;

  Logical_Operator_out8426_out1 <= Logical_Operator_out4218_out1 XOR Logical_Operator_out4346_out1;

  Logical_Operator_out8427_out1 <= Logical_Operator_out4219_out1 XOR Logical_Operator_out4347_out1;

  Logical_Operator_out8428_out1 <= Logical_Operator_out4220_out1 XOR Logical_Operator_out4348_out1;

  Logical_Operator_out8429_out1 <= Logical_Operator_out4221_out1 XOR Logical_Operator_out4349_out1;

  Logical_Operator_out8430_out1 <= Logical_Operator_out4222_out1 XOR Logical_Operator_out4350_out1;

  Logical_Operator_out8431_out1 <= Logical_Operator_out4223_out1 XOR Logical_Operator_out4351_out1;

  Logical_Operator_out8432_out1 <= Logical_Operator_out4224_out1 XOR Logical_Operator_out4352_out1;

  Logical_Operator_out8433_out1 <= Logical_Operator_out3193_out1 XOR Logical_Operator_out3321_out1;

  Logical_Operator_out8434_out1 <= Logical_Operator_out3194_out1 XOR Logical_Operator_out3322_out1;

  Logical_Operator_out8435_out1 <= Logical_Operator_out3195_out1 XOR Logical_Operator_out3323_out1;

  Logical_Operator_out8436_out1 <= Logical_Operator_out3196_out1 XOR Logical_Operator_out3324_out1;

  Logical_Operator_out8437_out1 <= Logical_Operator_out3197_out1 XOR Logical_Operator_out3325_out1;

  Logical_Operator_out8438_out1 <= Logical_Operator_out3198_out1 XOR Logical_Operator_out3326_out1;

  Logical_Operator_out8439_out1 <= Logical_Operator_out3199_out1 XOR Logical_Operator_out3327_out1;

  Logical_Operator_out8440_out1 <= Logical_Operator_out3200_out1 XOR Logical_Operator_out3328_out1;

  Logical_Operator_out8441_out1 <= Logical_Operator_out2173_out1 XOR Logical_Operator_out2301_out1;

  Logical_Operator_out8442_out1 <= Logical_Operator_out2174_out1 XOR Logical_Operator_out2302_out1;

  Logical_Operator_out8443_out1 <= Logical_Operator_out2175_out1 XOR Logical_Operator_out2303_out1;

  Logical_Operator_out8444_out1 <= Logical_Operator_out2176_out1 XOR Logical_Operator_out2304_out1;

  Logical_Operator_out8445_out1 <= Logical_Operator_out1151_out1 XOR Logical_Operator_out1279_out1;

  Logical_Operator_out8446_out1 <= Logical_Operator_out1152_out1 XOR Logical_Operator_out1280_out1;

  Logical_Operator_out8447_out1 <= Logical_Operator_out128_out1 XOR Logical_Operator_out256_out1;

  Logical_Operator_out8448_out1 <= in256 XOR in512;

  Logical_Operator_out8449_out1 <= Logical_Operator_out7425_out1 XOR Logical_Operator_out7553_out1;

  Logical_Operator_out8450_out1 <= Logical_Operator_out7426_out1 XOR Logical_Operator_out7554_out1;

  Logical_Operator_out8451_out1 <= Logical_Operator_out7427_out1 XOR Logical_Operator_out7555_out1;

  Logical_Operator_out8452_out1 <= Logical_Operator_out7428_out1 XOR Logical_Operator_out7556_out1;

  Logical_Operator_out8453_out1 <= Logical_Operator_out7429_out1 XOR Logical_Operator_out7557_out1;

  Logical_Operator_out8454_out1 <= Logical_Operator_out7430_out1 XOR Logical_Operator_out7558_out1;

  Logical_Operator_out8455_out1 <= Logical_Operator_out7431_out1 XOR Logical_Operator_out7559_out1;

  Logical_Operator_out8456_out1 <= Logical_Operator_out7432_out1 XOR Logical_Operator_out7560_out1;

  Logical_Operator_out8457_out1 <= Logical_Operator_out7433_out1 XOR Logical_Operator_out7561_out1;

  Logical_Operator_out8458_out1 <= Logical_Operator_out7434_out1 XOR Logical_Operator_out7562_out1;

  Logical_Operator_out8459_out1 <= Logical_Operator_out7435_out1 XOR Logical_Operator_out7563_out1;

  Logical_Operator_out8460_out1 <= Logical_Operator_out7436_out1 XOR Logical_Operator_out7564_out1;

  Logical_Operator_out8461_out1 <= Logical_Operator_out7437_out1 XOR Logical_Operator_out7565_out1;

  Logical_Operator_out8462_out1 <= Logical_Operator_out7438_out1 XOR Logical_Operator_out7566_out1;

  Logical_Operator_out8463_out1 <= Logical_Operator_out7439_out1 XOR Logical_Operator_out7567_out1;

  Logical_Operator_out8464_out1 <= Logical_Operator_out7440_out1 XOR Logical_Operator_out7568_out1;

  Logical_Operator_out8465_out1 <= Logical_Operator_out7441_out1 XOR Logical_Operator_out7569_out1;

  Logical_Operator_out8466_out1 <= Logical_Operator_out7442_out1 XOR Logical_Operator_out7570_out1;

  Logical_Operator_out8467_out1 <= Logical_Operator_out7443_out1 XOR Logical_Operator_out7571_out1;

  Logical_Operator_out8468_out1 <= Logical_Operator_out7444_out1 XOR Logical_Operator_out7572_out1;

  Logical_Operator_out8469_out1 <= Logical_Operator_out7445_out1 XOR Logical_Operator_out7573_out1;

  Logical_Operator_out8470_out1 <= Logical_Operator_out7446_out1 XOR Logical_Operator_out7574_out1;

  Logical_Operator_out8471_out1 <= Logical_Operator_out7447_out1 XOR Logical_Operator_out7575_out1;

  Logical_Operator_out8472_out1 <= Logical_Operator_out7448_out1 XOR Logical_Operator_out7576_out1;

  Logical_Operator_out8473_out1 <= Logical_Operator_out7449_out1 XOR Logical_Operator_out7577_out1;

  Logical_Operator_out8474_out1 <= Logical_Operator_out7450_out1 XOR Logical_Operator_out7578_out1;

  Logical_Operator_out8475_out1 <= Logical_Operator_out7451_out1 XOR Logical_Operator_out7579_out1;

  Logical_Operator_out8476_out1 <= Logical_Operator_out7452_out1 XOR Logical_Operator_out7580_out1;

  Logical_Operator_out8477_out1 <= Logical_Operator_out7453_out1 XOR Logical_Operator_out7581_out1;

  Logical_Operator_out8478_out1 <= Logical_Operator_out7454_out1 XOR Logical_Operator_out7582_out1;

  Logical_Operator_out8479_out1 <= Logical_Operator_out7455_out1 XOR Logical_Operator_out7583_out1;

  Logical_Operator_out8480_out1 <= Logical_Operator_out7456_out1 XOR Logical_Operator_out7584_out1;

  Logical_Operator_out8481_out1 <= Logical_Operator_out7457_out1 XOR Logical_Operator_out7585_out1;

  Logical_Operator_out8482_out1 <= Logical_Operator_out7458_out1 XOR Logical_Operator_out7586_out1;

  Logical_Operator_out8483_out1 <= Logical_Operator_out7459_out1 XOR Logical_Operator_out7587_out1;

  Logical_Operator_out8484_out1 <= Logical_Operator_out7460_out1 XOR Logical_Operator_out7588_out1;

  Logical_Operator_out8485_out1 <= Logical_Operator_out7461_out1 XOR Logical_Operator_out7589_out1;

  Logical_Operator_out8486_out1 <= Logical_Operator_out7462_out1 XOR Logical_Operator_out7590_out1;

  Logical_Operator_out8487_out1 <= Logical_Operator_out7463_out1 XOR Logical_Operator_out7591_out1;

  Logical_Operator_out8488_out1 <= Logical_Operator_out7464_out1 XOR Logical_Operator_out7592_out1;

  Logical_Operator_out8489_out1 <= Logical_Operator_out7465_out1 XOR Logical_Operator_out7593_out1;

  Logical_Operator_out8490_out1 <= Logical_Operator_out7466_out1 XOR Logical_Operator_out7594_out1;

  Logical_Operator_out8491_out1 <= Logical_Operator_out7467_out1 XOR Logical_Operator_out7595_out1;

  Logical_Operator_out8492_out1 <= Logical_Operator_out7468_out1 XOR Logical_Operator_out7596_out1;

  Logical_Operator_out8493_out1 <= Logical_Operator_out7469_out1 XOR Logical_Operator_out7597_out1;

  Logical_Operator_out8494_out1 <= Logical_Operator_out7470_out1 XOR Logical_Operator_out7598_out1;

  Logical_Operator_out8495_out1 <= Logical_Operator_out7471_out1 XOR Logical_Operator_out7599_out1;

  Logical_Operator_out8496_out1 <= Logical_Operator_out7472_out1 XOR Logical_Operator_out7600_out1;

  Logical_Operator_out8497_out1 <= Logical_Operator_out7473_out1 XOR Logical_Operator_out7601_out1;

  Logical_Operator_out8498_out1 <= Logical_Operator_out7474_out1 XOR Logical_Operator_out7602_out1;

  Logical_Operator_out8499_out1 <= Logical_Operator_out7475_out1 XOR Logical_Operator_out7603_out1;

  Logical_Operator_out8500_out1 <= Logical_Operator_out7476_out1 XOR Logical_Operator_out7604_out1;

  Logical_Operator_out8501_out1 <= Logical_Operator_out7477_out1 XOR Logical_Operator_out7605_out1;

  Logical_Operator_out8502_out1 <= Logical_Operator_out7478_out1 XOR Logical_Operator_out7606_out1;

  Logical_Operator_out8503_out1 <= Logical_Operator_out7479_out1 XOR Logical_Operator_out7607_out1;

  Logical_Operator_out8504_out1 <= Logical_Operator_out7480_out1 XOR Logical_Operator_out7608_out1;

  Logical_Operator_out8505_out1 <= Logical_Operator_out7481_out1 XOR Logical_Operator_out7609_out1;

  Logical_Operator_out8506_out1 <= Logical_Operator_out7482_out1 XOR Logical_Operator_out7610_out1;

  Logical_Operator_out8507_out1 <= Logical_Operator_out7483_out1 XOR Logical_Operator_out7611_out1;

  Logical_Operator_out8508_out1 <= Logical_Operator_out7484_out1 XOR Logical_Operator_out7612_out1;

  Logical_Operator_out8509_out1 <= Logical_Operator_out7485_out1 XOR Logical_Operator_out7613_out1;

  Logical_Operator_out8510_out1 <= Logical_Operator_out7486_out1 XOR Logical_Operator_out7614_out1;

  Logical_Operator_out8511_out1 <= Logical_Operator_out7487_out1 XOR Logical_Operator_out7615_out1;

  Logical_Operator_out8512_out1 <= Logical_Operator_out7488_out1 XOR Logical_Operator_out7616_out1;

  Logical_Operator_out8513_out1 <= Logical_Operator_out7489_out1 XOR Logical_Operator_out7617_out1;

  Logical_Operator_out8514_out1 <= Logical_Operator_out7490_out1 XOR Logical_Operator_out7618_out1;

  Logical_Operator_out8515_out1 <= Logical_Operator_out7491_out1 XOR Logical_Operator_out7619_out1;

  Logical_Operator_out8516_out1 <= Logical_Operator_out7492_out1 XOR Logical_Operator_out7620_out1;

  Logical_Operator_out8517_out1 <= Logical_Operator_out7493_out1 XOR Logical_Operator_out7621_out1;

  Logical_Operator_out8518_out1 <= Logical_Operator_out7494_out1 XOR Logical_Operator_out7622_out1;

  Logical_Operator_out8519_out1 <= Logical_Operator_out7495_out1 XOR Logical_Operator_out7623_out1;

  Logical_Operator_out8520_out1 <= Logical_Operator_out7496_out1 XOR Logical_Operator_out7624_out1;

  Logical_Operator_out8521_out1 <= Logical_Operator_out7497_out1 XOR Logical_Operator_out7625_out1;

  Logical_Operator_out8522_out1 <= Logical_Operator_out7498_out1 XOR Logical_Operator_out7626_out1;

  Logical_Operator_out8523_out1 <= Logical_Operator_out7499_out1 XOR Logical_Operator_out7627_out1;

  Logical_Operator_out8524_out1 <= Logical_Operator_out7500_out1 XOR Logical_Operator_out7628_out1;

  Logical_Operator_out8525_out1 <= Logical_Operator_out7501_out1 XOR Logical_Operator_out7629_out1;

  Logical_Operator_out8526_out1 <= Logical_Operator_out7502_out1 XOR Logical_Operator_out7630_out1;

  Logical_Operator_out8527_out1 <= Logical_Operator_out7503_out1 XOR Logical_Operator_out7631_out1;

  Logical_Operator_out8528_out1 <= Logical_Operator_out7504_out1 XOR Logical_Operator_out7632_out1;

  Logical_Operator_out8529_out1 <= Logical_Operator_out7505_out1 XOR Logical_Operator_out7633_out1;

  Logical_Operator_out8530_out1 <= Logical_Operator_out7506_out1 XOR Logical_Operator_out7634_out1;

  Logical_Operator_out8531_out1 <= Logical_Operator_out7507_out1 XOR Logical_Operator_out7635_out1;

  Logical_Operator_out8532_out1 <= Logical_Operator_out7508_out1 XOR Logical_Operator_out7636_out1;

  Logical_Operator_out8533_out1 <= Logical_Operator_out7509_out1 XOR Logical_Operator_out7637_out1;

  Logical_Operator_out8534_out1 <= Logical_Operator_out7510_out1 XOR Logical_Operator_out7638_out1;

  Logical_Operator_out8535_out1 <= Logical_Operator_out7511_out1 XOR Logical_Operator_out7639_out1;

  Logical_Operator_out8536_out1 <= Logical_Operator_out7512_out1 XOR Logical_Operator_out7640_out1;

  Logical_Operator_out8537_out1 <= Logical_Operator_out7513_out1 XOR Logical_Operator_out7641_out1;

  Logical_Operator_out8538_out1 <= Logical_Operator_out7514_out1 XOR Logical_Operator_out7642_out1;

  Logical_Operator_out8539_out1 <= Logical_Operator_out7515_out1 XOR Logical_Operator_out7643_out1;

  Logical_Operator_out8540_out1 <= Logical_Operator_out7516_out1 XOR Logical_Operator_out7644_out1;

  Logical_Operator_out8541_out1 <= Logical_Operator_out7517_out1 XOR Logical_Operator_out7645_out1;

  Logical_Operator_out8542_out1 <= Logical_Operator_out7518_out1 XOR Logical_Operator_out7646_out1;

  Logical_Operator_out8543_out1 <= Logical_Operator_out7519_out1 XOR Logical_Operator_out7647_out1;

  Logical_Operator_out8544_out1 <= Logical_Operator_out7520_out1 XOR Logical_Operator_out7648_out1;

  Logical_Operator_out8545_out1 <= Logical_Operator_out7521_out1 XOR Logical_Operator_out7649_out1;

  Logical_Operator_out8546_out1 <= Logical_Operator_out7522_out1 XOR Logical_Operator_out7650_out1;

  Logical_Operator_out8547_out1 <= Logical_Operator_out7523_out1 XOR Logical_Operator_out7651_out1;

  Logical_Operator_out8548_out1 <= Logical_Operator_out7524_out1 XOR Logical_Operator_out7652_out1;

  Logical_Operator_out8549_out1 <= Logical_Operator_out7525_out1 XOR Logical_Operator_out7653_out1;

  Logical_Operator_out8550_out1 <= Logical_Operator_out7526_out1 XOR Logical_Operator_out7654_out1;

  Logical_Operator_out8551_out1 <= Logical_Operator_out7527_out1 XOR Logical_Operator_out7655_out1;

  Logical_Operator_out8552_out1 <= Logical_Operator_out7528_out1 XOR Logical_Operator_out7656_out1;

  Logical_Operator_out8553_out1 <= Logical_Operator_out7529_out1 XOR Logical_Operator_out7657_out1;

  Logical_Operator_out8554_out1 <= Logical_Operator_out7530_out1 XOR Logical_Operator_out7658_out1;

  Logical_Operator_out8555_out1 <= Logical_Operator_out7531_out1 XOR Logical_Operator_out7659_out1;

  Logical_Operator_out8556_out1 <= Logical_Operator_out7532_out1 XOR Logical_Operator_out7660_out1;

  Logical_Operator_out8557_out1 <= Logical_Operator_out7533_out1 XOR Logical_Operator_out7661_out1;

  Logical_Operator_out8558_out1 <= Logical_Operator_out7534_out1 XOR Logical_Operator_out7662_out1;

  Logical_Operator_out8559_out1 <= Logical_Operator_out7535_out1 XOR Logical_Operator_out7663_out1;

  Logical_Operator_out8560_out1 <= Logical_Operator_out7536_out1 XOR Logical_Operator_out7664_out1;

  Logical_Operator_out8561_out1 <= Logical_Operator_out7537_out1 XOR Logical_Operator_out7665_out1;

  Logical_Operator_out8562_out1 <= Logical_Operator_out7538_out1 XOR Logical_Operator_out7666_out1;

  Logical_Operator_out8563_out1 <= Logical_Operator_out7539_out1 XOR Logical_Operator_out7667_out1;

  Logical_Operator_out8564_out1 <= Logical_Operator_out7540_out1 XOR Logical_Operator_out7668_out1;

  Logical_Operator_out8565_out1 <= Logical_Operator_out7541_out1 XOR Logical_Operator_out7669_out1;

  Logical_Operator_out8566_out1 <= Logical_Operator_out7542_out1 XOR Logical_Operator_out7670_out1;

  Logical_Operator_out8567_out1 <= Logical_Operator_out7543_out1 XOR Logical_Operator_out7671_out1;

  Logical_Operator_out8568_out1 <= Logical_Operator_out7544_out1 XOR Logical_Operator_out7672_out1;

  Logical_Operator_out8569_out1 <= Logical_Operator_out7545_out1 XOR Logical_Operator_out7673_out1;

  Logical_Operator_out8570_out1 <= Logical_Operator_out7546_out1 XOR Logical_Operator_out7674_out1;

  Logical_Operator_out8571_out1 <= Logical_Operator_out7547_out1 XOR Logical_Operator_out7675_out1;

  Logical_Operator_out8572_out1 <= Logical_Operator_out7548_out1 XOR Logical_Operator_out7676_out1;

  Logical_Operator_out8573_out1 <= Logical_Operator_out7549_out1 XOR Logical_Operator_out7677_out1;

  Logical_Operator_out8574_out1 <= Logical_Operator_out7550_out1 XOR Logical_Operator_out7678_out1;

  Logical_Operator_out8575_out1 <= Logical_Operator_out7551_out1 XOR Logical_Operator_out7679_out1;

  Logical_Operator_out8576_out1 <= Logical_Operator_out7552_out1 XOR Logical_Operator_out7680_out1;

  Logical_Operator_out8577_out1 <= Logical_Operator_out6465_out1 XOR Logical_Operator_out6593_out1;

  Logical_Operator_out8578_out1 <= Logical_Operator_out6466_out1 XOR Logical_Operator_out6594_out1;

  Logical_Operator_out8579_out1 <= Logical_Operator_out6467_out1 XOR Logical_Operator_out6595_out1;

  Logical_Operator_out8580_out1 <= Logical_Operator_out6468_out1 XOR Logical_Operator_out6596_out1;

  Logical_Operator_out8581_out1 <= Logical_Operator_out6469_out1 XOR Logical_Operator_out6597_out1;

  Logical_Operator_out8582_out1 <= Logical_Operator_out6470_out1 XOR Logical_Operator_out6598_out1;

  Logical_Operator_out8583_out1 <= Logical_Operator_out6471_out1 XOR Logical_Operator_out6599_out1;

  Logical_Operator_out8584_out1 <= Logical_Operator_out6472_out1 XOR Logical_Operator_out6600_out1;

  Logical_Operator_out8585_out1 <= Logical_Operator_out6473_out1 XOR Logical_Operator_out6601_out1;

  Logical_Operator_out8586_out1 <= Logical_Operator_out6474_out1 XOR Logical_Operator_out6602_out1;

  Logical_Operator_out8587_out1 <= Logical_Operator_out6475_out1 XOR Logical_Operator_out6603_out1;

  Logical_Operator_out8588_out1 <= Logical_Operator_out6476_out1 XOR Logical_Operator_out6604_out1;

  Logical_Operator_out8589_out1 <= Logical_Operator_out6477_out1 XOR Logical_Operator_out6605_out1;

  Logical_Operator_out8590_out1 <= Logical_Operator_out6478_out1 XOR Logical_Operator_out6606_out1;

  Logical_Operator_out8591_out1 <= Logical_Operator_out6479_out1 XOR Logical_Operator_out6607_out1;

  Logical_Operator_out8592_out1 <= Logical_Operator_out6480_out1 XOR Logical_Operator_out6608_out1;

  Logical_Operator_out8593_out1 <= Logical_Operator_out6481_out1 XOR Logical_Operator_out6609_out1;

  Logical_Operator_out8594_out1 <= Logical_Operator_out6482_out1 XOR Logical_Operator_out6610_out1;

  Logical_Operator_out8595_out1 <= Logical_Operator_out6483_out1 XOR Logical_Operator_out6611_out1;

  Logical_Operator_out8596_out1 <= Logical_Operator_out6484_out1 XOR Logical_Operator_out6612_out1;

  Logical_Operator_out8597_out1 <= Logical_Operator_out6485_out1 XOR Logical_Operator_out6613_out1;

  Logical_Operator_out8598_out1 <= Logical_Operator_out6486_out1 XOR Logical_Operator_out6614_out1;

  Logical_Operator_out8599_out1 <= Logical_Operator_out6487_out1 XOR Logical_Operator_out6615_out1;

  Logical_Operator_out8600_out1 <= Logical_Operator_out6488_out1 XOR Logical_Operator_out6616_out1;

  Logical_Operator_out8601_out1 <= Logical_Operator_out6489_out1 XOR Logical_Operator_out6617_out1;

  Logical_Operator_out8602_out1 <= Logical_Operator_out6490_out1 XOR Logical_Operator_out6618_out1;

  Logical_Operator_out8603_out1 <= Logical_Operator_out6491_out1 XOR Logical_Operator_out6619_out1;

  Logical_Operator_out8604_out1 <= Logical_Operator_out6492_out1 XOR Logical_Operator_out6620_out1;

  Logical_Operator_out8605_out1 <= Logical_Operator_out6493_out1 XOR Logical_Operator_out6621_out1;

  Logical_Operator_out8606_out1 <= Logical_Operator_out6494_out1 XOR Logical_Operator_out6622_out1;

  Logical_Operator_out8607_out1 <= Logical_Operator_out6495_out1 XOR Logical_Operator_out6623_out1;

  Logical_Operator_out8608_out1 <= Logical_Operator_out6496_out1 XOR Logical_Operator_out6624_out1;

  Logical_Operator_out8609_out1 <= Logical_Operator_out6497_out1 XOR Logical_Operator_out6625_out1;

  Logical_Operator_out8610_out1 <= Logical_Operator_out6498_out1 XOR Logical_Operator_out6626_out1;

  Logical_Operator_out8611_out1 <= Logical_Operator_out6499_out1 XOR Logical_Operator_out6627_out1;

  Logical_Operator_out8612_out1 <= Logical_Operator_out6500_out1 XOR Logical_Operator_out6628_out1;

  Logical_Operator_out8613_out1 <= Logical_Operator_out6501_out1 XOR Logical_Operator_out6629_out1;

  Logical_Operator_out8614_out1 <= Logical_Operator_out6502_out1 XOR Logical_Operator_out6630_out1;

  Logical_Operator_out8615_out1 <= Logical_Operator_out6503_out1 XOR Logical_Operator_out6631_out1;

  Logical_Operator_out8616_out1 <= Logical_Operator_out6504_out1 XOR Logical_Operator_out6632_out1;

  Logical_Operator_out8617_out1 <= Logical_Operator_out6505_out1 XOR Logical_Operator_out6633_out1;

  Logical_Operator_out8618_out1 <= Logical_Operator_out6506_out1 XOR Logical_Operator_out6634_out1;

  Logical_Operator_out8619_out1 <= Logical_Operator_out6507_out1 XOR Logical_Operator_out6635_out1;

  Logical_Operator_out8620_out1 <= Logical_Operator_out6508_out1 XOR Logical_Operator_out6636_out1;

  Logical_Operator_out8621_out1 <= Logical_Operator_out6509_out1 XOR Logical_Operator_out6637_out1;

  Logical_Operator_out8622_out1 <= Logical_Operator_out6510_out1 XOR Logical_Operator_out6638_out1;

  Logical_Operator_out8623_out1 <= Logical_Operator_out6511_out1 XOR Logical_Operator_out6639_out1;

  Logical_Operator_out8624_out1 <= Logical_Operator_out6512_out1 XOR Logical_Operator_out6640_out1;

  Logical_Operator_out8625_out1 <= Logical_Operator_out6513_out1 XOR Logical_Operator_out6641_out1;

  Logical_Operator_out8626_out1 <= Logical_Operator_out6514_out1 XOR Logical_Operator_out6642_out1;

  Logical_Operator_out8627_out1 <= Logical_Operator_out6515_out1 XOR Logical_Operator_out6643_out1;

  Logical_Operator_out8628_out1 <= Logical_Operator_out6516_out1 XOR Logical_Operator_out6644_out1;

  Logical_Operator_out8629_out1 <= Logical_Operator_out6517_out1 XOR Logical_Operator_out6645_out1;

  Logical_Operator_out8630_out1 <= Logical_Operator_out6518_out1 XOR Logical_Operator_out6646_out1;

  Logical_Operator_out8631_out1 <= Logical_Operator_out6519_out1 XOR Logical_Operator_out6647_out1;

  Logical_Operator_out8632_out1 <= Logical_Operator_out6520_out1 XOR Logical_Operator_out6648_out1;

  Logical_Operator_out8633_out1 <= Logical_Operator_out6521_out1 XOR Logical_Operator_out6649_out1;

  Logical_Operator_out8634_out1 <= Logical_Operator_out6522_out1 XOR Logical_Operator_out6650_out1;

  Logical_Operator_out8635_out1 <= Logical_Operator_out6523_out1 XOR Logical_Operator_out6651_out1;

  Logical_Operator_out8636_out1 <= Logical_Operator_out6524_out1 XOR Logical_Operator_out6652_out1;

  Logical_Operator_out8637_out1 <= Logical_Operator_out6525_out1 XOR Logical_Operator_out6653_out1;

  Logical_Operator_out8638_out1 <= Logical_Operator_out6526_out1 XOR Logical_Operator_out6654_out1;

  Logical_Operator_out8639_out1 <= Logical_Operator_out6527_out1 XOR Logical_Operator_out6655_out1;

  Logical_Operator_out8640_out1 <= Logical_Operator_out6528_out1 XOR Logical_Operator_out6656_out1;

  Logical_Operator_out8641_out1 <= Logical_Operator_out5473_out1 XOR Logical_Operator_out5601_out1;

  Logical_Operator_out8642_out1 <= Logical_Operator_out5474_out1 XOR Logical_Operator_out5602_out1;

  Logical_Operator_out8643_out1 <= Logical_Operator_out5475_out1 XOR Logical_Operator_out5603_out1;

  Logical_Operator_out8644_out1 <= Logical_Operator_out5476_out1 XOR Logical_Operator_out5604_out1;

  Logical_Operator_out8645_out1 <= Logical_Operator_out5477_out1 XOR Logical_Operator_out5605_out1;

  Logical_Operator_out8646_out1 <= Logical_Operator_out5478_out1 XOR Logical_Operator_out5606_out1;

  Logical_Operator_out8647_out1 <= Logical_Operator_out5479_out1 XOR Logical_Operator_out5607_out1;

  Logical_Operator_out8648_out1 <= Logical_Operator_out5480_out1 XOR Logical_Operator_out5608_out1;

  Logical_Operator_out8649_out1 <= Logical_Operator_out5481_out1 XOR Logical_Operator_out5609_out1;

  Logical_Operator_out8650_out1 <= Logical_Operator_out5482_out1 XOR Logical_Operator_out5610_out1;

  Logical_Operator_out8651_out1 <= Logical_Operator_out5483_out1 XOR Logical_Operator_out5611_out1;

  Logical_Operator_out8652_out1 <= Logical_Operator_out5484_out1 XOR Logical_Operator_out5612_out1;

  Logical_Operator_out8653_out1 <= Logical_Operator_out5485_out1 XOR Logical_Operator_out5613_out1;

  Logical_Operator_out8654_out1 <= Logical_Operator_out5486_out1 XOR Logical_Operator_out5614_out1;

  Logical_Operator_out8655_out1 <= Logical_Operator_out5487_out1 XOR Logical_Operator_out5615_out1;

  Logical_Operator_out8656_out1 <= Logical_Operator_out5488_out1 XOR Logical_Operator_out5616_out1;

  Logical_Operator_out8657_out1 <= Logical_Operator_out5489_out1 XOR Logical_Operator_out5617_out1;

  Logical_Operator_out8658_out1 <= Logical_Operator_out5490_out1 XOR Logical_Operator_out5618_out1;

  Logical_Operator_out8659_out1 <= Logical_Operator_out5491_out1 XOR Logical_Operator_out5619_out1;

  Logical_Operator_out8660_out1 <= Logical_Operator_out5492_out1 XOR Logical_Operator_out5620_out1;

  Logical_Operator_out8661_out1 <= Logical_Operator_out5493_out1 XOR Logical_Operator_out5621_out1;

  Logical_Operator_out8662_out1 <= Logical_Operator_out5494_out1 XOR Logical_Operator_out5622_out1;

  Logical_Operator_out8663_out1 <= Logical_Operator_out5495_out1 XOR Logical_Operator_out5623_out1;

  Logical_Operator_out8664_out1 <= Logical_Operator_out5496_out1 XOR Logical_Operator_out5624_out1;

  Logical_Operator_out8665_out1 <= Logical_Operator_out5497_out1 XOR Logical_Operator_out5625_out1;

  Logical_Operator_out8666_out1 <= Logical_Operator_out5498_out1 XOR Logical_Operator_out5626_out1;

  Logical_Operator_out8667_out1 <= Logical_Operator_out5499_out1 XOR Logical_Operator_out5627_out1;

  Logical_Operator_out8668_out1 <= Logical_Operator_out5500_out1 XOR Logical_Operator_out5628_out1;

  Logical_Operator_out8669_out1 <= Logical_Operator_out5501_out1 XOR Logical_Operator_out5629_out1;

  Logical_Operator_out8670_out1 <= Logical_Operator_out5502_out1 XOR Logical_Operator_out5630_out1;

  Logical_Operator_out8671_out1 <= Logical_Operator_out5503_out1 XOR Logical_Operator_out5631_out1;

  Logical_Operator_out8672_out1 <= Logical_Operator_out5504_out1 XOR Logical_Operator_out5632_out1;

  Logical_Operator_out8673_out1 <= Logical_Operator_out4465_out1 XOR Logical_Operator_out4593_out1;

  Logical_Operator_out8674_out1 <= Logical_Operator_out4466_out1 XOR Logical_Operator_out4594_out1;

  Logical_Operator_out8675_out1 <= Logical_Operator_out4467_out1 XOR Logical_Operator_out4595_out1;

  Logical_Operator_out8676_out1 <= Logical_Operator_out4468_out1 XOR Logical_Operator_out4596_out1;

  Logical_Operator_out8677_out1 <= Logical_Operator_out4469_out1 XOR Logical_Operator_out4597_out1;

  Logical_Operator_out8678_out1 <= Logical_Operator_out4470_out1 XOR Logical_Operator_out4598_out1;

  Logical_Operator_out8679_out1 <= Logical_Operator_out4471_out1 XOR Logical_Operator_out4599_out1;

  Logical_Operator_out8680_out1 <= Logical_Operator_out4472_out1 XOR Logical_Operator_out4600_out1;

  Logical_Operator_out8681_out1 <= Logical_Operator_out4473_out1 XOR Logical_Operator_out4601_out1;

  Logical_Operator_out8682_out1 <= Logical_Operator_out4474_out1 XOR Logical_Operator_out4602_out1;

  Logical_Operator_out8683_out1 <= Logical_Operator_out4475_out1 XOR Logical_Operator_out4603_out1;

  Logical_Operator_out8684_out1 <= Logical_Operator_out4476_out1 XOR Logical_Operator_out4604_out1;

  Logical_Operator_out8685_out1 <= Logical_Operator_out4477_out1 XOR Logical_Operator_out4605_out1;

  Logical_Operator_out8686_out1 <= Logical_Operator_out4478_out1 XOR Logical_Operator_out4606_out1;

  Logical_Operator_out8687_out1 <= Logical_Operator_out4479_out1 XOR Logical_Operator_out4607_out1;

  Logical_Operator_out8688_out1 <= Logical_Operator_out4480_out1 XOR Logical_Operator_out4608_out1;

  Logical_Operator_out8689_out1 <= Logical_Operator_out3449_out1 XOR Logical_Operator_out3577_out1;

  Logical_Operator_out8690_out1 <= Logical_Operator_out3450_out1 XOR Logical_Operator_out3578_out1;

  Logical_Operator_out8691_out1 <= Logical_Operator_out3451_out1 XOR Logical_Operator_out3579_out1;

  Logical_Operator_out8692_out1 <= Logical_Operator_out3452_out1 XOR Logical_Operator_out3580_out1;

  Logical_Operator_out8693_out1 <= Logical_Operator_out3453_out1 XOR Logical_Operator_out3581_out1;

  Logical_Operator_out8694_out1 <= Logical_Operator_out3454_out1 XOR Logical_Operator_out3582_out1;

  Logical_Operator_out8695_out1 <= Logical_Operator_out3455_out1 XOR Logical_Operator_out3583_out1;

  Logical_Operator_out8696_out1 <= Logical_Operator_out3456_out1 XOR Logical_Operator_out3584_out1;

  Logical_Operator_out8697_out1 <= Logical_Operator_out2429_out1 XOR Logical_Operator_out2557_out1;

  Logical_Operator_out8698_out1 <= Logical_Operator_out2430_out1 XOR Logical_Operator_out2558_out1;

  Logical_Operator_out8699_out1 <= Logical_Operator_out2431_out1 XOR Logical_Operator_out2559_out1;

  Logical_Operator_out8700_out1 <= Logical_Operator_out2432_out1 XOR Logical_Operator_out2560_out1;

  Logical_Operator_out8701_out1 <= Logical_Operator_out1407_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out8702_out1 <= Logical_Operator_out1408_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out8703_out1 <= Logical_Operator_out384_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out8704_out1 <= in768 XOR in1024;

  Logical_Operator_out8705_out1 <= Logical_Operator_out7681_out1 XOR Logical_Operator_out7809_out1;

  Logical_Operator_out8706_out1 <= Logical_Operator_out7682_out1 XOR Logical_Operator_out7810_out1;

  Logical_Operator_out8707_out1 <= Logical_Operator_out7683_out1 XOR Logical_Operator_out7811_out1;

  Logical_Operator_out8708_out1 <= Logical_Operator_out7684_out1 XOR Logical_Operator_out7812_out1;

  Logical_Operator_out8709_out1 <= Logical_Operator_out7685_out1 XOR Logical_Operator_out7813_out1;

  Logical_Operator_out8710_out1 <= Logical_Operator_out7686_out1 XOR Logical_Operator_out7814_out1;

  Logical_Operator_out8711_out1 <= Logical_Operator_out7687_out1 XOR Logical_Operator_out7815_out1;

  Logical_Operator_out8712_out1 <= Logical_Operator_out7688_out1 XOR Logical_Operator_out7816_out1;

  Logical_Operator_out8713_out1 <= Logical_Operator_out7689_out1 XOR Logical_Operator_out7817_out1;

  Logical_Operator_out8714_out1 <= Logical_Operator_out7690_out1 XOR Logical_Operator_out7818_out1;

  Logical_Operator_out8715_out1 <= Logical_Operator_out7691_out1 XOR Logical_Operator_out7819_out1;

  Logical_Operator_out8716_out1 <= Logical_Operator_out7692_out1 XOR Logical_Operator_out7820_out1;

  Logical_Operator_out8717_out1 <= Logical_Operator_out7693_out1 XOR Logical_Operator_out7821_out1;

  Logical_Operator_out8718_out1 <= Logical_Operator_out7694_out1 XOR Logical_Operator_out7822_out1;

  Logical_Operator_out8719_out1 <= Logical_Operator_out7695_out1 XOR Logical_Operator_out7823_out1;

  Logical_Operator_out8720_out1 <= Logical_Operator_out7696_out1 XOR Logical_Operator_out7824_out1;

  Logical_Operator_out8721_out1 <= Logical_Operator_out7697_out1 XOR Logical_Operator_out7825_out1;

  Logical_Operator_out8722_out1 <= Logical_Operator_out7698_out1 XOR Logical_Operator_out7826_out1;

  Logical_Operator_out8723_out1 <= Logical_Operator_out7699_out1 XOR Logical_Operator_out7827_out1;

  Logical_Operator_out8724_out1 <= Logical_Operator_out7700_out1 XOR Logical_Operator_out7828_out1;

  Logical_Operator_out8725_out1 <= Logical_Operator_out7701_out1 XOR Logical_Operator_out7829_out1;

  Logical_Operator_out8726_out1 <= Logical_Operator_out7702_out1 XOR Logical_Operator_out7830_out1;

  Logical_Operator_out8727_out1 <= Logical_Operator_out7703_out1 XOR Logical_Operator_out7831_out1;

  Logical_Operator_out8728_out1 <= Logical_Operator_out7704_out1 XOR Logical_Operator_out7832_out1;

  Logical_Operator_out8729_out1 <= Logical_Operator_out7705_out1 XOR Logical_Operator_out7833_out1;

  Logical_Operator_out8730_out1 <= Logical_Operator_out7706_out1 XOR Logical_Operator_out7834_out1;

  Logical_Operator_out8731_out1 <= Logical_Operator_out7707_out1 XOR Logical_Operator_out7835_out1;

  Logical_Operator_out8732_out1 <= Logical_Operator_out7708_out1 XOR Logical_Operator_out7836_out1;

  Logical_Operator_out8733_out1 <= Logical_Operator_out7709_out1 XOR Logical_Operator_out7837_out1;

  Logical_Operator_out8734_out1 <= Logical_Operator_out7710_out1 XOR Logical_Operator_out7838_out1;

  Logical_Operator_out8735_out1 <= Logical_Operator_out7711_out1 XOR Logical_Operator_out7839_out1;

  Logical_Operator_out8736_out1 <= Logical_Operator_out7712_out1 XOR Logical_Operator_out7840_out1;

  Logical_Operator_out8737_out1 <= Logical_Operator_out7713_out1 XOR Logical_Operator_out7841_out1;

  Logical_Operator_out8738_out1 <= Logical_Operator_out7714_out1 XOR Logical_Operator_out7842_out1;

  Logical_Operator_out8739_out1 <= Logical_Operator_out7715_out1 XOR Logical_Operator_out7843_out1;

  Logical_Operator_out8740_out1 <= Logical_Operator_out7716_out1 XOR Logical_Operator_out7844_out1;

  Logical_Operator_out8741_out1 <= Logical_Operator_out7717_out1 XOR Logical_Operator_out7845_out1;

  Logical_Operator_out8742_out1 <= Logical_Operator_out7718_out1 XOR Logical_Operator_out7846_out1;

  Logical_Operator_out8743_out1 <= Logical_Operator_out7719_out1 XOR Logical_Operator_out7847_out1;

  Logical_Operator_out8744_out1 <= Logical_Operator_out7720_out1 XOR Logical_Operator_out7848_out1;

  Logical_Operator_out8745_out1 <= Logical_Operator_out7721_out1 XOR Logical_Operator_out7849_out1;

  Logical_Operator_out8746_out1 <= Logical_Operator_out7722_out1 XOR Logical_Operator_out7850_out1;

  Logical_Operator_out8747_out1 <= Logical_Operator_out7723_out1 XOR Logical_Operator_out7851_out1;

  Logical_Operator_out8748_out1 <= Logical_Operator_out7724_out1 XOR Logical_Operator_out7852_out1;

  Logical_Operator_out8749_out1 <= Logical_Operator_out7725_out1 XOR Logical_Operator_out7853_out1;

  Logical_Operator_out8750_out1 <= Logical_Operator_out7726_out1 XOR Logical_Operator_out7854_out1;

  Logical_Operator_out8751_out1 <= Logical_Operator_out7727_out1 XOR Logical_Operator_out7855_out1;

  Logical_Operator_out8752_out1 <= Logical_Operator_out7728_out1 XOR Logical_Operator_out7856_out1;

  Logical_Operator_out8753_out1 <= Logical_Operator_out7729_out1 XOR Logical_Operator_out7857_out1;

  Logical_Operator_out8754_out1 <= Logical_Operator_out7730_out1 XOR Logical_Operator_out7858_out1;

  Logical_Operator_out8755_out1 <= Logical_Operator_out7731_out1 XOR Logical_Operator_out7859_out1;

  Logical_Operator_out8756_out1 <= Logical_Operator_out7732_out1 XOR Logical_Operator_out7860_out1;

  Logical_Operator_out8757_out1 <= Logical_Operator_out7733_out1 XOR Logical_Operator_out7861_out1;

  Logical_Operator_out8758_out1 <= Logical_Operator_out7734_out1 XOR Logical_Operator_out7862_out1;

  Logical_Operator_out8759_out1 <= Logical_Operator_out7735_out1 XOR Logical_Operator_out7863_out1;

  Logical_Operator_out8760_out1 <= Logical_Operator_out7736_out1 XOR Logical_Operator_out7864_out1;

  Logical_Operator_out8761_out1 <= Logical_Operator_out7737_out1 XOR Logical_Operator_out7865_out1;

  Logical_Operator_out8762_out1 <= Logical_Operator_out7738_out1 XOR Logical_Operator_out7866_out1;

  Logical_Operator_out8763_out1 <= Logical_Operator_out7739_out1 XOR Logical_Operator_out7867_out1;

  Logical_Operator_out8764_out1 <= Logical_Operator_out7740_out1 XOR Logical_Operator_out7868_out1;

  Logical_Operator_out8765_out1 <= Logical_Operator_out7741_out1 XOR Logical_Operator_out7869_out1;

  Logical_Operator_out8766_out1 <= Logical_Operator_out7742_out1 XOR Logical_Operator_out7870_out1;

  Logical_Operator_out8767_out1 <= Logical_Operator_out7743_out1 XOR Logical_Operator_out7871_out1;

  Logical_Operator_out8768_out1 <= Logical_Operator_out7744_out1 XOR Logical_Operator_out7872_out1;

  Logical_Operator_out8769_out1 <= Logical_Operator_out7745_out1 XOR Logical_Operator_out7873_out1;

  Logical_Operator_out8770_out1 <= Logical_Operator_out7746_out1 XOR Logical_Operator_out7874_out1;

  Logical_Operator_out8771_out1 <= Logical_Operator_out7747_out1 XOR Logical_Operator_out7875_out1;

  Logical_Operator_out8772_out1 <= Logical_Operator_out7748_out1 XOR Logical_Operator_out7876_out1;

  Logical_Operator_out8773_out1 <= Logical_Operator_out7749_out1 XOR Logical_Operator_out7877_out1;

  Logical_Operator_out8774_out1 <= Logical_Operator_out7750_out1 XOR Logical_Operator_out7878_out1;

  Logical_Operator_out8775_out1 <= Logical_Operator_out7751_out1 XOR Logical_Operator_out7879_out1;

  Logical_Operator_out8776_out1 <= Logical_Operator_out7752_out1 XOR Logical_Operator_out7880_out1;

  Logical_Operator_out8777_out1 <= Logical_Operator_out7753_out1 XOR Logical_Operator_out7881_out1;

  Logical_Operator_out8778_out1 <= Logical_Operator_out7754_out1 XOR Logical_Operator_out7882_out1;

  Logical_Operator_out8779_out1 <= Logical_Operator_out7755_out1 XOR Logical_Operator_out7883_out1;

  Logical_Operator_out8780_out1 <= Logical_Operator_out7756_out1 XOR Logical_Operator_out7884_out1;

  Logical_Operator_out8781_out1 <= Logical_Operator_out7757_out1 XOR Logical_Operator_out7885_out1;

  Logical_Operator_out8782_out1 <= Logical_Operator_out7758_out1 XOR Logical_Operator_out7886_out1;

  Logical_Operator_out8783_out1 <= Logical_Operator_out7759_out1 XOR Logical_Operator_out7887_out1;

  Logical_Operator_out8784_out1 <= Logical_Operator_out7760_out1 XOR Logical_Operator_out7888_out1;

  Logical_Operator_out8785_out1 <= Logical_Operator_out7761_out1 XOR Logical_Operator_out7889_out1;

  Logical_Operator_out8786_out1 <= Logical_Operator_out7762_out1 XOR Logical_Operator_out7890_out1;

  Logical_Operator_out8787_out1 <= Logical_Operator_out7763_out1 XOR Logical_Operator_out7891_out1;

  Logical_Operator_out8788_out1 <= Logical_Operator_out7764_out1 XOR Logical_Operator_out7892_out1;

  Logical_Operator_out8789_out1 <= Logical_Operator_out7765_out1 XOR Logical_Operator_out7893_out1;

  Logical_Operator_out8790_out1 <= Logical_Operator_out7766_out1 XOR Logical_Operator_out7894_out1;

  Logical_Operator_out8791_out1 <= Logical_Operator_out7767_out1 XOR Logical_Operator_out7895_out1;

  Logical_Operator_out8792_out1 <= Logical_Operator_out7768_out1 XOR Logical_Operator_out7896_out1;

  Logical_Operator_out8793_out1 <= Logical_Operator_out7769_out1 XOR Logical_Operator_out7897_out1;

  Logical_Operator_out8794_out1 <= Logical_Operator_out7770_out1 XOR Logical_Operator_out7898_out1;

  Logical_Operator_out8795_out1 <= Logical_Operator_out7771_out1 XOR Logical_Operator_out7899_out1;

  Logical_Operator_out8796_out1 <= Logical_Operator_out7772_out1 XOR Logical_Operator_out7900_out1;

  Logical_Operator_out8797_out1 <= Logical_Operator_out7773_out1 XOR Logical_Operator_out7901_out1;

  Logical_Operator_out8798_out1 <= Logical_Operator_out7774_out1 XOR Logical_Operator_out7902_out1;

  Logical_Operator_out8799_out1 <= Logical_Operator_out7775_out1 XOR Logical_Operator_out7903_out1;

  Logical_Operator_out8800_out1 <= Logical_Operator_out7776_out1 XOR Logical_Operator_out7904_out1;

  Logical_Operator_out8801_out1 <= Logical_Operator_out7777_out1 XOR Logical_Operator_out7905_out1;

  Logical_Operator_out8802_out1 <= Logical_Operator_out7778_out1 XOR Logical_Operator_out7906_out1;

  Logical_Operator_out8803_out1 <= Logical_Operator_out7779_out1 XOR Logical_Operator_out7907_out1;

  Logical_Operator_out8804_out1 <= Logical_Operator_out7780_out1 XOR Logical_Operator_out7908_out1;

  Logical_Operator_out8805_out1 <= Logical_Operator_out7781_out1 XOR Logical_Operator_out7909_out1;

  Logical_Operator_out8806_out1 <= Logical_Operator_out7782_out1 XOR Logical_Operator_out7910_out1;

  Logical_Operator_out8807_out1 <= Logical_Operator_out7783_out1 XOR Logical_Operator_out7911_out1;

  Logical_Operator_out8808_out1 <= Logical_Operator_out7784_out1 XOR Logical_Operator_out7912_out1;

  Logical_Operator_out8809_out1 <= Logical_Operator_out7785_out1 XOR Logical_Operator_out7913_out1;

  Logical_Operator_out8810_out1 <= Logical_Operator_out7786_out1 XOR Logical_Operator_out7914_out1;

  Logical_Operator_out8811_out1 <= Logical_Operator_out7787_out1 XOR Logical_Operator_out7915_out1;

  Logical_Operator_out8812_out1 <= Logical_Operator_out7788_out1 XOR Logical_Operator_out7916_out1;

  Logical_Operator_out8813_out1 <= Logical_Operator_out7789_out1 XOR Logical_Operator_out7917_out1;

  Logical_Operator_out8814_out1 <= Logical_Operator_out7790_out1 XOR Logical_Operator_out7918_out1;

  Logical_Operator_out8815_out1 <= Logical_Operator_out7791_out1 XOR Logical_Operator_out7919_out1;

  Logical_Operator_out8816_out1 <= Logical_Operator_out7792_out1 XOR Logical_Operator_out7920_out1;

  Logical_Operator_out8817_out1 <= Logical_Operator_out7793_out1 XOR Logical_Operator_out7921_out1;

  Logical_Operator_out8818_out1 <= Logical_Operator_out7794_out1 XOR Logical_Operator_out7922_out1;

  Logical_Operator_out8819_out1 <= Logical_Operator_out7795_out1 XOR Logical_Operator_out7923_out1;

  Logical_Operator_out8820_out1 <= Logical_Operator_out7796_out1 XOR Logical_Operator_out7924_out1;

  Logical_Operator_out8821_out1 <= Logical_Operator_out7797_out1 XOR Logical_Operator_out7925_out1;

  Logical_Operator_out8822_out1 <= Logical_Operator_out7798_out1 XOR Logical_Operator_out7926_out1;

  Logical_Operator_out8823_out1 <= Logical_Operator_out7799_out1 XOR Logical_Operator_out7927_out1;

  Logical_Operator_out8824_out1 <= Logical_Operator_out7800_out1 XOR Logical_Operator_out7928_out1;

  Logical_Operator_out8825_out1 <= Logical_Operator_out7801_out1 XOR Logical_Operator_out7929_out1;

  Logical_Operator_out8826_out1 <= Logical_Operator_out7802_out1 XOR Logical_Operator_out7930_out1;

  Logical_Operator_out8827_out1 <= Logical_Operator_out7803_out1 XOR Logical_Operator_out7931_out1;

  Logical_Operator_out8828_out1 <= Logical_Operator_out7804_out1 XOR Logical_Operator_out7932_out1;

  Logical_Operator_out8829_out1 <= Logical_Operator_out7805_out1 XOR Logical_Operator_out7933_out1;

  Logical_Operator_out8830_out1 <= Logical_Operator_out7806_out1 XOR Logical_Operator_out7934_out1;

  Logical_Operator_out8831_out1 <= Logical_Operator_out7807_out1 XOR Logical_Operator_out7935_out1;

  Logical_Operator_out8832_out1 <= Logical_Operator_out7808_out1 XOR Logical_Operator_out7936_out1;

  Logical_Operator_out8833_out1 <= Logical_Operator_out6721_out1 XOR Logical_Operator_out6849_out1;

  Logical_Operator_out8834_out1 <= Logical_Operator_out6722_out1 XOR Logical_Operator_out6850_out1;

  Logical_Operator_out8835_out1 <= Logical_Operator_out6723_out1 XOR Logical_Operator_out6851_out1;

  Logical_Operator_out8836_out1 <= Logical_Operator_out6724_out1 XOR Logical_Operator_out6852_out1;

  Logical_Operator_out8837_out1 <= Logical_Operator_out6725_out1 XOR Logical_Operator_out6853_out1;

  Logical_Operator_out8838_out1 <= Logical_Operator_out6726_out1 XOR Logical_Operator_out6854_out1;

  Logical_Operator_out8839_out1 <= Logical_Operator_out6727_out1 XOR Logical_Operator_out6855_out1;

  Logical_Operator_out8840_out1 <= Logical_Operator_out6728_out1 XOR Logical_Operator_out6856_out1;

  Logical_Operator_out8841_out1 <= Logical_Operator_out6729_out1 XOR Logical_Operator_out6857_out1;

  Logical_Operator_out8842_out1 <= Logical_Operator_out6730_out1 XOR Logical_Operator_out6858_out1;

  Logical_Operator_out8843_out1 <= Logical_Operator_out6731_out1 XOR Logical_Operator_out6859_out1;

  Logical_Operator_out8844_out1 <= Logical_Operator_out6732_out1 XOR Logical_Operator_out6860_out1;

  Logical_Operator_out8845_out1 <= Logical_Operator_out6733_out1 XOR Logical_Operator_out6861_out1;

  Logical_Operator_out8846_out1 <= Logical_Operator_out6734_out1 XOR Logical_Operator_out6862_out1;

  Logical_Operator_out8847_out1 <= Logical_Operator_out6735_out1 XOR Logical_Operator_out6863_out1;

  Logical_Operator_out8848_out1 <= Logical_Operator_out6736_out1 XOR Logical_Operator_out6864_out1;

  Logical_Operator_out8849_out1 <= Logical_Operator_out6737_out1 XOR Logical_Operator_out6865_out1;

  Logical_Operator_out8850_out1 <= Logical_Operator_out6738_out1 XOR Logical_Operator_out6866_out1;

  Logical_Operator_out8851_out1 <= Logical_Operator_out6739_out1 XOR Logical_Operator_out6867_out1;

  Logical_Operator_out8852_out1 <= Logical_Operator_out6740_out1 XOR Logical_Operator_out6868_out1;

  Logical_Operator_out8853_out1 <= Logical_Operator_out6741_out1 XOR Logical_Operator_out6869_out1;

  Logical_Operator_out8854_out1 <= Logical_Operator_out6742_out1 XOR Logical_Operator_out6870_out1;

  Logical_Operator_out8855_out1 <= Logical_Operator_out6743_out1 XOR Logical_Operator_out6871_out1;

  Logical_Operator_out8856_out1 <= Logical_Operator_out6744_out1 XOR Logical_Operator_out6872_out1;

  Logical_Operator_out8857_out1 <= Logical_Operator_out6745_out1 XOR Logical_Operator_out6873_out1;

  Logical_Operator_out8858_out1 <= Logical_Operator_out6746_out1 XOR Logical_Operator_out6874_out1;

  Logical_Operator_out8859_out1 <= Logical_Operator_out6747_out1 XOR Logical_Operator_out6875_out1;

  Logical_Operator_out8860_out1 <= Logical_Operator_out6748_out1 XOR Logical_Operator_out6876_out1;

  Logical_Operator_out8861_out1 <= Logical_Operator_out6749_out1 XOR Logical_Operator_out6877_out1;

  Logical_Operator_out8862_out1 <= Logical_Operator_out6750_out1 XOR Logical_Operator_out6878_out1;

  Logical_Operator_out8863_out1 <= Logical_Operator_out6751_out1 XOR Logical_Operator_out6879_out1;

  Logical_Operator_out8864_out1 <= Logical_Operator_out6752_out1 XOR Logical_Operator_out6880_out1;

  Logical_Operator_out8865_out1 <= Logical_Operator_out6753_out1 XOR Logical_Operator_out6881_out1;

  Logical_Operator_out8866_out1 <= Logical_Operator_out6754_out1 XOR Logical_Operator_out6882_out1;

  Logical_Operator_out8867_out1 <= Logical_Operator_out6755_out1 XOR Logical_Operator_out6883_out1;

  Logical_Operator_out8868_out1 <= Logical_Operator_out6756_out1 XOR Logical_Operator_out6884_out1;

  Logical_Operator_out8869_out1 <= Logical_Operator_out6757_out1 XOR Logical_Operator_out6885_out1;

  Logical_Operator_out8870_out1 <= Logical_Operator_out6758_out1 XOR Logical_Operator_out6886_out1;

  Logical_Operator_out8871_out1 <= Logical_Operator_out6759_out1 XOR Logical_Operator_out6887_out1;

  Logical_Operator_out8872_out1 <= Logical_Operator_out6760_out1 XOR Logical_Operator_out6888_out1;

  Logical_Operator_out8873_out1 <= Logical_Operator_out6761_out1 XOR Logical_Operator_out6889_out1;

  Logical_Operator_out8874_out1 <= Logical_Operator_out6762_out1 XOR Logical_Operator_out6890_out1;

  Logical_Operator_out8875_out1 <= Logical_Operator_out6763_out1 XOR Logical_Operator_out6891_out1;

  Logical_Operator_out8876_out1 <= Logical_Operator_out6764_out1 XOR Logical_Operator_out6892_out1;

  Logical_Operator_out8877_out1 <= Logical_Operator_out6765_out1 XOR Logical_Operator_out6893_out1;

  Logical_Operator_out8878_out1 <= Logical_Operator_out6766_out1 XOR Logical_Operator_out6894_out1;

  Logical_Operator_out8879_out1 <= Logical_Operator_out6767_out1 XOR Logical_Operator_out6895_out1;

  Logical_Operator_out8880_out1 <= Logical_Operator_out6768_out1 XOR Logical_Operator_out6896_out1;

  Logical_Operator_out8881_out1 <= Logical_Operator_out6769_out1 XOR Logical_Operator_out6897_out1;

  Logical_Operator_out8882_out1 <= Logical_Operator_out6770_out1 XOR Logical_Operator_out6898_out1;

  Logical_Operator_out8883_out1 <= Logical_Operator_out6771_out1 XOR Logical_Operator_out6899_out1;

  Logical_Operator_out8884_out1 <= Logical_Operator_out6772_out1 XOR Logical_Operator_out6900_out1;

  Logical_Operator_out8885_out1 <= Logical_Operator_out6773_out1 XOR Logical_Operator_out6901_out1;

  Logical_Operator_out8886_out1 <= Logical_Operator_out6774_out1 XOR Logical_Operator_out6902_out1;

  Logical_Operator_out8887_out1 <= Logical_Operator_out6775_out1 XOR Logical_Operator_out6903_out1;

  Logical_Operator_out8888_out1 <= Logical_Operator_out6776_out1 XOR Logical_Operator_out6904_out1;

  Logical_Operator_out8889_out1 <= Logical_Operator_out6777_out1 XOR Logical_Operator_out6905_out1;

  Logical_Operator_out8890_out1 <= Logical_Operator_out6778_out1 XOR Logical_Operator_out6906_out1;

  Logical_Operator_out8891_out1 <= Logical_Operator_out6779_out1 XOR Logical_Operator_out6907_out1;

  Logical_Operator_out8892_out1 <= Logical_Operator_out6780_out1 XOR Logical_Operator_out6908_out1;

  Logical_Operator_out8893_out1 <= Logical_Operator_out6781_out1 XOR Logical_Operator_out6909_out1;

  Logical_Operator_out8894_out1 <= Logical_Operator_out6782_out1 XOR Logical_Operator_out6910_out1;

  Logical_Operator_out8895_out1 <= Logical_Operator_out6783_out1 XOR Logical_Operator_out6911_out1;

  Logical_Operator_out8896_out1 <= Logical_Operator_out6784_out1 XOR Logical_Operator_out6912_out1;

  Logical_Operator_out8897_out1 <= Logical_Operator_out5729_out1 XOR Logical_Operator_out5857_out1;

  Logical_Operator_out8898_out1 <= Logical_Operator_out5730_out1 XOR Logical_Operator_out5858_out1;

  Logical_Operator_out8899_out1 <= Logical_Operator_out5731_out1 XOR Logical_Operator_out5859_out1;

  Logical_Operator_out8900_out1 <= Logical_Operator_out5732_out1 XOR Logical_Operator_out5860_out1;

  Logical_Operator_out8901_out1 <= Logical_Operator_out5733_out1 XOR Logical_Operator_out5861_out1;

  Logical_Operator_out8902_out1 <= Logical_Operator_out5734_out1 XOR Logical_Operator_out5862_out1;

  Logical_Operator_out8903_out1 <= Logical_Operator_out5735_out1 XOR Logical_Operator_out5863_out1;

  Logical_Operator_out8904_out1 <= Logical_Operator_out5736_out1 XOR Logical_Operator_out5864_out1;

  Logical_Operator_out8905_out1 <= Logical_Operator_out5737_out1 XOR Logical_Operator_out5865_out1;

  Logical_Operator_out8906_out1 <= Logical_Operator_out5738_out1 XOR Logical_Operator_out5866_out1;

  Logical_Operator_out8907_out1 <= Logical_Operator_out5739_out1 XOR Logical_Operator_out5867_out1;

  Logical_Operator_out8908_out1 <= Logical_Operator_out5740_out1 XOR Logical_Operator_out5868_out1;

  Logical_Operator_out8909_out1 <= Logical_Operator_out5741_out1 XOR Logical_Operator_out5869_out1;

  Logical_Operator_out8910_out1 <= Logical_Operator_out5742_out1 XOR Logical_Operator_out5870_out1;

  Logical_Operator_out8911_out1 <= Logical_Operator_out5743_out1 XOR Logical_Operator_out5871_out1;

  Logical_Operator_out8912_out1 <= Logical_Operator_out5744_out1 XOR Logical_Operator_out5872_out1;

  Logical_Operator_out8913_out1 <= Logical_Operator_out5745_out1 XOR Logical_Operator_out5873_out1;

  Logical_Operator_out8914_out1 <= Logical_Operator_out5746_out1 XOR Logical_Operator_out5874_out1;

  Logical_Operator_out8915_out1 <= Logical_Operator_out5747_out1 XOR Logical_Operator_out5875_out1;

  Logical_Operator_out8916_out1 <= Logical_Operator_out5748_out1 XOR Logical_Operator_out5876_out1;

  Logical_Operator_out8917_out1 <= Logical_Operator_out5749_out1 XOR Logical_Operator_out5877_out1;

  Logical_Operator_out8918_out1 <= Logical_Operator_out5750_out1 XOR Logical_Operator_out5878_out1;

  Logical_Operator_out8919_out1 <= Logical_Operator_out5751_out1 XOR Logical_Operator_out5879_out1;

  Logical_Operator_out8920_out1 <= Logical_Operator_out5752_out1 XOR Logical_Operator_out5880_out1;

  Logical_Operator_out8921_out1 <= Logical_Operator_out5753_out1 XOR Logical_Operator_out5881_out1;

  Logical_Operator_out8922_out1 <= Logical_Operator_out5754_out1 XOR Logical_Operator_out5882_out1;

  Logical_Operator_out8923_out1 <= Logical_Operator_out5755_out1 XOR Logical_Operator_out5883_out1;

  Logical_Operator_out8924_out1 <= Logical_Operator_out5756_out1 XOR Logical_Operator_out5884_out1;

  Logical_Operator_out8925_out1 <= Logical_Operator_out5757_out1 XOR Logical_Operator_out5885_out1;

  Logical_Operator_out8926_out1 <= Logical_Operator_out5758_out1 XOR Logical_Operator_out5886_out1;

  Logical_Operator_out8927_out1 <= Logical_Operator_out5759_out1 XOR Logical_Operator_out5887_out1;

  Logical_Operator_out8928_out1 <= Logical_Operator_out5760_out1 XOR Logical_Operator_out5888_out1;

  Logical_Operator_out8929_out1 <= Logical_Operator_out4721_out1 XOR Logical_Operator_out4849_out1;

  Logical_Operator_out8930_out1 <= Logical_Operator_out4722_out1 XOR Logical_Operator_out4850_out1;

  Logical_Operator_out8931_out1 <= Logical_Operator_out4723_out1 XOR Logical_Operator_out4851_out1;

  Logical_Operator_out8932_out1 <= Logical_Operator_out4724_out1 XOR Logical_Operator_out4852_out1;

  Logical_Operator_out8933_out1 <= Logical_Operator_out4725_out1 XOR Logical_Operator_out4853_out1;

  Logical_Operator_out8934_out1 <= Logical_Operator_out4726_out1 XOR Logical_Operator_out4854_out1;

  Logical_Operator_out8935_out1 <= Logical_Operator_out4727_out1 XOR Logical_Operator_out4855_out1;

  Logical_Operator_out8936_out1 <= Logical_Operator_out4728_out1 XOR Logical_Operator_out4856_out1;

  Logical_Operator_out8937_out1 <= Logical_Operator_out4729_out1 XOR Logical_Operator_out4857_out1;

  Logical_Operator_out8938_out1 <= Logical_Operator_out4730_out1 XOR Logical_Operator_out4858_out1;

  Logical_Operator_out8939_out1 <= Logical_Operator_out4731_out1 XOR Logical_Operator_out4859_out1;

  Logical_Operator_out8940_out1 <= Logical_Operator_out4732_out1 XOR Logical_Operator_out4860_out1;

  Logical_Operator_out8941_out1 <= Logical_Operator_out4733_out1 XOR Logical_Operator_out4861_out1;

  Logical_Operator_out8942_out1 <= Logical_Operator_out4734_out1 XOR Logical_Operator_out4862_out1;

  Logical_Operator_out8943_out1 <= Logical_Operator_out4735_out1 XOR Logical_Operator_out4863_out1;

  Logical_Operator_out8944_out1 <= Logical_Operator_out4736_out1 XOR Logical_Operator_out4864_out1;

  Logical_Operator_out8945_out1 <= Logical_Operator_out3705_out1 XOR Logical_Operator_out3833_out1;

  Logical_Operator_out8946_out1 <= Logical_Operator_out3706_out1 XOR Logical_Operator_out3834_out1;

  Logical_Operator_out8947_out1 <= Logical_Operator_out3707_out1 XOR Logical_Operator_out3835_out1;

  Logical_Operator_out8948_out1 <= Logical_Operator_out3708_out1 XOR Logical_Operator_out3836_out1;

  Logical_Operator_out8949_out1 <= Logical_Operator_out3709_out1 XOR Logical_Operator_out3837_out1;

  Logical_Operator_out8950_out1 <= Logical_Operator_out3710_out1 XOR Logical_Operator_out3838_out1;

  Logical_Operator_out8951_out1 <= Logical_Operator_out3711_out1 XOR Logical_Operator_out3839_out1;

  Logical_Operator_out8952_out1 <= Logical_Operator_out3712_out1 XOR Logical_Operator_out3840_out1;

  Logical_Operator_out8953_out1 <= Logical_Operator_out2685_out1 XOR Logical_Operator_out2813_out1;

  Logical_Operator_out8954_out1 <= Logical_Operator_out2686_out1 XOR Logical_Operator_out2814_out1;

  Logical_Operator_out8955_out1 <= Logical_Operator_out2687_out1 XOR Logical_Operator_out2815_out1;

  Logical_Operator_out8956_out1 <= Logical_Operator_out2688_out1 XOR Logical_Operator_out2816_out1;

  Logical_Operator_out8957_out1 <= Logical_Operator_out1663_out1 XOR Logical_Operator_out1791_out1;

  Logical_Operator_out8958_out1 <= Logical_Operator_out1664_out1 XOR Logical_Operator_out1792_out1;

  Logical_Operator_out8959_out1 <= Logical_Operator_out640_out1 XOR Logical_Operator_out768_out1;

  Logical_Operator_out8960_out1 <= in1280 XOR in1536;

  Logical_Operator_out8961_out1 <= Logical_Operator_out7937_out1 XOR Logical_Operator_out8065_out1;

  Logical_Operator_out8962_out1 <= Logical_Operator_out7938_out1 XOR Logical_Operator_out8066_out1;

  Logical_Operator_out8963_out1 <= Logical_Operator_out7939_out1 XOR Logical_Operator_out8067_out1;

  Logical_Operator_out8964_out1 <= Logical_Operator_out7940_out1 XOR Logical_Operator_out8068_out1;

  Logical_Operator_out8965_out1 <= Logical_Operator_out7941_out1 XOR Logical_Operator_out8069_out1;

  Logical_Operator_out8966_out1 <= Logical_Operator_out7942_out1 XOR Logical_Operator_out8070_out1;

  Logical_Operator_out8967_out1 <= Logical_Operator_out7943_out1 XOR Logical_Operator_out8071_out1;

  Logical_Operator_out8968_out1 <= Logical_Operator_out7944_out1 XOR Logical_Operator_out8072_out1;

  Logical_Operator_out8969_out1 <= Logical_Operator_out7945_out1 XOR Logical_Operator_out8073_out1;

  Logical_Operator_out8970_out1 <= Logical_Operator_out7946_out1 XOR Logical_Operator_out8074_out1;

  Logical_Operator_out8971_out1 <= Logical_Operator_out7947_out1 XOR Logical_Operator_out8075_out1;

  Logical_Operator_out8972_out1 <= Logical_Operator_out7948_out1 XOR Logical_Operator_out8076_out1;

  Logical_Operator_out8973_out1 <= Logical_Operator_out7949_out1 XOR Logical_Operator_out8077_out1;

  Logical_Operator_out8974_out1 <= Logical_Operator_out7950_out1 XOR Logical_Operator_out8078_out1;

  Logical_Operator_out8975_out1 <= Logical_Operator_out7951_out1 XOR Logical_Operator_out8079_out1;

  Logical_Operator_out8976_out1 <= Logical_Operator_out7952_out1 XOR Logical_Operator_out8080_out1;

  Logical_Operator_out8977_out1 <= Logical_Operator_out7953_out1 XOR Logical_Operator_out8081_out1;

  Logical_Operator_out8978_out1 <= Logical_Operator_out7954_out1 XOR Logical_Operator_out8082_out1;

  Logical_Operator_out8979_out1 <= Logical_Operator_out7955_out1 XOR Logical_Operator_out8083_out1;

  Logical_Operator_out8980_out1 <= Logical_Operator_out7956_out1 XOR Logical_Operator_out8084_out1;

  Logical_Operator_out8981_out1 <= Logical_Operator_out7957_out1 XOR Logical_Operator_out8085_out1;

  Logical_Operator_out8982_out1 <= Logical_Operator_out7958_out1 XOR Logical_Operator_out8086_out1;

  Logical_Operator_out8983_out1 <= Logical_Operator_out7959_out1 XOR Logical_Operator_out8087_out1;

  Logical_Operator_out8984_out1 <= Logical_Operator_out7960_out1 XOR Logical_Operator_out8088_out1;

  Logical_Operator_out8985_out1 <= Logical_Operator_out7961_out1 XOR Logical_Operator_out8089_out1;

  Logical_Operator_out8986_out1 <= Logical_Operator_out7962_out1 XOR Logical_Operator_out8090_out1;

  Logical_Operator_out8987_out1 <= Logical_Operator_out7963_out1 XOR Logical_Operator_out8091_out1;

  Logical_Operator_out8988_out1 <= Logical_Operator_out7964_out1 XOR Logical_Operator_out8092_out1;

  Logical_Operator_out8989_out1 <= Logical_Operator_out7965_out1 XOR Logical_Operator_out8093_out1;

  Logical_Operator_out8990_out1 <= Logical_Operator_out7966_out1 XOR Logical_Operator_out8094_out1;

  Logical_Operator_out8991_out1 <= Logical_Operator_out7967_out1 XOR Logical_Operator_out8095_out1;

  Logical_Operator_out8992_out1 <= Logical_Operator_out7968_out1 XOR Logical_Operator_out8096_out1;

  Logical_Operator_out8993_out1 <= Logical_Operator_out7969_out1 XOR Logical_Operator_out8097_out1;

  Logical_Operator_out8994_out1 <= Logical_Operator_out7970_out1 XOR Logical_Operator_out8098_out1;

  Logical_Operator_out8995_out1 <= Logical_Operator_out7971_out1 XOR Logical_Operator_out8099_out1;

  Logical_Operator_out8996_out1 <= Logical_Operator_out7972_out1 XOR Logical_Operator_out8100_out1;

  Logical_Operator_out8997_out1 <= Logical_Operator_out7973_out1 XOR Logical_Operator_out8101_out1;

  Logical_Operator_out8998_out1 <= Logical_Operator_out7974_out1 XOR Logical_Operator_out8102_out1;

  Logical_Operator_out8999_out1 <= Logical_Operator_out7975_out1 XOR Logical_Operator_out8103_out1;

  Logical_Operator_out9000_out1 <= Logical_Operator_out7976_out1 XOR Logical_Operator_out8104_out1;

  Logical_Operator_out9001_out1 <= Logical_Operator_out7977_out1 XOR Logical_Operator_out8105_out1;

  Logical_Operator_out9002_out1 <= Logical_Operator_out7978_out1 XOR Logical_Operator_out8106_out1;

  Logical_Operator_out9003_out1 <= Logical_Operator_out7979_out1 XOR Logical_Operator_out8107_out1;

  Logical_Operator_out9004_out1 <= Logical_Operator_out7980_out1 XOR Logical_Operator_out8108_out1;

  Logical_Operator_out9005_out1 <= Logical_Operator_out7981_out1 XOR Logical_Operator_out8109_out1;

  Logical_Operator_out9006_out1 <= Logical_Operator_out7982_out1 XOR Logical_Operator_out8110_out1;

  Logical_Operator_out9007_out1 <= Logical_Operator_out7983_out1 XOR Logical_Operator_out8111_out1;

  Logical_Operator_out9008_out1 <= Logical_Operator_out7984_out1 XOR Logical_Operator_out8112_out1;

  Logical_Operator_out9009_out1 <= Logical_Operator_out7985_out1 XOR Logical_Operator_out8113_out1;

  Logical_Operator_out9010_out1 <= Logical_Operator_out7986_out1 XOR Logical_Operator_out8114_out1;

  Logical_Operator_out9011_out1 <= Logical_Operator_out7987_out1 XOR Logical_Operator_out8115_out1;

  Logical_Operator_out9012_out1 <= Logical_Operator_out7988_out1 XOR Logical_Operator_out8116_out1;

  Logical_Operator_out9013_out1 <= Logical_Operator_out7989_out1 XOR Logical_Operator_out8117_out1;

  Logical_Operator_out9014_out1 <= Logical_Operator_out7990_out1 XOR Logical_Operator_out8118_out1;

  Logical_Operator_out9015_out1 <= Logical_Operator_out7991_out1 XOR Logical_Operator_out8119_out1;

  Logical_Operator_out9016_out1 <= Logical_Operator_out7992_out1 XOR Logical_Operator_out8120_out1;

  Logical_Operator_out9017_out1 <= Logical_Operator_out7993_out1 XOR Logical_Operator_out8121_out1;

  Logical_Operator_out9018_out1 <= Logical_Operator_out7994_out1 XOR Logical_Operator_out8122_out1;

  Logical_Operator_out9019_out1 <= Logical_Operator_out7995_out1 XOR Logical_Operator_out8123_out1;

  Logical_Operator_out9020_out1 <= Logical_Operator_out7996_out1 XOR Logical_Operator_out8124_out1;

  Logical_Operator_out9021_out1 <= Logical_Operator_out7997_out1 XOR Logical_Operator_out8125_out1;

  Logical_Operator_out9022_out1 <= Logical_Operator_out7998_out1 XOR Logical_Operator_out8126_out1;

  Logical_Operator_out9023_out1 <= Logical_Operator_out7999_out1 XOR Logical_Operator_out8127_out1;

  Logical_Operator_out9024_out1 <= Logical_Operator_out8000_out1 XOR Logical_Operator_out8128_out1;

  Logical_Operator_out9025_out1 <= Logical_Operator_out8001_out1 XOR Logical_Operator_out8129_out1;

  Logical_Operator_out9026_out1 <= Logical_Operator_out8002_out1 XOR Logical_Operator_out8130_out1;

  Logical_Operator_out9027_out1 <= Logical_Operator_out8003_out1 XOR Logical_Operator_out8131_out1;

  Logical_Operator_out9028_out1 <= Logical_Operator_out8004_out1 XOR Logical_Operator_out8132_out1;

  Logical_Operator_out9029_out1 <= Logical_Operator_out8005_out1 XOR Logical_Operator_out8133_out1;

  Logical_Operator_out9030_out1 <= Logical_Operator_out8006_out1 XOR Logical_Operator_out8134_out1;

  Logical_Operator_out9031_out1 <= Logical_Operator_out8007_out1 XOR Logical_Operator_out8135_out1;

  Logical_Operator_out9032_out1 <= Logical_Operator_out8008_out1 XOR Logical_Operator_out8136_out1;

  Logical_Operator_out9033_out1 <= Logical_Operator_out8009_out1 XOR Logical_Operator_out8137_out1;

  Logical_Operator_out9034_out1 <= Logical_Operator_out8010_out1 XOR Logical_Operator_out8138_out1;

  Logical_Operator_out9035_out1 <= Logical_Operator_out8011_out1 XOR Logical_Operator_out8139_out1;

  Logical_Operator_out9036_out1 <= Logical_Operator_out8012_out1 XOR Logical_Operator_out8140_out1;

  Logical_Operator_out9037_out1 <= Logical_Operator_out8013_out1 XOR Logical_Operator_out8141_out1;

  Logical_Operator_out9038_out1 <= Logical_Operator_out8014_out1 XOR Logical_Operator_out8142_out1;

  Logical_Operator_out9039_out1 <= Logical_Operator_out8015_out1 XOR Logical_Operator_out8143_out1;

  Logical_Operator_out9040_out1 <= Logical_Operator_out8016_out1 XOR Logical_Operator_out8144_out1;

  Logical_Operator_out9041_out1 <= Logical_Operator_out8017_out1 XOR Logical_Operator_out8145_out1;

  Logical_Operator_out9042_out1 <= Logical_Operator_out8018_out1 XOR Logical_Operator_out8146_out1;

  Logical_Operator_out9043_out1 <= Logical_Operator_out8019_out1 XOR Logical_Operator_out8147_out1;

  Logical_Operator_out9044_out1 <= Logical_Operator_out8020_out1 XOR Logical_Operator_out8148_out1;

  Logical_Operator_out9045_out1 <= Logical_Operator_out8021_out1 XOR Logical_Operator_out8149_out1;

  Logical_Operator_out9046_out1 <= Logical_Operator_out8022_out1 XOR Logical_Operator_out8150_out1;

  Logical_Operator_out9047_out1 <= Logical_Operator_out8023_out1 XOR Logical_Operator_out8151_out1;

  Logical_Operator_out9048_out1 <= Logical_Operator_out8024_out1 XOR Logical_Operator_out8152_out1;

  Logical_Operator_out9049_out1 <= Logical_Operator_out8025_out1 XOR Logical_Operator_out8153_out1;

  Logical_Operator_out9050_out1 <= Logical_Operator_out8026_out1 XOR Logical_Operator_out8154_out1;

  Logical_Operator_out9051_out1 <= Logical_Operator_out8027_out1 XOR Logical_Operator_out8155_out1;

  Logical_Operator_out9052_out1 <= Logical_Operator_out8028_out1 XOR Logical_Operator_out8156_out1;

  Logical_Operator_out9053_out1 <= Logical_Operator_out8029_out1 XOR Logical_Operator_out8157_out1;

  Logical_Operator_out9054_out1 <= Logical_Operator_out8030_out1 XOR Logical_Operator_out8158_out1;

  Logical_Operator_out9055_out1 <= Logical_Operator_out8031_out1 XOR Logical_Operator_out8159_out1;

  Logical_Operator_out9056_out1 <= Logical_Operator_out8032_out1 XOR Logical_Operator_out8160_out1;

  Logical_Operator_out9057_out1 <= Logical_Operator_out8033_out1 XOR Logical_Operator_out8161_out1;

  Logical_Operator_out9058_out1 <= Logical_Operator_out8034_out1 XOR Logical_Operator_out8162_out1;

  Logical_Operator_out9059_out1 <= Logical_Operator_out8035_out1 XOR Logical_Operator_out8163_out1;

  Logical_Operator_out9060_out1 <= Logical_Operator_out8036_out1 XOR Logical_Operator_out8164_out1;

  Logical_Operator_out9061_out1 <= Logical_Operator_out8037_out1 XOR Logical_Operator_out8165_out1;

  Logical_Operator_out9062_out1 <= Logical_Operator_out8038_out1 XOR Logical_Operator_out8166_out1;

  Logical_Operator_out9063_out1 <= Logical_Operator_out8039_out1 XOR Logical_Operator_out8167_out1;

  Logical_Operator_out9064_out1 <= Logical_Operator_out8040_out1 XOR Logical_Operator_out8168_out1;

  Logical_Operator_out9065_out1 <= Logical_Operator_out8041_out1 XOR Logical_Operator_out8169_out1;

  Logical_Operator_out9066_out1 <= Logical_Operator_out8042_out1 XOR Logical_Operator_out8170_out1;

  Logical_Operator_out9067_out1 <= Logical_Operator_out8043_out1 XOR Logical_Operator_out8171_out1;

  Logical_Operator_out9068_out1 <= Logical_Operator_out8044_out1 XOR Logical_Operator_out8172_out1;

  Logical_Operator_out9069_out1 <= Logical_Operator_out8045_out1 XOR Logical_Operator_out8173_out1;

  Logical_Operator_out9070_out1 <= Logical_Operator_out8046_out1 XOR Logical_Operator_out8174_out1;

  Logical_Operator_out9071_out1 <= Logical_Operator_out8047_out1 XOR Logical_Operator_out8175_out1;

  Logical_Operator_out9072_out1 <= Logical_Operator_out8048_out1 XOR Logical_Operator_out8176_out1;

  Logical_Operator_out9073_out1 <= Logical_Operator_out8049_out1 XOR Logical_Operator_out8177_out1;

  Logical_Operator_out9074_out1 <= Logical_Operator_out8050_out1 XOR Logical_Operator_out8178_out1;

  Logical_Operator_out9075_out1 <= Logical_Operator_out8051_out1 XOR Logical_Operator_out8179_out1;

  Logical_Operator_out9076_out1 <= Logical_Operator_out8052_out1 XOR Logical_Operator_out8180_out1;

  Logical_Operator_out9077_out1 <= Logical_Operator_out8053_out1 XOR Logical_Operator_out8181_out1;

  Logical_Operator_out9078_out1 <= Logical_Operator_out8054_out1 XOR Logical_Operator_out8182_out1;

  Logical_Operator_out9079_out1 <= Logical_Operator_out8055_out1 XOR Logical_Operator_out8183_out1;

  Logical_Operator_out9080_out1 <= Logical_Operator_out8056_out1 XOR Logical_Operator_out8184_out1;

  Logical_Operator_out9081_out1 <= Logical_Operator_out8057_out1 XOR Logical_Operator_out8185_out1;

  Logical_Operator_out9082_out1 <= Logical_Operator_out8058_out1 XOR Logical_Operator_out8186_out1;

  Logical_Operator_out9083_out1 <= Logical_Operator_out8059_out1 XOR Logical_Operator_out8187_out1;

  Logical_Operator_out9084_out1 <= Logical_Operator_out8060_out1 XOR Logical_Operator_out8188_out1;

  Logical_Operator_out9085_out1 <= Logical_Operator_out8061_out1 XOR Logical_Operator_out8189_out1;

  Logical_Operator_out9086_out1 <= Logical_Operator_out8062_out1 XOR Logical_Operator_out8190_out1;

  Logical_Operator_out9087_out1 <= Logical_Operator_out8063_out1 XOR Logical_Operator_out8191_out1;

  Logical_Operator_out9088_out1 <= Logical_Operator_out8064_out1 XOR Logical_Operator_out8192_out1;

  Logical_Operator_out9089_out1 <= Logical_Operator_out6977_out1 XOR Logical_Operator_out7105_out1;

  Logical_Operator_out9090_out1 <= Logical_Operator_out6978_out1 XOR Logical_Operator_out7106_out1;

  Logical_Operator_out9091_out1 <= Logical_Operator_out6979_out1 XOR Logical_Operator_out7107_out1;

  Logical_Operator_out9092_out1 <= Logical_Operator_out6980_out1 XOR Logical_Operator_out7108_out1;

  Logical_Operator_out9093_out1 <= Logical_Operator_out6981_out1 XOR Logical_Operator_out7109_out1;

  Logical_Operator_out9094_out1 <= Logical_Operator_out6982_out1 XOR Logical_Operator_out7110_out1;

  Logical_Operator_out9095_out1 <= Logical_Operator_out6983_out1 XOR Logical_Operator_out7111_out1;

  Logical_Operator_out9096_out1 <= Logical_Operator_out6984_out1 XOR Logical_Operator_out7112_out1;

  Logical_Operator_out9097_out1 <= Logical_Operator_out6985_out1 XOR Logical_Operator_out7113_out1;

  Logical_Operator_out9098_out1 <= Logical_Operator_out6986_out1 XOR Logical_Operator_out7114_out1;

  Logical_Operator_out9099_out1 <= Logical_Operator_out6987_out1 XOR Logical_Operator_out7115_out1;

  Logical_Operator_out9100_out1 <= Logical_Operator_out6988_out1 XOR Logical_Operator_out7116_out1;

  Logical_Operator_out9101_out1 <= Logical_Operator_out6989_out1 XOR Logical_Operator_out7117_out1;

  Logical_Operator_out9102_out1 <= Logical_Operator_out6990_out1 XOR Logical_Operator_out7118_out1;

  Logical_Operator_out9103_out1 <= Logical_Operator_out6991_out1 XOR Logical_Operator_out7119_out1;

  Logical_Operator_out9104_out1 <= Logical_Operator_out6992_out1 XOR Logical_Operator_out7120_out1;

  Logical_Operator_out9105_out1 <= Logical_Operator_out6993_out1 XOR Logical_Operator_out7121_out1;

  Logical_Operator_out9106_out1 <= Logical_Operator_out6994_out1 XOR Logical_Operator_out7122_out1;

  Logical_Operator_out9107_out1 <= Logical_Operator_out6995_out1 XOR Logical_Operator_out7123_out1;

  Logical_Operator_out9108_out1 <= Logical_Operator_out6996_out1 XOR Logical_Operator_out7124_out1;

  Logical_Operator_out9109_out1 <= Logical_Operator_out6997_out1 XOR Logical_Operator_out7125_out1;

  Logical_Operator_out9110_out1 <= Logical_Operator_out6998_out1 XOR Logical_Operator_out7126_out1;

  Logical_Operator_out9111_out1 <= Logical_Operator_out6999_out1 XOR Logical_Operator_out7127_out1;

  Logical_Operator_out9112_out1 <= Logical_Operator_out7000_out1 XOR Logical_Operator_out7128_out1;

  Logical_Operator_out9113_out1 <= Logical_Operator_out7001_out1 XOR Logical_Operator_out7129_out1;

  Logical_Operator_out9114_out1 <= Logical_Operator_out7002_out1 XOR Logical_Operator_out7130_out1;

  Logical_Operator_out9115_out1 <= Logical_Operator_out7003_out1 XOR Logical_Operator_out7131_out1;

  Logical_Operator_out9116_out1 <= Logical_Operator_out7004_out1 XOR Logical_Operator_out7132_out1;

  Logical_Operator_out9117_out1 <= Logical_Operator_out7005_out1 XOR Logical_Operator_out7133_out1;

  Logical_Operator_out9118_out1 <= Logical_Operator_out7006_out1 XOR Logical_Operator_out7134_out1;

  Logical_Operator_out9119_out1 <= Logical_Operator_out7007_out1 XOR Logical_Operator_out7135_out1;

  Logical_Operator_out9120_out1 <= Logical_Operator_out7008_out1 XOR Logical_Operator_out7136_out1;

  Logical_Operator_out9121_out1 <= Logical_Operator_out7009_out1 XOR Logical_Operator_out7137_out1;

  Logical_Operator_out9122_out1 <= Logical_Operator_out7010_out1 XOR Logical_Operator_out7138_out1;

  Logical_Operator_out9123_out1 <= Logical_Operator_out7011_out1 XOR Logical_Operator_out7139_out1;

  Logical_Operator_out9124_out1 <= Logical_Operator_out7012_out1 XOR Logical_Operator_out7140_out1;

  Logical_Operator_out9125_out1 <= Logical_Operator_out7013_out1 XOR Logical_Operator_out7141_out1;

  Logical_Operator_out9126_out1 <= Logical_Operator_out7014_out1 XOR Logical_Operator_out7142_out1;

  Logical_Operator_out9127_out1 <= Logical_Operator_out7015_out1 XOR Logical_Operator_out7143_out1;

  Logical_Operator_out9128_out1 <= Logical_Operator_out7016_out1 XOR Logical_Operator_out7144_out1;

  Logical_Operator_out9129_out1 <= Logical_Operator_out7017_out1 XOR Logical_Operator_out7145_out1;

  Logical_Operator_out9130_out1 <= Logical_Operator_out7018_out1 XOR Logical_Operator_out7146_out1;

  Logical_Operator_out9131_out1 <= Logical_Operator_out7019_out1 XOR Logical_Operator_out7147_out1;

  Logical_Operator_out9132_out1 <= Logical_Operator_out7020_out1 XOR Logical_Operator_out7148_out1;

  Logical_Operator_out9133_out1 <= Logical_Operator_out7021_out1 XOR Logical_Operator_out7149_out1;

  Logical_Operator_out9134_out1 <= Logical_Operator_out7022_out1 XOR Logical_Operator_out7150_out1;

  Logical_Operator_out9135_out1 <= Logical_Operator_out7023_out1 XOR Logical_Operator_out7151_out1;

  Logical_Operator_out9136_out1 <= Logical_Operator_out7024_out1 XOR Logical_Operator_out7152_out1;

  Logical_Operator_out9137_out1 <= Logical_Operator_out7025_out1 XOR Logical_Operator_out7153_out1;

  Logical_Operator_out9138_out1 <= Logical_Operator_out7026_out1 XOR Logical_Operator_out7154_out1;

  Logical_Operator_out9139_out1 <= Logical_Operator_out7027_out1 XOR Logical_Operator_out7155_out1;

  Logical_Operator_out9140_out1 <= Logical_Operator_out7028_out1 XOR Logical_Operator_out7156_out1;

  Logical_Operator_out9141_out1 <= Logical_Operator_out7029_out1 XOR Logical_Operator_out7157_out1;

  Logical_Operator_out9142_out1 <= Logical_Operator_out7030_out1 XOR Logical_Operator_out7158_out1;

  Logical_Operator_out9143_out1 <= Logical_Operator_out7031_out1 XOR Logical_Operator_out7159_out1;

  Logical_Operator_out9144_out1 <= Logical_Operator_out7032_out1 XOR Logical_Operator_out7160_out1;

  Logical_Operator_out9145_out1 <= Logical_Operator_out7033_out1 XOR Logical_Operator_out7161_out1;

  Logical_Operator_out9146_out1 <= Logical_Operator_out7034_out1 XOR Logical_Operator_out7162_out1;

  Logical_Operator_out9147_out1 <= Logical_Operator_out7035_out1 XOR Logical_Operator_out7163_out1;

  Logical_Operator_out9148_out1 <= Logical_Operator_out7036_out1 XOR Logical_Operator_out7164_out1;

  Logical_Operator_out9149_out1 <= Logical_Operator_out7037_out1 XOR Logical_Operator_out7165_out1;

  Logical_Operator_out9150_out1 <= Logical_Operator_out7038_out1 XOR Logical_Operator_out7166_out1;

  Logical_Operator_out9151_out1 <= Logical_Operator_out7039_out1 XOR Logical_Operator_out7167_out1;

  Logical_Operator_out9152_out1 <= Logical_Operator_out7040_out1 XOR Logical_Operator_out7168_out1;

  Logical_Operator_out9153_out1 <= Logical_Operator_out5985_out1 XOR Logical_Operator_out6113_out1;

  Logical_Operator_out9154_out1 <= Logical_Operator_out5986_out1 XOR Logical_Operator_out6114_out1;

  Logical_Operator_out9155_out1 <= Logical_Operator_out5987_out1 XOR Logical_Operator_out6115_out1;

  Logical_Operator_out9156_out1 <= Logical_Operator_out5988_out1 XOR Logical_Operator_out6116_out1;

  Logical_Operator_out9157_out1 <= Logical_Operator_out5989_out1 XOR Logical_Operator_out6117_out1;

  Logical_Operator_out9158_out1 <= Logical_Operator_out5990_out1 XOR Logical_Operator_out6118_out1;

  Logical_Operator_out9159_out1 <= Logical_Operator_out5991_out1 XOR Logical_Operator_out6119_out1;

  Logical_Operator_out9160_out1 <= Logical_Operator_out5992_out1 XOR Logical_Operator_out6120_out1;

  Logical_Operator_out9161_out1 <= Logical_Operator_out5993_out1 XOR Logical_Operator_out6121_out1;

  Logical_Operator_out9162_out1 <= Logical_Operator_out5994_out1 XOR Logical_Operator_out6122_out1;

  Logical_Operator_out9163_out1 <= Logical_Operator_out5995_out1 XOR Logical_Operator_out6123_out1;

  Logical_Operator_out9164_out1 <= Logical_Operator_out5996_out1 XOR Logical_Operator_out6124_out1;

  Logical_Operator_out9165_out1 <= Logical_Operator_out5997_out1 XOR Logical_Operator_out6125_out1;

  Logical_Operator_out9166_out1 <= Logical_Operator_out5998_out1 XOR Logical_Operator_out6126_out1;

  Logical_Operator_out9167_out1 <= Logical_Operator_out5999_out1 XOR Logical_Operator_out6127_out1;

  Logical_Operator_out9168_out1 <= Logical_Operator_out6000_out1 XOR Logical_Operator_out6128_out1;

  Logical_Operator_out9169_out1 <= Logical_Operator_out6001_out1 XOR Logical_Operator_out6129_out1;

  Logical_Operator_out9170_out1 <= Logical_Operator_out6002_out1 XOR Logical_Operator_out6130_out1;

  Logical_Operator_out9171_out1 <= Logical_Operator_out6003_out1 XOR Logical_Operator_out6131_out1;

  Logical_Operator_out9172_out1 <= Logical_Operator_out6004_out1 XOR Logical_Operator_out6132_out1;

  Logical_Operator_out9173_out1 <= Logical_Operator_out6005_out1 XOR Logical_Operator_out6133_out1;

  Logical_Operator_out9174_out1 <= Logical_Operator_out6006_out1 XOR Logical_Operator_out6134_out1;

  Logical_Operator_out9175_out1 <= Logical_Operator_out6007_out1 XOR Logical_Operator_out6135_out1;

  Logical_Operator_out9176_out1 <= Logical_Operator_out6008_out1 XOR Logical_Operator_out6136_out1;

  Logical_Operator_out9177_out1 <= Logical_Operator_out6009_out1 XOR Logical_Operator_out6137_out1;

  Logical_Operator_out9178_out1 <= Logical_Operator_out6010_out1 XOR Logical_Operator_out6138_out1;

  Logical_Operator_out9179_out1 <= Logical_Operator_out6011_out1 XOR Logical_Operator_out6139_out1;

  Logical_Operator_out9180_out1 <= Logical_Operator_out6012_out1 XOR Logical_Operator_out6140_out1;

  Logical_Operator_out9181_out1 <= Logical_Operator_out6013_out1 XOR Logical_Operator_out6141_out1;

  Logical_Operator_out9182_out1 <= Logical_Operator_out6014_out1 XOR Logical_Operator_out6142_out1;

  Logical_Operator_out9183_out1 <= Logical_Operator_out6015_out1 XOR Logical_Operator_out6143_out1;

  Logical_Operator_out9184_out1 <= Logical_Operator_out6016_out1 XOR Logical_Operator_out6144_out1;

  Logical_Operator_out9185_out1 <= Logical_Operator_out4977_out1 XOR Logical_Operator_out5105_out1;

  Logical_Operator_out9186_out1 <= Logical_Operator_out4978_out1 XOR Logical_Operator_out5106_out1;

  Logical_Operator_out9187_out1 <= Logical_Operator_out4979_out1 XOR Logical_Operator_out5107_out1;

  Logical_Operator_out9188_out1 <= Logical_Operator_out4980_out1 XOR Logical_Operator_out5108_out1;

  Logical_Operator_out9189_out1 <= Logical_Operator_out4981_out1 XOR Logical_Operator_out5109_out1;

  Logical_Operator_out9190_out1 <= Logical_Operator_out4982_out1 XOR Logical_Operator_out5110_out1;

  Logical_Operator_out9191_out1 <= Logical_Operator_out4983_out1 XOR Logical_Operator_out5111_out1;

  Logical_Operator_out9192_out1 <= Logical_Operator_out4984_out1 XOR Logical_Operator_out5112_out1;

  Logical_Operator_out9193_out1 <= Logical_Operator_out4985_out1 XOR Logical_Operator_out5113_out1;

  Logical_Operator_out9194_out1 <= Logical_Operator_out4986_out1 XOR Logical_Operator_out5114_out1;

  Logical_Operator_out9195_out1 <= Logical_Operator_out4987_out1 XOR Logical_Operator_out5115_out1;

  Logical_Operator_out9196_out1 <= Logical_Operator_out4988_out1 XOR Logical_Operator_out5116_out1;

  Logical_Operator_out9197_out1 <= Logical_Operator_out4989_out1 XOR Logical_Operator_out5117_out1;

  Logical_Operator_out9198_out1 <= Logical_Operator_out4990_out1 XOR Logical_Operator_out5118_out1;

  Logical_Operator_out9199_out1 <= Logical_Operator_out4991_out1 XOR Logical_Operator_out5119_out1;

  Logical_Operator_out9200_out1 <= Logical_Operator_out4992_out1 XOR Logical_Operator_out5120_out1;

  Logical_Operator_out9201_out1 <= Logical_Operator_out3961_out1 XOR Logical_Operator_out4089_out1;

  Logical_Operator_out9202_out1 <= Logical_Operator_out3962_out1 XOR Logical_Operator_out4090_out1;

  Logical_Operator_out9203_out1 <= Logical_Operator_out3963_out1 XOR Logical_Operator_out4091_out1;

  Logical_Operator_out9204_out1 <= Logical_Operator_out3964_out1 XOR Logical_Operator_out4092_out1;

  Logical_Operator_out9205_out1 <= Logical_Operator_out3965_out1 XOR Logical_Operator_out4093_out1;

  Logical_Operator_out9206_out1 <= Logical_Operator_out3966_out1 XOR Logical_Operator_out4094_out1;

  Logical_Operator_out9207_out1 <= Logical_Operator_out3967_out1 XOR Logical_Operator_out4095_out1;

  Logical_Operator_out9208_out1 <= Logical_Operator_out3968_out1 XOR Logical_Operator_out4096_out1;

  Logical_Operator_out9209_out1 <= Logical_Operator_out2941_out1 XOR Logical_Operator_out3069_out1;

  Logical_Operator_out9210_out1 <= Logical_Operator_out2942_out1 XOR Logical_Operator_out3070_out1;

  Logical_Operator_out9211_out1 <= Logical_Operator_out2943_out1 XOR Logical_Operator_out3071_out1;

  Logical_Operator_out9212_out1 <= Logical_Operator_out2944_out1 XOR Logical_Operator_out3072_out1;

  Logical_Operator_out9213_out1 <= Logical_Operator_out1919_out1 XOR Logical_Operator_out2047_out1;

  Logical_Operator_out9214_out1 <= Logical_Operator_out1920_out1 XOR Logical_Operator_out2048_out1;

  Logical_Operator_out9215_out1 <= Logical_Operator_out896_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out9216_out1 <= in1792 XOR in2048;

  Logical_Operator_out9217_out1 <= Logical_Operator_out8193_out1 XOR Logical_Operator_out8449_out1;

  Logical_Operator_out9218_out1 <= Logical_Operator_out8194_out1 XOR Logical_Operator_out8450_out1;

  Logical_Operator_out9219_out1 <= Logical_Operator_out8195_out1 XOR Logical_Operator_out8451_out1;

  Logical_Operator_out9220_out1 <= Logical_Operator_out8196_out1 XOR Logical_Operator_out8452_out1;

  Logical_Operator_out9221_out1 <= Logical_Operator_out8197_out1 XOR Logical_Operator_out8453_out1;

  Logical_Operator_out9222_out1 <= Logical_Operator_out8198_out1 XOR Logical_Operator_out8454_out1;

  Logical_Operator_out9223_out1 <= Logical_Operator_out8199_out1 XOR Logical_Operator_out8455_out1;

  Logical_Operator_out9224_out1 <= Logical_Operator_out8200_out1 XOR Logical_Operator_out8456_out1;

  Logical_Operator_out9225_out1 <= Logical_Operator_out8201_out1 XOR Logical_Operator_out8457_out1;

  Logical_Operator_out9226_out1 <= Logical_Operator_out8202_out1 XOR Logical_Operator_out8458_out1;

  Logical_Operator_out9227_out1 <= Logical_Operator_out8203_out1 XOR Logical_Operator_out8459_out1;

  Logical_Operator_out9228_out1 <= Logical_Operator_out8204_out1 XOR Logical_Operator_out8460_out1;

  Logical_Operator_out9229_out1 <= Logical_Operator_out8205_out1 XOR Logical_Operator_out8461_out1;

  Logical_Operator_out9230_out1 <= Logical_Operator_out8206_out1 XOR Logical_Operator_out8462_out1;

  Logical_Operator_out9231_out1 <= Logical_Operator_out8207_out1 XOR Logical_Operator_out8463_out1;

  Logical_Operator_out9232_out1 <= Logical_Operator_out8208_out1 XOR Logical_Operator_out8464_out1;

  Logical_Operator_out9233_out1 <= Logical_Operator_out8209_out1 XOR Logical_Operator_out8465_out1;

  Logical_Operator_out9234_out1 <= Logical_Operator_out8210_out1 XOR Logical_Operator_out8466_out1;

  Logical_Operator_out9235_out1 <= Logical_Operator_out8211_out1 XOR Logical_Operator_out8467_out1;

  Logical_Operator_out9236_out1 <= Logical_Operator_out8212_out1 XOR Logical_Operator_out8468_out1;

  Logical_Operator_out9237_out1 <= Logical_Operator_out8213_out1 XOR Logical_Operator_out8469_out1;

  Logical_Operator_out9238_out1 <= Logical_Operator_out8214_out1 XOR Logical_Operator_out8470_out1;

  Logical_Operator_out9239_out1 <= Logical_Operator_out8215_out1 XOR Logical_Operator_out8471_out1;

  Logical_Operator_out9240_out1 <= Logical_Operator_out8216_out1 XOR Logical_Operator_out8472_out1;

  Logical_Operator_out9241_out1 <= Logical_Operator_out8217_out1 XOR Logical_Operator_out8473_out1;

  Logical_Operator_out9242_out1 <= Logical_Operator_out8218_out1 XOR Logical_Operator_out8474_out1;

  Logical_Operator_out9243_out1 <= Logical_Operator_out8219_out1 XOR Logical_Operator_out8475_out1;

  Logical_Operator_out9244_out1 <= Logical_Operator_out8220_out1 XOR Logical_Operator_out8476_out1;

  Logical_Operator_out9245_out1 <= Logical_Operator_out8221_out1 XOR Logical_Operator_out8477_out1;

  Logical_Operator_out9246_out1 <= Logical_Operator_out8222_out1 XOR Logical_Operator_out8478_out1;

  Logical_Operator_out9247_out1 <= Logical_Operator_out8223_out1 XOR Logical_Operator_out8479_out1;

  Logical_Operator_out9248_out1 <= Logical_Operator_out8224_out1 XOR Logical_Operator_out8480_out1;

  Logical_Operator_out9249_out1 <= Logical_Operator_out8225_out1 XOR Logical_Operator_out8481_out1;

  Logical_Operator_out9250_out1 <= Logical_Operator_out8226_out1 XOR Logical_Operator_out8482_out1;

  Logical_Operator_out9251_out1 <= Logical_Operator_out8227_out1 XOR Logical_Operator_out8483_out1;

  Logical_Operator_out9252_out1 <= Logical_Operator_out8228_out1 XOR Logical_Operator_out8484_out1;

  Logical_Operator_out9253_out1 <= Logical_Operator_out8229_out1 XOR Logical_Operator_out8485_out1;

  Logical_Operator_out9254_out1 <= Logical_Operator_out8230_out1 XOR Logical_Operator_out8486_out1;

  Logical_Operator_out9255_out1 <= Logical_Operator_out8231_out1 XOR Logical_Operator_out8487_out1;

  Logical_Operator_out9256_out1 <= Logical_Operator_out8232_out1 XOR Logical_Operator_out8488_out1;

  Logical_Operator_out9257_out1 <= Logical_Operator_out8233_out1 XOR Logical_Operator_out8489_out1;

  Logical_Operator_out9258_out1 <= Logical_Operator_out8234_out1 XOR Logical_Operator_out8490_out1;

  Logical_Operator_out9259_out1 <= Logical_Operator_out8235_out1 XOR Logical_Operator_out8491_out1;

  Logical_Operator_out9260_out1 <= Logical_Operator_out8236_out1 XOR Logical_Operator_out8492_out1;

  Logical_Operator_out9261_out1 <= Logical_Operator_out8237_out1 XOR Logical_Operator_out8493_out1;

  Logical_Operator_out9262_out1 <= Logical_Operator_out8238_out1 XOR Logical_Operator_out8494_out1;

  Logical_Operator_out9263_out1 <= Logical_Operator_out8239_out1 XOR Logical_Operator_out8495_out1;

  Logical_Operator_out9264_out1 <= Logical_Operator_out8240_out1 XOR Logical_Operator_out8496_out1;

  Logical_Operator_out9265_out1 <= Logical_Operator_out8241_out1 XOR Logical_Operator_out8497_out1;

  Logical_Operator_out9266_out1 <= Logical_Operator_out8242_out1 XOR Logical_Operator_out8498_out1;

  Logical_Operator_out9267_out1 <= Logical_Operator_out8243_out1 XOR Logical_Operator_out8499_out1;

  Logical_Operator_out9268_out1 <= Logical_Operator_out8244_out1 XOR Logical_Operator_out8500_out1;

  Logical_Operator_out9269_out1 <= Logical_Operator_out8245_out1 XOR Logical_Operator_out8501_out1;

  Logical_Operator_out9270_out1 <= Logical_Operator_out8246_out1 XOR Logical_Operator_out8502_out1;

  Logical_Operator_out9271_out1 <= Logical_Operator_out8247_out1 XOR Logical_Operator_out8503_out1;

  Logical_Operator_out9272_out1 <= Logical_Operator_out8248_out1 XOR Logical_Operator_out8504_out1;

  Logical_Operator_out9273_out1 <= Logical_Operator_out8249_out1 XOR Logical_Operator_out8505_out1;

  Logical_Operator_out9274_out1 <= Logical_Operator_out8250_out1 XOR Logical_Operator_out8506_out1;

  Logical_Operator_out9275_out1 <= Logical_Operator_out8251_out1 XOR Logical_Operator_out8507_out1;

  Logical_Operator_out9276_out1 <= Logical_Operator_out8252_out1 XOR Logical_Operator_out8508_out1;

  Logical_Operator_out9277_out1 <= Logical_Operator_out8253_out1 XOR Logical_Operator_out8509_out1;

  Logical_Operator_out9278_out1 <= Logical_Operator_out8254_out1 XOR Logical_Operator_out8510_out1;

  Logical_Operator_out9279_out1 <= Logical_Operator_out8255_out1 XOR Logical_Operator_out8511_out1;

  Logical_Operator_out9280_out1 <= Logical_Operator_out8256_out1 XOR Logical_Operator_out8512_out1;

  Logical_Operator_out9281_out1 <= Logical_Operator_out8257_out1 XOR Logical_Operator_out8513_out1;

  Logical_Operator_out9282_out1 <= Logical_Operator_out8258_out1 XOR Logical_Operator_out8514_out1;

  Logical_Operator_out9283_out1 <= Logical_Operator_out8259_out1 XOR Logical_Operator_out8515_out1;

  Logical_Operator_out9284_out1 <= Logical_Operator_out8260_out1 XOR Logical_Operator_out8516_out1;

  Logical_Operator_out9285_out1 <= Logical_Operator_out8261_out1 XOR Logical_Operator_out8517_out1;

  Logical_Operator_out9286_out1 <= Logical_Operator_out8262_out1 XOR Logical_Operator_out8518_out1;

  Logical_Operator_out9287_out1 <= Logical_Operator_out8263_out1 XOR Logical_Operator_out8519_out1;

  Logical_Operator_out9288_out1 <= Logical_Operator_out8264_out1 XOR Logical_Operator_out8520_out1;

  Logical_Operator_out9289_out1 <= Logical_Operator_out8265_out1 XOR Logical_Operator_out8521_out1;

  Logical_Operator_out9290_out1 <= Logical_Operator_out8266_out1 XOR Logical_Operator_out8522_out1;

  Logical_Operator_out9291_out1 <= Logical_Operator_out8267_out1 XOR Logical_Operator_out8523_out1;

  Logical_Operator_out9292_out1 <= Logical_Operator_out8268_out1 XOR Logical_Operator_out8524_out1;

  Logical_Operator_out9293_out1 <= Logical_Operator_out8269_out1 XOR Logical_Operator_out8525_out1;

  Logical_Operator_out9294_out1 <= Logical_Operator_out8270_out1 XOR Logical_Operator_out8526_out1;

  Logical_Operator_out9295_out1 <= Logical_Operator_out8271_out1 XOR Logical_Operator_out8527_out1;

  Logical_Operator_out9296_out1 <= Logical_Operator_out8272_out1 XOR Logical_Operator_out8528_out1;

  Logical_Operator_out9297_out1 <= Logical_Operator_out8273_out1 XOR Logical_Operator_out8529_out1;

  Logical_Operator_out9298_out1 <= Logical_Operator_out8274_out1 XOR Logical_Operator_out8530_out1;

  Logical_Operator_out9299_out1 <= Logical_Operator_out8275_out1 XOR Logical_Operator_out8531_out1;

  Logical_Operator_out9300_out1 <= Logical_Operator_out8276_out1 XOR Logical_Operator_out8532_out1;

  Logical_Operator_out9301_out1 <= Logical_Operator_out8277_out1 XOR Logical_Operator_out8533_out1;

  Logical_Operator_out9302_out1 <= Logical_Operator_out8278_out1 XOR Logical_Operator_out8534_out1;

  Logical_Operator_out9303_out1 <= Logical_Operator_out8279_out1 XOR Logical_Operator_out8535_out1;

  Logical_Operator_out9304_out1 <= Logical_Operator_out8280_out1 XOR Logical_Operator_out8536_out1;

  Logical_Operator_out9305_out1 <= Logical_Operator_out8281_out1 XOR Logical_Operator_out8537_out1;

  Logical_Operator_out9306_out1 <= Logical_Operator_out8282_out1 XOR Logical_Operator_out8538_out1;

  Logical_Operator_out9307_out1 <= Logical_Operator_out8283_out1 XOR Logical_Operator_out8539_out1;

  Logical_Operator_out9308_out1 <= Logical_Operator_out8284_out1 XOR Logical_Operator_out8540_out1;

  Logical_Operator_out9309_out1 <= Logical_Operator_out8285_out1 XOR Logical_Operator_out8541_out1;

  Logical_Operator_out9310_out1 <= Logical_Operator_out8286_out1 XOR Logical_Operator_out8542_out1;

  Logical_Operator_out9311_out1 <= Logical_Operator_out8287_out1 XOR Logical_Operator_out8543_out1;

  Logical_Operator_out9312_out1 <= Logical_Operator_out8288_out1 XOR Logical_Operator_out8544_out1;

  Logical_Operator_out9313_out1 <= Logical_Operator_out8289_out1 XOR Logical_Operator_out8545_out1;

  Logical_Operator_out9314_out1 <= Logical_Operator_out8290_out1 XOR Logical_Operator_out8546_out1;

  Logical_Operator_out9315_out1 <= Logical_Operator_out8291_out1 XOR Logical_Operator_out8547_out1;

  Logical_Operator_out9316_out1 <= Logical_Operator_out8292_out1 XOR Logical_Operator_out8548_out1;

  Logical_Operator_out9317_out1 <= Logical_Operator_out8293_out1 XOR Logical_Operator_out8549_out1;

  Logical_Operator_out9318_out1 <= Logical_Operator_out8294_out1 XOR Logical_Operator_out8550_out1;

  Logical_Operator_out9319_out1 <= Logical_Operator_out8295_out1 XOR Logical_Operator_out8551_out1;

  Logical_Operator_out9320_out1 <= Logical_Operator_out8296_out1 XOR Logical_Operator_out8552_out1;

  Logical_Operator_out9321_out1 <= Logical_Operator_out8297_out1 XOR Logical_Operator_out8553_out1;

  Logical_Operator_out9322_out1 <= Logical_Operator_out8298_out1 XOR Logical_Operator_out8554_out1;

  Logical_Operator_out9323_out1 <= Logical_Operator_out8299_out1 XOR Logical_Operator_out8555_out1;

  Logical_Operator_out9324_out1 <= Logical_Operator_out8300_out1 XOR Logical_Operator_out8556_out1;

  Logical_Operator_out9325_out1 <= Logical_Operator_out8301_out1 XOR Logical_Operator_out8557_out1;

  Logical_Operator_out9326_out1 <= Logical_Operator_out8302_out1 XOR Logical_Operator_out8558_out1;

  Logical_Operator_out9327_out1 <= Logical_Operator_out8303_out1 XOR Logical_Operator_out8559_out1;

  Logical_Operator_out9328_out1 <= Logical_Operator_out8304_out1 XOR Logical_Operator_out8560_out1;

  Logical_Operator_out9329_out1 <= Logical_Operator_out8305_out1 XOR Logical_Operator_out8561_out1;

  Logical_Operator_out9330_out1 <= Logical_Operator_out8306_out1 XOR Logical_Operator_out8562_out1;

  Logical_Operator_out9331_out1 <= Logical_Operator_out8307_out1 XOR Logical_Operator_out8563_out1;

  Logical_Operator_out9332_out1 <= Logical_Operator_out8308_out1 XOR Logical_Operator_out8564_out1;

  Logical_Operator_out9333_out1 <= Logical_Operator_out8309_out1 XOR Logical_Operator_out8565_out1;

  Logical_Operator_out9334_out1 <= Logical_Operator_out8310_out1 XOR Logical_Operator_out8566_out1;

  Logical_Operator_out9335_out1 <= Logical_Operator_out8311_out1 XOR Logical_Operator_out8567_out1;

  Logical_Operator_out9336_out1 <= Logical_Operator_out8312_out1 XOR Logical_Operator_out8568_out1;

  Logical_Operator_out9337_out1 <= Logical_Operator_out8313_out1 XOR Logical_Operator_out8569_out1;

  Logical_Operator_out9338_out1 <= Logical_Operator_out8314_out1 XOR Logical_Operator_out8570_out1;

  Logical_Operator_out9339_out1 <= Logical_Operator_out8315_out1 XOR Logical_Operator_out8571_out1;

  Logical_Operator_out9340_out1 <= Logical_Operator_out8316_out1 XOR Logical_Operator_out8572_out1;

  Logical_Operator_out9341_out1 <= Logical_Operator_out8317_out1 XOR Logical_Operator_out8573_out1;

  Logical_Operator_out9342_out1 <= Logical_Operator_out8318_out1 XOR Logical_Operator_out8574_out1;

  Logical_Operator_out9343_out1 <= Logical_Operator_out8319_out1 XOR Logical_Operator_out8575_out1;

  Logical_Operator_out9344_out1 <= Logical_Operator_out8320_out1 XOR Logical_Operator_out8576_out1;

  Logical_Operator_out9345_out1 <= Logical_Operator_out8321_out1 XOR Logical_Operator_out8577_out1;

  Logical_Operator_out9346_out1 <= Logical_Operator_out8322_out1 XOR Logical_Operator_out8578_out1;

  Logical_Operator_out9347_out1 <= Logical_Operator_out8323_out1 XOR Logical_Operator_out8579_out1;

  Logical_Operator_out9348_out1 <= Logical_Operator_out8324_out1 XOR Logical_Operator_out8580_out1;

  Logical_Operator_out9349_out1 <= Logical_Operator_out8325_out1 XOR Logical_Operator_out8581_out1;

  Logical_Operator_out9350_out1 <= Logical_Operator_out8326_out1 XOR Logical_Operator_out8582_out1;

  Logical_Operator_out9351_out1 <= Logical_Operator_out8327_out1 XOR Logical_Operator_out8583_out1;

  Logical_Operator_out9352_out1 <= Logical_Operator_out8328_out1 XOR Logical_Operator_out8584_out1;

  Logical_Operator_out9353_out1 <= Logical_Operator_out8329_out1 XOR Logical_Operator_out8585_out1;

  Logical_Operator_out9354_out1 <= Logical_Operator_out8330_out1 XOR Logical_Operator_out8586_out1;

  Logical_Operator_out9355_out1 <= Logical_Operator_out8331_out1 XOR Logical_Operator_out8587_out1;

  Logical_Operator_out9356_out1 <= Logical_Operator_out8332_out1 XOR Logical_Operator_out8588_out1;

  Logical_Operator_out9357_out1 <= Logical_Operator_out8333_out1 XOR Logical_Operator_out8589_out1;

  Logical_Operator_out9358_out1 <= Logical_Operator_out8334_out1 XOR Logical_Operator_out8590_out1;

  Logical_Operator_out9359_out1 <= Logical_Operator_out8335_out1 XOR Logical_Operator_out8591_out1;

  Logical_Operator_out9360_out1 <= Logical_Operator_out8336_out1 XOR Logical_Operator_out8592_out1;

  Logical_Operator_out9361_out1 <= Logical_Operator_out8337_out1 XOR Logical_Operator_out8593_out1;

  Logical_Operator_out9362_out1 <= Logical_Operator_out8338_out1 XOR Logical_Operator_out8594_out1;

  Logical_Operator_out9363_out1 <= Logical_Operator_out8339_out1 XOR Logical_Operator_out8595_out1;

  Logical_Operator_out9364_out1 <= Logical_Operator_out8340_out1 XOR Logical_Operator_out8596_out1;

  Logical_Operator_out9365_out1 <= Logical_Operator_out8341_out1 XOR Logical_Operator_out8597_out1;

  Logical_Operator_out9366_out1 <= Logical_Operator_out8342_out1 XOR Logical_Operator_out8598_out1;

  Logical_Operator_out9367_out1 <= Logical_Operator_out8343_out1 XOR Logical_Operator_out8599_out1;

  Logical_Operator_out9368_out1 <= Logical_Operator_out8344_out1 XOR Logical_Operator_out8600_out1;

  Logical_Operator_out9369_out1 <= Logical_Operator_out8345_out1 XOR Logical_Operator_out8601_out1;

  Logical_Operator_out9370_out1 <= Logical_Operator_out8346_out1 XOR Logical_Operator_out8602_out1;

  Logical_Operator_out9371_out1 <= Logical_Operator_out8347_out1 XOR Logical_Operator_out8603_out1;

  Logical_Operator_out9372_out1 <= Logical_Operator_out8348_out1 XOR Logical_Operator_out8604_out1;

  Logical_Operator_out9373_out1 <= Logical_Operator_out8349_out1 XOR Logical_Operator_out8605_out1;

  Logical_Operator_out9374_out1 <= Logical_Operator_out8350_out1 XOR Logical_Operator_out8606_out1;

  Logical_Operator_out9375_out1 <= Logical_Operator_out8351_out1 XOR Logical_Operator_out8607_out1;

  Logical_Operator_out9376_out1 <= Logical_Operator_out8352_out1 XOR Logical_Operator_out8608_out1;

  Logical_Operator_out9377_out1 <= Logical_Operator_out8353_out1 XOR Logical_Operator_out8609_out1;

  Logical_Operator_out9378_out1 <= Logical_Operator_out8354_out1 XOR Logical_Operator_out8610_out1;

  Logical_Operator_out9379_out1 <= Logical_Operator_out8355_out1 XOR Logical_Operator_out8611_out1;

  Logical_Operator_out9380_out1 <= Logical_Operator_out8356_out1 XOR Logical_Operator_out8612_out1;

  Logical_Operator_out9381_out1 <= Logical_Operator_out8357_out1 XOR Logical_Operator_out8613_out1;

  Logical_Operator_out9382_out1 <= Logical_Operator_out8358_out1 XOR Logical_Operator_out8614_out1;

  Logical_Operator_out9383_out1 <= Logical_Operator_out8359_out1 XOR Logical_Operator_out8615_out1;

  Logical_Operator_out9384_out1 <= Logical_Operator_out8360_out1 XOR Logical_Operator_out8616_out1;

  Logical_Operator_out9385_out1 <= Logical_Operator_out8361_out1 XOR Logical_Operator_out8617_out1;

  Logical_Operator_out9386_out1 <= Logical_Operator_out8362_out1 XOR Logical_Operator_out8618_out1;

  Logical_Operator_out9387_out1 <= Logical_Operator_out8363_out1 XOR Logical_Operator_out8619_out1;

  Logical_Operator_out9388_out1 <= Logical_Operator_out8364_out1 XOR Logical_Operator_out8620_out1;

  Logical_Operator_out9389_out1 <= Logical_Operator_out8365_out1 XOR Logical_Operator_out8621_out1;

  Logical_Operator_out9390_out1 <= Logical_Operator_out8366_out1 XOR Logical_Operator_out8622_out1;

  Logical_Operator_out9391_out1 <= Logical_Operator_out8367_out1 XOR Logical_Operator_out8623_out1;

  Logical_Operator_out9392_out1 <= Logical_Operator_out8368_out1 XOR Logical_Operator_out8624_out1;

  Logical_Operator_out9393_out1 <= Logical_Operator_out8369_out1 XOR Logical_Operator_out8625_out1;

  Logical_Operator_out9394_out1 <= Logical_Operator_out8370_out1 XOR Logical_Operator_out8626_out1;

  Logical_Operator_out9395_out1 <= Logical_Operator_out8371_out1 XOR Logical_Operator_out8627_out1;

  Logical_Operator_out9396_out1 <= Logical_Operator_out8372_out1 XOR Logical_Operator_out8628_out1;

  Logical_Operator_out9397_out1 <= Logical_Operator_out8373_out1 XOR Logical_Operator_out8629_out1;

  Logical_Operator_out9398_out1 <= Logical_Operator_out8374_out1 XOR Logical_Operator_out8630_out1;

  Logical_Operator_out9399_out1 <= Logical_Operator_out8375_out1 XOR Logical_Operator_out8631_out1;

  Logical_Operator_out9400_out1 <= Logical_Operator_out8376_out1 XOR Logical_Operator_out8632_out1;

  Logical_Operator_out9401_out1 <= Logical_Operator_out8377_out1 XOR Logical_Operator_out8633_out1;

  Logical_Operator_out9402_out1 <= Logical_Operator_out8378_out1 XOR Logical_Operator_out8634_out1;

  Logical_Operator_out9403_out1 <= Logical_Operator_out8379_out1 XOR Logical_Operator_out8635_out1;

  Logical_Operator_out9404_out1 <= Logical_Operator_out8380_out1 XOR Logical_Operator_out8636_out1;

  Logical_Operator_out9405_out1 <= Logical_Operator_out8381_out1 XOR Logical_Operator_out8637_out1;

  Logical_Operator_out9406_out1 <= Logical_Operator_out8382_out1 XOR Logical_Operator_out8638_out1;

  Logical_Operator_out9407_out1 <= Logical_Operator_out8383_out1 XOR Logical_Operator_out8639_out1;

  Logical_Operator_out9408_out1 <= Logical_Operator_out8384_out1 XOR Logical_Operator_out8640_out1;

  Logical_Operator_out9409_out1 <= Logical_Operator_out8385_out1 XOR Logical_Operator_out8641_out1;

  Logical_Operator_out9410_out1 <= Logical_Operator_out8386_out1 XOR Logical_Operator_out8642_out1;

  Logical_Operator_out9411_out1 <= Logical_Operator_out8387_out1 XOR Logical_Operator_out8643_out1;

  Logical_Operator_out9412_out1 <= Logical_Operator_out8388_out1 XOR Logical_Operator_out8644_out1;

  Logical_Operator_out9413_out1 <= Logical_Operator_out8389_out1 XOR Logical_Operator_out8645_out1;

  Logical_Operator_out9414_out1 <= Logical_Operator_out8390_out1 XOR Logical_Operator_out8646_out1;

  Logical_Operator_out9415_out1 <= Logical_Operator_out8391_out1 XOR Logical_Operator_out8647_out1;

  Logical_Operator_out9416_out1 <= Logical_Operator_out8392_out1 XOR Logical_Operator_out8648_out1;

  Logical_Operator_out9417_out1 <= Logical_Operator_out8393_out1 XOR Logical_Operator_out8649_out1;

  Logical_Operator_out9418_out1 <= Logical_Operator_out8394_out1 XOR Logical_Operator_out8650_out1;

  Logical_Operator_out9419_out1 <= Logical_Operator_out8395_out1 XOR Logical_Operator_out8651_out1;

  Logical_Operator_out9420_out1 <= Logical_Operator_out8396_out1 XOR Logical_Operator_out8652_out1;

  Logical_Operator_out9421_out1 <= Logical_Operator_out8397_out1 XOR Logical_Operator_out8653_out1;

  Logical_Operator_out9422_out1 <= Logical_Operator_out8398_out1 XOR Logical_Operator_out8654_out1;

  Logical_Operator_out9423_out1 <= Logical_Operator_out8399_out1 XOR Logical_Operator_out8655_out1;

  Logical_Operator_out9424_out1 <= Logical_Operator_out8400_out1 XOR Logical_Operator_out8656_out1;

  Logical_Operator_out9425_out1 <= Logical_Operator_out8401_out1 XOR Logical_Operator_out8657_out1;

  Logical_Operator_out9426_out1 <= Logical_Operator_out8402_out1 XOR Logical_Operator_out8658_out1;

  Logical_Operator_out9427_out1 <= Logical_Operator_out8403_out1 XOR Logical_Operator_out8659_out1;

  Logical_Operator_out9428_out1 <= Logical_Operator_out8404_out1 XOR Logical_Operator_out8660_out1;

  Logical_Operator_out9429_out1 <= Logical_Operator_out8405_out1 XOR Logical_Operator_out8661_out1;

  Logical_Operator_out9430_out1 <= Logical_Operator_out8406_out1 XOR Logical_Operator_out8662_out1;

  Logical_Operator_out9431_out1 <= Logical_Operator_out8407_out1 XOR Logical_Operator_out8663_out1;

  Logical_Operator_out9432_out1 <= Logical_Operator_out8408_out1 XOR Logical_Operator_out8664_out1;

  Logical_Operator_out9433_out1 <= Logical_Operator_out8409_out1 XOR Logical_Operator_out8665_out1;

  Logical_Operator_out9434_out1 <= Logical_Operator_out8410_out1 XOR Logical_Operator_out8666_out1;

  Logical_Operator_out9435_out1 <= Logical_Operator_out8411_out1 XOR Logical_Operator_out8667_out1;

  Logical_Operator_out9436_out1 <= Logical_Operator_out8412_out1 XOR Logical_Operator_out8668_out1;

  Logical_Operator_out9437_out1 <= Logical_Operator_out8413_out1 XOR Logical_Operator_out8669_out1;

  Logical_Operator_out9438_out1 <= Logical_Operator_out8414_out1 XOR Logical_Operator_out8670_out1;

  Logical_Operator_out9439_out1 <= Logical_Operator_out8415_out1 XOR Logical_Operator_out8671_out1;

  Logical_Operator_out9440_out1 <= Logical_Operator_out8416_out1 XOR Logical_Operator_out8672_out1;

  Logical_Operator_out9441_out1 <= Logical_Operator_out8417_out1 XOR Logical_Operator_out8673_out1;

  Logical_Operator_out9442_out1 <= Logical_Operator_out8418_out1 XOR Logical_Operator_out8674_out1;

  Logical_Operator_out9443_out1 <= Logical_Operator_out8419_out1 XOR Logical_Operator_out8675_out1;

  Logical_Operator_out9444_out1 <= Logical_Operator_out8420_out1 XOR Logical_Operator_out8676_out1;

  Logical_Operator_out9445_out1 <= Logical_Operator_out8421_out1 XOR Logical_Operator_out8677_out1;

  Logical_Operator_out9446_out1 <= Logical_Operator_out8422_out1 XOR Logical_Operator_out8678_out1;

  Logical_Operator_out9447_out1 <= Logical_Operator_out8423_out1 XOR Logical_Operator_out8679_out1;

  Logical_Operator_out9448_out1 <= Logical_Operator_out8424_out1 XOR Logical_Operator_out8680_out1;

  Logical_Operator_out9449_out1 <= Logical_Operator_out8425_out1 XOR Logical_Operator_out8681_out1;

  Logical_Operator_out9450_out1 <= Logical_Operator_out8426_out1 XOR Logical_Operator_out8682_out1;

  Logical_Operator_out9451_out1 <= Logical_Operator_out8427_out1 XOR Logical_Operator_out8683_out1;

  Logical_Operator_out9452_out1 <= Logical_Operator_out8428_out1 XOR Logical_Operator_out8684_out1;

  Logical_Operator_out9453_out1 <= Logical_Operator_out8429_out1 XOR Logical_Operator_out8685_out1;

  Logical_Operator_out9454_out1 <= Logical_Operator_out8430_out1 XOR Logical_Operator_out8686_out1;

  Logical_Operator_out9455_out1 <= Logical_Operator_out8431_out1 XOR Logical_Operator_out8687_out1;

  Logical_Operator_out9456_out1 <= Logical_Operator_out8432_out1 XOR Logical_Operator_out8688_out1;

  Logical_Operator_out9457_out1 <= Logical_Operator_out8433_out1 XOR Logical_Operator_out8689_out1;

  Logical_Operator_out9458_out1 <= Logical_Operator_out8434_out1 XOR Logical_Operator_out8690_out1;

  Logical_Operator_out9459_out1 <= Logical_Operator_out8435_out1 XOR Logical_Operator_out8691_out1;

  Logical_Operator_out9460_out1 <= Logical_Operator_out8436_out1 XOR Logical_Operator_out8692_out1;

  Logical_Operator_out9461_out1 <= Logical_Operator_out8437_out1 XOR Logical_Operator_out8693_out1;

  Logical_Operator_out9462_out1 <= Logical_Operator_out8438_out1 XOR Logical_Operator_out8694_out1;

  Logical_Operator_out9463_out1 <= Logical_Operator_out8439_out1 XOR Logical_Operator_out8695_out1;

  Logical_Operator_out9464_out1 <= Logical_Operator_out8440_out1 XOR Logical_Operator_out8696_out1;

  Logical_Operator_out9465_out1 <= Logical_Operator_out8441_out1 XOR Logical_Operator_out8697_out1;

  Logical_Operator_out9466_out1 <= Logical_Operator_out8442_out1 XOR Logical_Operator_out8698_out1;

  Logical_Operator_out9467_out1 <= Logical_Operator_out8443_out1 XOR Logical_Operator_out8699_out1;

  Logical_Operator_out9468_out1 <= Logical_Operator_out8444_out1 XOR Logical_Operator_out8700_out1;

  Logical_Operator_out9469_out1 <= Logical_Operator_out8445_out1 XOR Logical_Operator_out8701_out1;

  Logical_Operator_out9470_out1 <= Logical_Operator_out8446_out1 XOR Logical_Operator_out8702_out1;

  Logical_Operator_out9471_out1 <= Logical_Operator_out8447_out1 XOR Logical_Operator_out8703_out1;

  Logical_Operator_out9472_out1 <= Logical_Operator_out8448_out1 XOR Logical_Operator_out8704_out1;

  Logical_Operator_out9473_out1 <= Logical_Operator_out7297_out1 XOR Logical_Operator_out7553_out1;

  Logical_Operator_out9474_out1 <= Logical_Operator_out7298_out1 XOR Logical_Operator_out7554_out1;

  Logical_Operator_out9475_out1 <= Logical_Operator_out7299_out1 XOR Logical_Operator_out7555_out1;

  Logical_Operator_out9476_out1 <= Logical_Operator_out7300_out1 XOR Logical_Operator_out7556_out1;

  Logical_Operator_out9477_out1 <= Logical_Operator_out7301_out1 XOR Logical_Operator_out7557_out1;

  Logical_Operator_out9478_out1 <= Logical_Operator_out7302_out1 XOR Logical_Operator_out7558_out1;

  Logical_Operator_out9479_out1 <= Logical_Operator_out7303_out1 XOR Logical_Operator_out7559_out1;

  Logical_Operator_out9480_out1 <= Logical_Operator_out7304_out1 XOR Logical_Operator_out7560_out1;

  Logical_Operator_out9481_out1 <= Logical_Operator_out7305_out1 XOR Logical_Operator_out7561_out1;

  Logical_Operator_out9482_out1 <= Logical_Operator_out7306_out1 XOR Logical_Operator_out7562_out1;

  Logical_Operator_out9483_out1 <= Logical_Operator_out7307_out1 XOR Logical_Operator_out7563_out1;

  Logical_Operator_out9484_out1 <= Logical_Operator_out7308_out1 XOR Logical_Operator_out7564_out1;

  Logical_Operator_out9485_out1 <= Logical_Operator_out7309_out1 XOR Logical_Operator_out7565_out1;

  Logical_Operator_out9486_out1 <= Logical_Operator_out7310_out1 XOR Logical_Operator_out7566_out1;

  Logical_Operator_out9487_out1 <= Logical_Operator_out7311_out1 XOR Logical_Operator_out7567_out1;

  Logical_Operator_out9488_out1 <= Logical_Operator_out7312_out1 XOR Logical_Operator_out7568_out1;

  Logical_Operator_out9489_out1 <= Logical_Operator_out7313_out1 XOR Logical_Operator_out7569_out1;

  Logical_Operator_out9490_out1 <= Logical_Operator_out7314_out1 XOR Logical_Operator_out7570_out1;

  Logical_Operator_out9491_out1 <= Logical_Operator_out7315_out1 XOR Logical_Operator_out7571_out1;

  Logical_Operator_out9492_out1 <= Logical_Operator_out7316_out1 XOR Logical_Operator_out7572_out1;

  Logical_Operator_out9493_out1 <= Logical_Operator_out7317_out1 XOR Logical_Operator_out7573_out1;

  Logical_Operator_out9494_out1 <= Logical_Operator_out7318_out1 XOR Logical_Operator_out7574_out1;

  Logical_Operator_out9495_out1 <= Logical_Operator_out7319_out1 XOR Logical_Operator_out7575_out1;

  Logical_Operator_out9496_out1 <= Logical_Operator_out7320_out1 XOR Logical_Operator_out7576_out1;

  Logical_Operator_out9497_out1 <= Logical_Operator_out7321_out1 XOR Logical_Operator_out7577_out1;

  Logical_Operator_out9498_out1 <= Logical_Operator_out7322_out1 XOR Logical_Operator_out7578_out1;

  Logical_Operator_out9499_out1 <= Logical_Operator_out7323_out1 XOR Logical_Operator_out7579_out1;

  Logical_Operator_out9500_out1 <= Logical_Operator_out7324_out1 XOR Logical_Operator_out7580_out1;

  Logical_Operator_out9501_out1 <= Logical_Operator_out7325_out1 XOR Logical_Operator_out7581_out1;

  Logical_Operator_out9502_out1 <= Logical_Operator_out7326_out1 XOR Logical_Operator_out7582_out1;

  Logical_Operator_out9503_out1 <= Logical_Operator_out7327_out1 XOR Logical_Operator_out7583_out1;

  Logical_Operator_out9504_out1 <= Logical_Operator_out7328_out1 XOR Logical_Operator_out7584_out1;

  Logical_Operator_out9505_out1 <= Logical_Operator_out7329_out1 XOR Logical_Operator_out7585_out1;

  Logical_Operator_out9506_out1 <= Logical_Operator_out7330_out1 XOR Logical_Operator_out7586_out1;

  Logical_Operator_out9507_out1 <= Logical_Operator_out7331_out1 XOR Logical_Operator_out7587_out1;

  Logical_Operator_out9508_out1 <= Logical_Operator_out7332_out1 XOR Logical_Operator_out7588_out1;

  Logical_Operator_out9509_out1 <= Logical_Operator_out7333_out1 XOR Logical_Operator_out7589_out1;

  Logical_Operator_out9510_out1 <= Logical_Operator_out7334_out1 XOR Logical_Operator_out7590_out1;

  Logical_Operator_out9511_out1 <= Logical_Operator_out7335_out1 XOR Logical_Operator_out7591_out1;

  Logical_Operator_out9512_out1 <= Logical_Operator_out7336_out1 XOR Logical_Operator_out7592_out1;

  Logical_Operator_out9513_out1 <= Logical_Operator_out7337_out1 XOR Logical_Operator_out7593_out1;

  Logical_Operator_out9514_out1 <= Logical_Operator_out7338_out1 XOR Logical_Operator_out7594_out1;

  Logical_Operator_out9515_out1 <= Logical_Operator_out7339_out1 XOR Logical_Operator_out7595_out1;

  Logical_Operator_out9516_out1 <= Logical_Operator_out7340_out1 XOR Logical_Operator_out7596_out1;

  Logical_Operator_out9517_out1 <= Logical_Operator_out7341_out1 XOR Logical_Operator_out7597_out1;

  Logical_Operator_out9518_out1 <= Logical_Operator_out7342_out1 XOR Logical_Operator_out7598_out1;

  Logical_Operator_out9519_out1 <= Logical_Operator_out7343_out1 XOR Logical_Operator_out7599_out1;

  Logical_Operator_out9520_out1 <= Logical_Operator_out7344_out1 XOR Logical_Operator_out7600_out1;

  Logical_Operator_out9521_out1 <= Logical_Operator_out7345_out1 XOR Logical_Operator_out7601_out1;

  Logical_Operator_out9522_out1 <= Logical_Operator_out7346_out1 XOR Logical_Operator_out7602_out1;

  Logical_Operator_out9523_out1 <= Logical_Operator_out7347_out1 XOR Logical_Operator_out7603_out1;

  Logical_Operator_out9524_out1 <= Logical_Operator_out7348_out1 XOR Logical_Operator_out7604_out1;

  Logical_Operator_out9525_out1 <= Logical_Operator_out7349_out1 XOR Logical_Operator_out7605_out1;

  Logical_Operator_out9526_out1 <= Logical_Operator_out7350_out1 XOR Logical_Operator_out7606_out1;

  Logical_Operator_out9527_out1 <= Logical_Operator_out7351_out1 XOR Logical_Operator_out7607_out1;

  Logical_Operator_out9528_out1 <= Logical_Operator_out7352_out1 XOR Logical_Operator_out7608_out1;

  Logical_Operator_out9529_out1 <= Logical_Operator_out7353_out1 XOR Logical_Operator_out7609_out1;

  Logical_Operator_out9530_out1 <= Logical_Operator_out7354_out1 XOR Logical_Operator_out7610_out1;

  Logical_Operator_out9531_out1 <= Logical_Operator_out7355_out1 XOR Logical_Operator_out7611_out1;

  Logical_Operator_out9532_out1 <= Logical_Operator_out7356_out1 XOR Logical_Operator_out7612_out1;

  Logical_Operator_out9533_out1 <= Logical_Operator_out7357_out1 XOR Logical_Operator_out7613_out1;

  Logical_Operator_out9534_out1 <= Logical_Operator_out7358_out1 XOR Logical_Operator_out7614_out1;

  Logical_Operator_out9535_out1 <= Logical_Operator_out7359_out1 XOR Logical_Operator_out7615_out1;

  Logical_Operator_out9536_out1 <= Logical_Operator_out7360_out1 XOR Logical_Operator_out7616_out1;

  Logical_Operator_out9537_out1 <= Logical_Operator_out7361_out1 XOR Logical_Operator_out7617_out1;

  Logical_Operator_out9538_out1 <= Logical_Operator_out7362_out1 XOR Logical_Operator_out7618_out1;

  Logical_Operator_out9539_out1 <= Logical_Operator_out7363_out1 XOR Logical_Operator_out7619_out1;

  Logical_Operator_out9540_out1 <= Logical_Operator_out7364_out1 XOR Logical_Operator_out7620_out1;

  Logical_Operator_out9541_out1 <= Logical_Operator_out7365_out1 XOR Logical_Operator_out7621_out1;

  Logical_Operator_out9542_out1 <= Logical_Operator_out7366_out1 XOR Logical_Operator_out7622_out1;

  Logical_Operator_out9543_out1 <= Logical_Operator_out7367_out1 XOR Logical_Operator_out7623_out1;

  Logical_Operator_out9544_out1 <= Logical_Operator_out7368_out1 XOR Logical_Operator_out7624_out1;

  Logical_Operator_out9545_out1 <= Logical_Operator_out7369_out1 XOR Logical_Operator_out7625_out1;

  Logical_Operator_out9546_out1 <= Logical_Operator_out7370_out1 XOR Logical_Operator_out7626_out1;

  Logical_Operator_out9547_out1 <= Logical_Operator_out7371_out1 XOR Logical_Operator_out7627_out1;

  Logical_Operator_out9548_out1 <= Logical_Operator_out7372_out1 XOR Logical_Operator_out7628_out1;

  Logical_Operator_out9549_out1 <= Logical_Operator_out7373_out1 XOR Logical_Operator_out7629_out1;

  Logical_Operator_out9550_out1 <= Logical_Operator_out7374_out1 XOR Logical_Operator_out7630_out1;

  Logical_Operator_out9551_out1 <= Logical_Operator_out7375_out1 XOR Logical_Operator_out7631_out1;

  Logical_Operator_out9552_out1 <= Logical_Operator_out7376_out1 XOR Logical_Operator_out7632_out1;

  Logical_Operator_out9553_out1 <= Logical_Operator_out7377_out1 XOR Logical_Operator_out7633_out1;

  Logical_Operator_out9554_out1 <= Logical_Operator_out7378_out1 XOR Logical_Operator_out7634_out1;

  Logical_Operator_out9555_out1 <= Logical_Operator_out7379_out1 XOR Logical_Operator_out7635_out1;

  Logical_Operator_out9556_out1 <= Logical_Operator_out7380_out1 XOR Logical_Operator_out7636_out1;

  Logical_Operator_out9557_out1 <= Logical_Operator_out7381_out1 XOR Logical_Operator_out7637_out1;

  Logical_Operator_out9558_out1 <= Logical_Operator_out7382_out1 XOR Logical_Operator_out7638_out1;

  Logical_Operator_out9559_out1 <= Logical_Operator_out7383_out1 XOR Logical_Operator_out7639_out1;

  Logical_Operator_out9560_out1 <= Logical_Operator_out7384_out1 XOR Logical_Operator_out7640_out1;

  Logical_Operator_out9561_out1 <= Logical_Operator_out7385_out1 XOR Logical_Operator_out7641_out1;

  Logical_Operator_out9562_out1 <= Logical_Operator_out7386_out1 XOR Logical_Operator_out7642_out1;

  Logical_Operator_out9563_out1 <= Logical_Operator_out7387_out1 XOR Logical_Operator_out7643_out1;

  Logical_Operator_out9564_out1 <= Logical_Operator_out7388_out1 XOR Logical_Operator_out7644_out1;

  Logical_Operator_out9565_out1 <= Logical_Operator_out7389_out1 XOR Logical_Operator_out7645_out1;

  Logical_Operator_out9566_out1 <= Logical_Operator_out7390_out1 XOR Logical_Operator_out7646_out1;

  Logical_Operator_out9567_out1 <= Logical_Operator_out7391_out1 XOR Logical_Operator_out7647_out1;

  Logical_Operator_out9568_out1 <= Logical_Operator_out7392_out1 XOR Logical_Operator_out7648_out1;

  Logical_Operator_out9569_out1 <= Logical_Operator_out7393_out1 XOR Logical_Operator_out7649_out1;

  Logical_Operator_out9570_out1 <= Logical_Operator_out7394_out1 XOR Logical_Operator_out7650_out1;

  Logical_Operator_out9571_out1 <= Logical_Operator_out7395_out1 XOR Logical_Operator_out7651_out1;

  Logical_Operator_out9572_out1 <= Logical_Operator_out7396_out1 XOR Logical_Operator_out7652_out1;

  Logical_Operator_out9573_out1 <= Logical_Operator_out7397_out1 XOR Logical_Operator_out7653_out1;

  Logical_Operator_out9574_out1 <= Logical_Operator_out7398_out1 XOR Logical_Operator_out7654_out1;

  Logical_Operator_out9575_out1 <= Logical_Operator_out7399_out1 XOR Logical_Operator_out7655_out1;

  Logical_Operator_out9576_out1 <= Logical_Operator_out7400_out1 XOR Logical_Operator_out7656_out1;

  Logical_Operator_out9577_out1 <= Logical_Operator_out7401_out1 XOR Logical_Operator_out7657_out1;

  Logical_Operator_out9578_out1 <= Logical_Operator_out7402_out1 XOR Logical_Operator_out7658_out1;

  Logical_Operator_out9579_out1 <= Logical_Operator_out7403_out1 XOR Logical_Operator_out7659_out1;

  Logical_Operator_out9580_out1 <= Logical_Operator_out7404_out1 XOR Logical_Operator_out7660_out1;

  Logical_Operator_out9581_out1 <= Logical_Operator_out7405_out1 XOR Logical_Operator_out7661_out1;

  Logical_Operator_out9582_out1 <= Logical_Operator_out7406_out1 XOR Logical_Operator_out7662_out1;

  Logical_Operator_out9583_out1 <= Logical_Operator_out7407_out1 XOR Logical_Operator_out7663_out1;

  Logical_Operator_out9584_out1 <= Logical_Operator_out7408_out1 XOR Logical_Operator_out7664_out1;

  Logical_Operator_out9585_out1 <= Logical_Operator_out7409_out1 XOR Logical_Operator_out7665_out1;

  Logical_Operator_out9586_out1 <= Logical_Operator_out7410_out1 XOR Logical_Operator_out7666_out1;

  Logical_Operator_out9587_out1 <= Logical_Operator_out7411_out1 XOR Logical_Operator_out7667_out1;

  Logical_Operator_out9588_out1 <= Logical_Operator_out7412_out1 XOR Logical_Operator_out7668_out1;

  Logical_Operator_out9589_out1 <= Logical_Operator_out7413_out1 XOR Logical_Operator_out7669_out1;

  Logical_Operator_out9590_out1 <= Logical_Operator_out7414_out1 XOR Logical_Operator_out7670_out1;

  Logical_Operator_out9591_out1 <= Logical_Operator_out7415_out1 XOR Logical_Operator_out7671_out1;

  Logical_Operator_out9592_out1 <= Logical_Operator_out7416_out1 XOR Logical_Operator_out7672_out1;

  Logical_Operator_out9593_out1 <= Logical_Operator_out7417_out1 XOR Logical_Operator_out7673_out1;

  Logical_Operator_out9594_out1 <= Logical_Operator_out7418_out1 XOR Logical_Operator_out7674_out1;

  Logical_Operator_out9595_out1 <= Logical_Operator_out7419_out1 XOR Logical_Operator_out7675_out1;

  Logical_Operator_out9596_out1 <= Logical_Operator_out7420_out1 XOR Logical_Operator_out7676_out1;

  Logical_Operator_out9597_out1 <= Logical_Operator_out7421_out1 XOR Logical_Operator_out7677_out1;

  Logical_Operator_out9598_out1 <= Logical_Operator_out7422_out1 XOR Logical_Operator_out7678_out1;

  Logical_Operator_out9599_out1 <= Logical_Operator_out7423_out1 XOR Logical_Operator_out7679_out1;

  Logical_Operator_out9600_out1 <= Logical_Operator_out7424_out1 XOR Logical_Operator_out7680_out1;

  Logical_Operator_out9601_out1 <= Logical_Operator_out6337_out1 XOR Logical_Operator_out6593_out1;

  Logical_Operator_out9602_out1 <= Logical_Operator_out6338_out1 XOR Logical_Operator_out6594_out1;

  Logical_Operator_out9603_out1 <= Logical_Operator_out6339_out1 XOR Logical_Operator_out6595_out1;

  Logical_Operator_out9604_out1 <= Logical_Operator_out6340_out1 XOR Logical_Operator_out6596_out1;

  Logical_Operator_out9605_out1 <= Logical_Operator_out6341_out1 XOR Logical_Operator_out6597_out1;

  Logical_Operator_out9606_out1 <= Logical_Operator_out6342_out1 XOR Logical_Operator_out6598_out1;

  Logical_Operator_out9607_out1 <= Logical_Operator_out6343_out1 XOR Logical_Operator_out6599_out1;

  Logical_Operator_out9608_out1 <= Logical_Operator_out6344_out1 XOR Logical_Operator_out6600_out1;

  Logical_Operator_out9609_out1 <= Logical_Operator_out6345_out1 XOR Logical_Operator_out6601_out1;

  Logical_Operator_out9610_out1 <= Logical_Operator_out6346_out1 XOR Logical_Operator_out6602_out1;

  Logical_Operator_out9611_out1 <= Logical_Operator_out6347_out1 XOR Logical_Operator_out6603_out1;

  Logical_Operator_out9612_out1 <= Logical_Operator_out6348_out1 XOR Logical_Operator_out6604_out1;

  Logical_Operator_out9613_out1 <= Logical_Operator_out6349_out1 XOR Logical_Operator_out6605_out1;

  Logical_Operator_out9614_out1 <= Logical_Operator_out6350_out1 XOR Logical_Operator_out6606_out1;

  Logical_Operator_out9615_out1 <= Logical_Operator_out6351_out1 XOR Logical_Operator_out6607_out1;

  Logical_Operator_out9616_out1 <= Logical_Operator_out6352_out1 XOR Logical_Operator_out6608_out1;

  Logical_Operator_out9617_out1 <= Logical_Operator_out6353_out1 XOR Logical_Operator_out6609_out1;

  Logical_Operator_out9618_out1 <= Logical_Operator_out6354_out1 XOR Logical_Operator_out6610_out1;

  Logical_Operator_out9619_out1 <= Logical_Operator_out6355_out1 XOR Logical_Operator_out6611_out1;

  Logical_Operator_out9620_out1 <= Logical_Operator_out6356_out1 XOR Logical_Operator_out6612_out1;

  Logical_Operator_out9621_out1 <= Logical_Operator_out6357_out1 XOR Logical_Operator_out6613_out1;

  Logical_Operator_out9622_out1 <= Logical_Operator_out6358_out1 XOR Logical_Operator_out6614_out1;

  Logical_Operator_out9623_out1 <= Logical_Operator_out6359_out1 XOR Logical_Operator_out6615_out1;

  Logical_Operator_out9624_out1 <= Logical_Operator_out6360_out1 XOR Logical_Operator_out6616_out1;

  Logical_Operator_out9625_out1 <= Logical_Operator_out6361_out1 XOR Logical_Operator_out6617_out1;

  Logical_Operator_out9626_out1 <= Logical_Operator_out6362_out1 XOR Logical_Operator_out6618_out1;

  Logical_Operator_out9627_out1 <= Logical_Operator_out6363_out1 XOR Logical_Operator_out6619_out1;

  Logical_Operator_out9628_out1 <= Logical_Operator_out6364_out1 XOR Logical_Operator_out6620_out1;

  Logical_Operator_out9629_out1 <= Logical_Operator_out6365_out1 XOR Logical_Operator_out6621_out1;

  Logical_Operator_out9630_out1 <= Logical_Operator_out6366_out1 XOR Logical_Operator_out6622_out1;

  Logical_Operator_out9631_out1 <= Logical_Operator_out6367_out1 XOR Logical_Operator_out6623_out1;

  Logical_Operator_out9632_out1 <= Logical_Operator_out6368_out1 XOR Logical_Operator_out6624_out1;

  Logical_Operator_out9633_out1 <= Logical_Operator_out6369_out1 XOR Logical_Operator_out6625_out1;

  Logical_Operator_out9634_out1 <= Logical_Operator_out6370_out1 XOR Logical_Operator_out6626_out1;

  Logical_Operator_out9635_out1 <= Logical_Operator_out6371_out1 XOR Logical_Operator_out6627_out1;

  Logical_Operator_out9636_out1 <= Logical_Operator_out6372_out1 XOR Logical_Operator_out6628_out1;

  Logical_Operator_out9637_out1 <= Logical_Operator_out6373_out1 XOR Logical_Operator_out6629_out1;

  Logical_Operator_out9638_out1 <= Logical_Operator_out6374_out1 XOR Logical_Operator_out6630_out1;

  Logical_Operator_out9639_out1 <= Logical_Operator_out6375_out1 XOR Logical_Operator_out6631_out1;

  Logical_Operator_out9640_out1 <= Logical_Operator_out6376_out1 XOR Logical_Operator_out6632_out1;

  Logical_Operator_out9641_out1 <= Logical_Operator_out6377_out1 XOR Logical_Operator_out6633_out1;

  Logical_Operator_out9642_out1 <= Logical_Operator_out6378_out1 XOR Logical_Operator_out6634_out1;

  Logical_Operator_out9643_out1 <= Logical_Operator_out6379_out1 XOR Logical_Operator_out6635_out1;

  Logical_Operator_out9644_out1 <= Logical_Operator_out6380_out1 XOR Logical_Operator_out6636_out1;

  Logical_Operator_out9645_out1 <= Logical_Operator_out6381_out1 XOR Logical_Operator_out6637_out1;

  Logical_Operator_out9646_out1 <= Logical_Operator_out6382_out1 XOR Logical_Operator_out6638_out1;

  Logical_Operator_out9647_out1 <= Logical_Operator_out6383_out1 XOR Logical_Operator_out6639_out1;

  Logical_Operator_out9648_out1 <= Logical_Operator_out6384_out1 XOR Logical_Operator_out6640_out1;

  Logical_Operator_out9649_out1 <= Logical_Operator_out6385_out1 XOR Logical_Operator_out6641_out1;

  Logical_Operator_out9650_out1 <= Logical_Operator_out6386_out1 XOR Logical_Operator_out6642_out1;

  Logical_Operator_out9651_out1 <= Logical_Operator_out6387_out1 XOR Logical_Operator_out6643_out1;

  Logical_Operator_out9652_out1 <= Logical_Operator_out6388_out1 XOR Logical_Operator_out6644_out1;

  Logical_Operator_out9653_out1 <= Logical_Operator_out6389_out1 XOR Logical_Operator_out6645_out1;

  Logical_Operator_out9654_out1 <= Logical_Operator_out6390_out1 XOR Logical_Operator_out6646_out1;

  Logical_Operator_out9655_out1 <= Logical_Operator_out6391_out1 XOR Logical_Operator_out6647_out1;

  Logical_Operator_out9656_out1 <= Logical_Operator_out6392_out1 XOR Logical_Operator_out6648_out1;

  Logical_Operator_out9657_out1 <= Logical_Operator_out6393_out1 XOR Logical_Operator_out6649_out1;

  Logical_Operator_out9658_out1 <= Logical_Operator_out6394_out1 XOR Logical_Operator_out6650_out1;

  Logical_Operator_out9659_out1 <= Logical_Operator_out6395_out1 XOR Logical_Operator_out6651_out1;

  Logical_Operator_out9660_out1 <= Logical_Operator_out6396_out1 XOR Logical_Operator_out6652_out1;

  Logical_Operator_out9661_out1 <= Logical_Operator_out6397_out1 XOR Logical_Operator_out6653_out1;

  Logical_Operator_out9662_out1 <= Logical_Operator_out6398_out1 XOR Logical_Operator_out6654_out1;

  Logical_Operator_out9663_out1 <= Logical_Operator_out6399_out1 XOR Logical_Operator_out6655_out1;

  Logical_Operator_out9664_out1 <= Logical_Operator_out6400_out1 XOR Logical_Operator_out6656_out1;

  Logical_Operator_out9665_out1 <= Logical_Operator_out5345_out1 XOR Logical_Operator_out5601_out1;

  Logical_Operator_out9666_out1 <= Logical_Operator_out5346_out1 XOR Logical_Operator_out5602_out1;

  Logical_Operator_out9667_out1 <= Logical_Operator_out5347_out1 XOR Logical_Operator_out5603_out1;

  Logical_Operator_out9668_out1 <= Logical_Operator_out5348_out1 XOR Logical_Operator_out5604_out1;

  Logical_Operator_out9669_out1 <= Logical_Operator_out5349_out1 XOR Logical_Operator_out5605_out1;

  Logical_Operator_out9670_out1 <= Logical_Operator_out5350_out1 XOR Logical_Operator_out5606_out1;

  Logical_Operator_out9671_out1 <= Logical_Operator_out5351_out1 XOR Logical_Operator_out5607_out1;

  Logical_Operator_out9672_out1 <= Logical_Operator_out5352_out1 XOR Logical_Operator_out5608_out1;

  Logical_Operator_out9673_out1 <= Logical_Operator_out5353_out1 XOR Logical_Operator_out5609_out1;

  Logical_Operator_out9674_out1 <= Logical_Operator_out5354_out1 XOR Logical_Operator_out5610_out1;

  Logical_Operator_out9675_out1 <= Logical_Operator_out5355_out1 XOR Logical_Operator_out5611_out1;

  Logical_Operator_out9676_out1 <= Logical_Operator_out5356_out1 XOR Logical_Operator_out5612_out1;

  Logical_Operator_out9677_out1 <= Logical_Operator_out5357_out1 XOR Logical_Operator_out5613_out1;

  Logical_Operator_out9678_out1 <= Logical_Operator_out5358_out1 XOR Logical_Operator_out5614_out1;

  Logical_Operator_out9679_out1 <= Logical_Operator_out5359_out1 XOR Logical_Operator_out5615_out1;

  Logical_Operator_out9680_out1 <= Logical_Operator_out5360_out1 XOR Logical_Operator_out5616_out1;

  Logical_Operator_out9681_out1 <= Logical_Operator_out5361_out1 XOR Logical_Operator_out5617_out1;

  Logical_Operator_out9682_out1 <= Logical_Operator_out5362_out1 XOR Logical_Operator_out5618_out1;

  Logical_Operator_out9683_out1 <= Logical_Operator_out5363_out1 XOR Logical_Operator_out5619_out1;

  Logical_Operator_out9684_out1 <= Logical_Operator_out5364_out1 XOR Logical_Operator_out5620_out1;

  Logical_Operator_out9685_out1 <= Logical_Operator_out5365_out1 XOR Logical_Operator_out5621_out1;

  Logical_Operator_out9686_out1 <= Logical_Operator_out5366_out1 XOR Logical_Operator_out5622_out1;

  Logical_Operator_out9687_out1 <= Logical_Operator_out5367_out1 XOR Logical_Operator_out5623_out1;

  Logical_Operator_out9688_out1 <= Logical_Operator_out5368_out1 XOR Logical_Operator_out5624_out1;

  Logical_Operator_out9689_out1 <= Logical_Operator_out5369_out1 XOR Logical_Operator_out5625_out1;

  Logical_Operator_out9690_out1 <= Logical_Operator_out5370_out1 XOR Logical_Operator_out5626_out1;

  Logical_Operator_out9691_out1 <= Logical_Operator_out5371_out1 XOR Logical_Operator_out5627_out1;

  Logical_Operator_out9692_out1 <= Logical_Operator_out5372_out1 XOR Logical_Operator_out5628_out1;

  Logical_Operator_out9693_out1 <= Logical_Operator_out5373_out1 XOR Logical_Operator_out5629_out1;

  Logical_Operator_out9694_out1 <= Logical_Operator_out5374_out1 XOR Logical_Operator_out5630_out1;

  Logical_Operator_out9695_out1 <= Logical_Operator_out5375_out1 XOR Logical_Operator_out5631_out1;

  Logical_Operator_out9696_out1 <= Logical_Operator_out5376_out1 XOR Logical_Operator_out5632_out1;

  Logical_Operator_out9697_out1 <= Logical_Operator_out4337_out1 XOR Logical_Operator_out4593_out1;

  Logical_Operator_out9698_out1 <= Logical_Operator_out4338_out1 XOR Logical_Operator_out4594_out1;

  Logical_Operator_out9699_out1 <= Logical_Operator_out4339_out1 XOR Logical_Operator_out4595_out1;

  Logical_Operator_out9700_out1 <= Logical_Operator_out4340_out1 XOR Logical_Operator_out4596_out1;

  Logical_Operator_out9701_out1 <= Logical_Operator_out4341_out1 XOR Logical_Operator_out4597_out1;

  Logical_Operator_out9702_out1 <= Logical_Operator_out4342_out1 XOR Logical_Operator_out4598_out1;

  Logical_Operator_out9703_out1 <= Logical_Operator_out4343_out1 XOR Logical_Operator_out4599_out1;

  Logical_Operator_out9704_out1 <= Logical_Operator_out4344_out1 XOR Logical_Operator_out4600_out1;

  Logical_Operator_out9705_out1 <= Logical_Operator_out4345_out1 XOR Logical_Operator_out4601_out1;

  Logical_Operator_out9706_out1 <= Logical_Operator_out4346_out1 XOR Logical_Operator_out4602_out1;

  Logical_Operator_out9707_out1 <= Logical_Operator_out4347_out1 XOR Logical_Operator_out4603_out1;

  Logical_Operator_out9708_out1 <= Logical_Operator_out4348_out1 XOR Logical_Operator_out4604_out1;

  Logical_Operator_out9709_out1 <= Logical_Operator_out4349_out1 XOR Logical_Operator_out4605_out1;

  Logical_Operator_out9710_out1 <= Logical_Operator_out4350_out1 XOR Logical_Operator_out4606_out1;

  Logical_Operator_out9711_out1 <= Logical_Operator_out4351_out1 XOR Logical_Operator_out4607_out1;

  Logical_Operator_out9712_out1 <= Logical_Operator_out4352_out1 XOR Logical_Operator_out4608_out1;

  Logical_Operator_out9713_out1 <= Logical_Operator_out3321_out1 XOR Logical_Operator_out3577_out1;

  Logical_Operator_out9714_out1 <= Logical_Operator_out3322_out1 XOR Logical_Operator_out3578_out1;

  Logical_Operator_out9715_out1 <= Logical_Operator_out3323_out1 XOR Logical_Operator_out3579_out1;

  Logical_Operator_out9716_out1 <= Logical_Operator_out3324_out1 XOR Logical_Operator_out3580_out1;

  Logical_Operator_out9717_out1 <= Logical_Operator_out3325_out1 XOR Logical_Operator_out3581_out1;

  Logical_Operator_out9718_out1 <= Logical_Operator_out3326_out1 XOR Logical_Operator_out3582_out1;

  Logical_Operator_out9719_out1 <= Logical_Operator_out3327_out1 XOR Logical_Operator_out3583_out1;

  Logical_Operator_out9720_out1 <= Logical_Operator_out3328_out1 XOR Logical_Operator_out3584_out1;

  Logical_Operator_out9721_out1 <= Logical_Operator_out2301_out1 XOR Logical_Operator_out2557_out1;

  Logical_Operator_out9722_out1 <= Logical_Operator_out2302_out1 XOR Logical_Operator_out2558_out1;

  Logical_Operator_out9723_out1 <= Logical_Operator_out2303_out1 XOR Logical_Operator_out2559_out1;

  Logical_Operator_out9724_out1 <= Logical_Operator_out2304_out1 XOR Logical_Operator_out2560_out1;

  Logical_Operator_out9725_out1 <= Logical_Operator_out1279_out1 XOR Logical_Operator_out1535_out1;

  Logical_Operator_out9726_out1 <= Logical_Operator_out1280_out1 XOR Logical_Operator_out1536_out1;

  Logical_Operator_out9727_out1 <= Logical_Operator_out256_out1 XOR Logical_Operator_out512_out1;

  Logical_Operator_out9728_out1 <= in512 XOR in1024;

  Logical_Operator_out9729_out1 <= Logical_Operator_out8705_out1 XOR Logical_Operator_out8961_out1;

  Logical_Operator_out9730_out1 <= Logical_Operator_out8706_out1 XOR Logical_Operator_out8962_out1;

  Logical_Operator_out9731_out1 <= Logical_Operator_out8707_out1 XOR Logical_Operator_out8963_out1;

  Logical_Operator_out9732_out1 <= Logical_Operator_out8708_out1 XOR Logical_Operator_out8964_out1;

  Logical_Operator_out9733_out1 <= Logical_Operator_out8709_out1 XOR Logical_Operator_out8965_out1;

  Logical_Operator_out9734_out1 <= Logical_Operator_out8710_out1 XOR Logical_Operator_out8966_out1;

  Logical_Operator_out9735_out1 <= Logical_Operator_out8711_out1 XOR Logical_Operator_out8967_out1;

  Logical_Operator_out9736_out1 <= Logical_Operator_out8712_out1 XOR Logical_Operator_out8968_out1;

  Logical_Operator_out9737_out1 <= Logical_Operator_out8713_out1 XOR Logical_Operator_out8969_out1;

  Logical_Operator_out9738_out1 <= Logical_Operator_out8714_out1 XOR Logical_Operator_out8970_out1;

  Logical_Operator_out9739_out1 <= Logical_Operator_out8715_out1 XOR Logical_Operator_out8971_out1;

  Logical_Operator_out9740_out1 <= Logical_Operator_out8716_out1 XOR Logical_Operator_out8972_out1;

  Logical_Operator_out9741_out1 <= Logical_Operator_out8717_out1 XOR Logical_Operator_out8973_out1;

  Logical_Operator_out9742_out1 <= Logical_Operator_out8718_out1 XOR Logical_Operator_out8974_out1;

  Logical_Operator_out9743_out1 <= Logical_Operator_out8719_out1 XOR Logical_Operator_out8975_out1;

  Logical_Operator_out9744_out1 <= Logical_Operator_out8720_out1 XOR Logical_Operator_out8976_out1;

  Logical_Operator_out9745_out1 <= Logical_Operator_out8721_out1 XOR Logical_Operator_out8977_out1;

  Logical_Operator_out9746_out1 <= Logical_Operator_out8722_out1 XOR Logical_Operator_out8978_out1;

  Logical_Operator_out9747_out1 <= Logical_Operator_out8723_out1 XOR Logical_Operator_out8979_out1;

  Logical_Operator_out9748_out1 <= Logical_Operator_out8724_out1 XOR Logical_Operator_out8980_out1;

  Logical_Operator_out9749_out1 <= Logical_Operator_out8725_out1 XOR Logical_Operator_out8981_out1;

  Logical_Operator_out9750_out1 <= Logical_Operator_out8726_out1 XOR Logical_Operator_out8982_out1;

  Logical_Operator_out9751_out1 <= Logical_Operator_out8727_out1 XOR Logical_Operator_out8983_out1;

  Logical_Operator_out9752_out1 <= Logical_Operator_out8728_out1 XOR Logical_Operator_out8984_out1;

  Logical_Operator_out9753_out1 <= Logical_Operator_out8729_out1 XOR Logical_Operator_out8985_out1;

  Logical_Operator_out9754_out1 <= Logical_Operator_out8730_out1 XOR Logical_Operator_out8986_out1;

  Logical_Operator_out9755_out1 <= Logical_Operator_out8731_out1 XOR Logical_Operator_out8987_out1;

  Logical_Operator_out9756_out1 <= Logical_Operator_out8732_out1 XOR Logical_Operator_out8988_out1;

  Logical_Operator_out9757_out1 <= Logical_Operator_out8733_out1 XOR Logical_Operator_out8989_out1;

  Logical_Operator_out9758_out1 <= Logical_Operator_out8734_out1 XOR Logical_Operator_out8990_out1;

  Logical_Operator_out9759_out1 <= Logical_Operator_out8735_out1 XOR Logical_Operator_out8991_out1;

  Logical_Operator_out9760_out1 <= Logical_Operator_out8736_out1 XOR Logical_Operator_out8992_out1;

  Logical_Operator_out9761_out1 <= Logical_Operator_out8737_out1 XOR Logical_Operator_out8993_out1;

  Logical_Operator_out9762_out1 <= Logical_Operator_out8738_out1 XOR Logical_Operator_out8994_out1;

  Logical_Operator_out9763_out1 <= Logical_Operator_out8739_out1 XOR Logical_Operator_out8995_out1;

  Logical_Operator_out9764_out1 <= Logical_Operator_out8740_out1 XOR Logical_Operator_out8996_out1;

  Logical_Operator_out9765_out1 <= Logical_Operator_out8741_out1 XOR Logical_Operator_out8997_out1;

  Logical_Operator_out9766_out1 <= Logical_Operator_out8742_out1 XOR Logical_Operator_out8998_out1;

  Logical_Operator_out9767_out1 <= Logical_Operator_out8743_out1 XOR Logical_Operator_out8999_out1;

  Logical_Operator_out9768_out1 <= Logical_Operator_out8744_out1 XOR Logical_Operator_out9000_out1;

  Logical_Operator_out9769_out1 <= Logical_Operator_out8745_out1 XOR Logical_Operator_out9001_out1;

  Logical_Operator_out9770_out1 <= Logical_Operator_out8746_out1 XOR Logical_Operator_out9002_out1;

  Logical_Operator_out9771_out1 <= Logical_Operator_out8747_out1 XOR Logical_Operator_out9003_out1;

  Logical_Operator_out9772_out1 <= Logical_Operator_out8748_out1 XOR Logical_Operator_out9004_out1;

  Logical_Operator_out9773_out1 <= Logical_Operator_out8749_out1 XOR Logical_Operator_out9005_out1;

  Logical_Operator_out9774_out1 <= Logical_Operator_out8750_out1 XOR Logical_Operator_out9006_out1;

  Logical_Operator_out9775_out1 <= Logical_Operator_out8751_out1 XOR Logical_Operator_out9007_out1;

  Logical_Operator_out9776_out1 <= Logical_Operator_out8752_out1 XOR Logical_Operator_out9008_out1;

  Logical_Operator_out9777_out1 <= Logical_Operator_out8753_out1 XOR Logical_Operator_out9009_out1;

  Logical_Operator_out9778_out1 <= Logical_Operator_out8754_out1 XOR Logical_Operator_out9010_out1;

  Logical_Operator_out9779_out1 <= Logical_Operator_out8755_out1 XOR Logical_Operator_out9011_out1;

  Logical_Operator_out9780_out1 <= Logical_Operator_out8756_out1 XOR Logical_Operator_out9012_out1;

  Logical_Operator_out9781_out1 <= Logical_Operator_out8757_out1 XOR Logical_Operator_out9013_out1;

  Logical_Operator_out9782_out1 <= Logical_Operator_out8758_out1 XOR Logical_Operator_out9014_out1;

  Logical_Operator_out9783_out1 <= Logical_Operator_out8759_out1 XOR Logical_Operator_out9015_out1;

  Logical_Operator_out9784_out1 <= Logical_Operator_out8760_out1 XOR Logical_Operator_out9016_out1;

  Logical_Operator_out9785_out1 <= Logical_Operator_out8761_out1 XOR Logical_Operator_out9017_out1;

  Logical_Operator_out9786_out1 <= Logical_Operator_out8762_out1 XOR Logical_Operator_out9018_out1;

  Logical_Operator_out9787_out1 <= Logical_Operator_out8763_out1 XOR Logical_Operator_out9019_out1;

  Logical_Operator_out9788_out1 <= Logical_Operator_out8764_out1 XOR Logical_Operator_out9020_out1;

  Logical_Operator_out9789_out1 <= Logical_Operator_out8765_out1 XOR Logical_Operator_out9021_out1;

  Logical_Operator_out9790_out1 <= Logical_Operator_out8766_out1 XOR Logical_Operator_out9022_out1;

  Logical_Operator_out9791_out1 <= Logical_Operator_out8767_out1 XOR Logical_Operator_out9023_out1;

  Logical_Operator_out9792_out1 <= Logical_Operator_out8768_out1 XOR Logical_Operator_out9024_out1;

  Logical_Operator_out9793_out1 <= Logical_Operator_out8769_out1 XOR Logical_Operator_out9025_out1;

  Logical_Operator_out9794_out1 <= Logical_Operator_out8770_out1 XOR Logical_Operator_out9026_out1;

  Logical_Operator_out9795_out1 <= Logical_Operator_out8771_out1 XOR Logical_Operator_out9027_out1;

  Logical_Operator_out9796_out1 <= Logical_Operator_out8772_out1 XOR Logical_Operator_out9028_out1;

  Logical_Operator_out9797_out1 <= Logical_Operator_out8773_out1 XOR Logical_Operator_out9029_out1;

  Logical_Operator_out9798_out1 <= Logical_Operator_out8774_out1 XOR Logical_Operator_out9030_out1;

  Logical_Operator_out9799_out1 <= Logical_Operator_out8775_out1 XOR Logical_Operator_out9031_out1;

  Logical_Operator_out9800_out1 <= Logical_Operator_out8776_out1 XOR Logical_Operator_out9032_out1;

  Logical_Operator_out9801_out1 <= Logical_Operator_out8777_out1 XOR Logical_Operator_out9033_out1;

  Logical_Operator_out9802_out1 <= Logical_Operator_out8778_out1 XOR Logical_Operator_out9034_out1;

  Logical_Operator_out9803_out1 <= Logical_Operator_out8779_out1 XOR Logical_Operator_out9035_out1;

  Logical_Operator_out9804_out1 <= Logical_Operator_out8780_out1 XOR Logical_Operator_out9036_out1;

  Logical_Operator_out9805_out1 <= Logical_Operator_out8781_out1 XOR Logical_Operator_out9037_out1;

  Logical_Operator_out9806_out1 <= Logical_Operator_out8782_out1 XOR Logical_Operator_out9038_out1;

  Logical_Operator_out9807_out1 <= Logical_Operator_out8783_out1 XOR Logical_Operator_out9039_out1;

  Logical_Operator_out9808_out1 <= Logical_Operator_out8784_out1 XOR Logical_Operator_out9040_out1;

  Logical_Operator_out9809_out1 <= Logical_Operator_out8785_out1 XOR Logical_Operator_out9041_out1;

  Logical_Operator_out9810_out1 <= Logical_Operator_out8786_out1 XOR Logical_Operator_out9042_out1;

  Logical_Operator_out9811_out1 <= Logical_Operator_out8787_out1 XOR Logical_Operator_out9043_out1;

  Logical_Operator_out9812_out1 <= Logical_Operator_out8788_out1 XOR Logical_Operator_out9044_out1;

  Logical_Operator_out9813_out1 <= Logical_Operator_out8789_out1 XOR Logical_Operator_out9045_out1;

  Logical_Operator_out9814_out1 <= Logical_Operator_out8790_out1 XOR Logical_Operator_out9046_out1;

  Logical_Operator_out9815_out1 <= Logical_Operator_out8791_out1 XOR Logical_Operator_out9047_out1;

  Logical_Operator_out9816_out1 <= Logical_Operator_out8792_out1 XOR Logical_Operator_out9048_out1;

  Logical_Operator_out9817_out1 <= Logical_Operator_out8793_out1 XOR Logical_Operator_out9049_out1;

  Logical_Operator_out9818_out1 <= Logical_Operator_out8794_out1 XOR Logical_Operator_out9050_out1;

  Logical_Operator_out9819_out1 <= Logical_Operator_out8795_out1 XOR Logical_Operator_out9051_out1;

  Logical_Operator_out9820_out1 <= Logical_Operator_out8796_out1 XOR Logical_Operator_out9052_out1;

  Logical_Operator_out9821_out1 <= Logical_Operator_out8797_out1 XOR Logical_Operator_out9053_out1;

  Logical_Operator_out9822_out1 <= Logical_Operator_out8798_out1 XOR Logical_Operator_out9054_out1;

  Logical_Operator_out9823_out1 <= Logical_Operator_out8799_out1 XOR Logical_Operator_out9055_out1;

  Logical_Operator_out9824_out1 <= Logical_Operator_out8800_out1 XOR Logical_Operator_out9056_out1;

  Logical_Operator_out9825_out1 <= Logical_Operator_out8801_out1 XOR Logical_Operator_out9057_out1;

  Logical_Operator_out9826_out1 <= Logical_Operator_out8802_out1 XOR Logical_Operator_out9058_out1;

  Logical_Operator_out9827_out1 <= Logical_Operator_out8803_out1 XOR Logical_Operator_out9059_out1;

  Logical_Operator_out9828_out1 <= Logical_Operator_out8804_out1 XOR Logical_Operator_out9060_out1;

  Logical_Operator_out9829_out1 <= Logical_Operator_out8805_out1 XOR Logical_Operator_out9061_out1;

  Logical_Operator_out9830_out1 <= Logical_Operator_out8806_out1 XOR Logical_Operator_out9062_out1;

  Logical_Operator_out9831_out1 <= Logical_Operator_out8807_out1 XOR Logical_Operator_out9063_out1;

  Logical_Operator_out9832_out1 <= Logical_Operator_out8808_out1 XOR Logical_Operator_out9064_out1;

  Logical_Operator_out9833_out1 <= Logical_Operator_out8809_out1 XOR Logical_Operator_out9065_out1;

  Logical_Operator_out9834_out1 <= Logical_Operator_out8810_out1 XOR Logical_Operator_out9066_out1;

  Logical_Operator_out9835_out1 <= Logical_Operator_out8811_out1 XOR Logical_Operator_out9067_out1;

  Logical_Operator_out9836_out1 <= Logical_Operator_out8812_out1 XOR Logical_Operator_out9068_out1;

  Logical_Operator_out9837_out1 <= Logical_Operator_out8813_out1 XOR Logical_Operator_out9069_out1;

  Logical_Operator_out9838_out1 <= Logical_Operator_out8814_out1 XOR Logical_Operator_out9070_out1;

  Logical_Operator_out9839_out1 <= Logical_Operator_out8815_out1 XOR Logical_Operator_out9071_out1;

  Logical_Operator_out9840_out1 <= Logical_Operator_out8816_out1 XOR Logical_Operator_out9072_out1;

  Logical_Operator_out9841_out1 <= Logical_Operator_out8817_out1 XOR Logical_Operator_out9073_out1;

  Logical_Operator_out9842_out1 <= Logical_Operator_out8818_out1 XOR Logical_Operator_out9074_out1;

  Logical_Operator_out9843_out1 <= Logical_Operator_out8819_out1 XOR Logical_Operator_out9075_out1;

  Logical_Operator_out9844_out1 <= Logical_Operator_out8820_out1 XOR Logical_Operator_out9076_out1;

  Logical_Operator_out9845_out1 <= Logical_Operator_out8821_out1 XOR Logical_Operator_out9077_out1;

  Logical_Operator_out9846_out1 <= Logical_Operator_out8822_out1 XOR Logical_Operator_out9078_out1;

  Logical_Operator_out9847_out1 <= Logical_Operator_out8823_out1 XOR Logical_Operator_out9079_out1;

  Logical_Operator_out9848_out1 <= Logical_Operator_out8824_out1 XOR Logical_Operator_out9080_out1;

  Logical_Operator_out9849_out1 <= Logical_Operator_out8825_out1 XOR Logical_Operator_out9081_out1;

  Logical_Operator_out9850_out1 <= Logical_Operator_out8826_out1 XOR Logical_Operator_out9082_out1;

  Logical_Operator_out9851_out1 <= Logical_Operator_out8827_out1 XOR Logical_Operator_out9083_out1;

  Logical_Operator_out9852_out1 <= Logical_Operator_out8828_out1 XOR Logical_Operator_out9084_out1;

  Logical_Operator_out9853_out1 <= Logical_Operator_out8829_out1 XOR Logical_Operator_out9085_out1;

  Logical_Operator_out9854_out1 <= Logical_Operator_out8830_out1 XOR Logical_Operator_out9086_out1;

  Logical_Operator_out9855_out1 <= Logical_Operator_out8831_out1 XOR Logical_Operator_out9087_out1;

  Logical_Operator_out9856_out1 <= Logical_Operator_out8832_out1 XOR Logical_Operator_out9088_out1;

  Logical_Operator_out9857_out1 <= Logical_Operator_out8833_out1 XOR Logical_Operator_out9089_out1;

  Logical_Operator_out9858_out1 <= Logical_Operator_out8834_out1 XOR Logical_Operator_out9090_out1;

  Logical_Operator_out9859_out1 <= Logical_Operator_out8835_out1 XOR Logical_Operator_out9091_out1;

  Logical_Operator_out9860_out1 <= Logical_Operator_out8836_out1 XOR Logical_Operator_out9092_out1;

  Logical_Operator_out9861_out1 <= Logical_Operator_out8837_out1 XOR Logical_Operator_out9093_out1;

  Logical_Operator_out9862_out1 <= Logical_Operator_out8838_out1 XOR Logical_Operator_out9094_out1;

  Logical_Operator_out9863_out1 <= Logical_Operator_out8839_out1 XOR Logical_Operator_out9095_out1;

  Logical_Operator_out9864_out1 <= Logical_Operator_out8840_out1 XOR Logical_Operator_out9096_out1;

  Logical_Operator_out9865_out1 <= Logical_Operator_out8841_out1 XOR Logical_Operator_out9097_out1;

  Logical_Operator_out9866_out1 <= Logical_Operator_out8842_out1 XOR Logical_Operator_out9098_out1;

  Logical_Operator_out9867_out1 <= Logical_Operator_out8843_out1 XOR Logical_Operator_out9099_out1;

  Logical_Operator_out9868_out1 <= Logical_Operator_out8844_out1 XOR Logical_Operator_out9100_out1;

  Logical_Operator_out9869_out1 <= Logical_Operator_out8845_out1 XOR Logical_Operator_out9101_out1;

  Logical_Operator_out9870_out1 <= Logical_Operator_out8846_out1 XOR Logical_Operator_out9102_out1;

  Logical_Operator_out9871_out1 <= Logical_Operator_out8847_out1 XOR Logical_Operator_out9103_out1;

  Logical_Operator_out9872_out1 <= Logical_Operator_out8848_out1 XOR Logical_Operator_out9104_out1;

  Logical_Operator_out9873_out1 <= Logical_Operator_out8849_out1 XOR Logical_Operator_out9105_out1;

  Logical_Operator_out9874_out1 <= Logical_Operator_out8850_out1 XOR Logical_Operator_out9106_out1;

  Logical_Operator_out9875_out1 <= Logical_Operator_out8851_out1 XOR Logical_Operator_out9107_out1;

  Logical_Operator_out9876_out1 <= Logical_Operator_out8852_out1 XOR Logical_Operator_out9108_out1;

  Logical_Operator_out9877_out1 <= Logical_Operator_out8853_out1 XOR Logical_Operator_out9109_out1;

  Logical_Operator_out9878_out1 <= Logical_Operator_out8854_out1 XOR Logical_Operator_out9110_out1;

  Logical_Operator_out9879_out1 <= Logical_Operator_out8855_out1 XOR Logical_Operator_out9111_out1;

  Logical_Operator_out9880_out1 <= Logical_Operator_out8856_out1 XOR Logical_Operator_out9112_out1;

  Logical_Operator_out9881_out1 <= Logical_Operator_out8857_out1 XOR Logical_Operator_out9113_out1;

  Logical_Operator_out9882_out1 <= Logical_Operator_out8858_out1 XOR Logical_Operator_out9114_out1;

  Logical_Operator_out9883_out1 <= Logical_Operator_out8859_out1 XOR Logical_Operator_out9115_out1;

  Logical_Operator_out9884_out1 <= Logical_Operator_out8860_out1 XOR Logical_Operator_out9116_out1;

  Logical_Operator_out9885_out1 <= Logical_Operator_out8861_out1 XOR Logical_Operator_out9117_out1;

  Logical_Operator_out9886_out1 <= Logical_Operator_out8862_out1 XOR Logical_Operator_out9118_out1;

  Logical_Operator_out9887_out1 <= Logical_Operator_out8863_out1 XOR Logical_Operator_out9119_out1;

  Logical_Operator_out9888_out1 <= Logical_Operator_out8864_out1 XOR Logical_Operator_out9120_out1;

  Logical_Operator_out9889_out1 <= Logical_Operator_out8865_out1 XOR Logical_Operator_out9121_out1;

  Logical_Operator_out9890_out1 <= Logical_Operator_out8866_out1 XOR Logical_Operator_out9122_out1;

  Logical_Operator_out9891_out1 <= Logical_Operator_out8867_out1 XOR Logical_Operator_out9123_out1;

  Logical_Operator_out9892_out1 <= Logical_Operator_out8868_out1 XOR Logical_Operator_out9124_out1;

  Logical_Operator_out9893_out1 <= Logical_Operator_out8869_out1 XOR Logical_Operator_out9125_out1;

  Logical_Operator_out9894_out1 <= Logical_Operator_out8870_out1 XOR Logical_Operator_out9126_out1;

  Logical_Operator_out9895_out1 <= Logical_Operator_out8871_out1 XOR Logical_Operator_out9127_out1;

  Logical_Operator_out9896_out1 <= Logical_Operator_out8872_out1 XOR Logical_Operator_out9128_out1;

  Logical_Operator_out9897_out1 <= Logical_Operator_out8873_out1 XOR Logical_Operator_out9129_out1;

  Logical_Operator_out9898_out1 <= Logical_Operator_out8874_out1 XOR Logical_Operator_out9130_out1;

  Logical_Operator_out9899_out1 <= Logical_Operator_out8875_out1 XOR Logical_Operator_out9131_out1;

  Logical_Operator_out9900_out1 <= Logical_Operator_out8876_out1 XOR Logical_Operator_out9132_out1;

  Logical_Operator_out9901_out1 <= Logical_Operator_out8877_out1 XOR Logical_Operator_out9133_out1;

  Logical_Operator_out9902_out1 <= Logical_Operator_out8878_out1 XOR Logical_Operator_out9134_out1;

  Logical_Operator_out9903_out1 <= Logical_Operator_out8879_out1 XOR Logical_Operator_out9135_out1;

  Logical_Operator_out9904_out1 <= Logical_Operator_out8880_out1 XOR Logical_Operator_out9136_out1;

  Logical_Operator_out9905_out1 <= Logical_Operator_out8881_out1 XOR Logical_Operator_out9137_out1;

  Logical_Operator_out9906_out1 <= Logical_Operator_out8882_out1 XOR Logical_Operator_out9138_out1;

  Logical_Operator_out9907_out1 <= Logical_Operator_out8883_out1 XOR Logical_Operator_out9139_out1;

  Logical_Operator_out9908_out1 <= Logical_Operator_out8884_out1 XOR Logical_Operator_out9140_out1;

  Logical_Operator_out9909_out1 <= Logical_Operator_out8885_out1 XOR Logical_Operator_out9141_out1;

  Logical_Operator_out9910_out1 <= Logical_Operator_out8886_out1 XOR Logical_Operator_out9142_out1;

  Logical_Operator_out9911_out1 <= Logical_Operator_out8887_out1 XOR Logical_Operator_out9143_out1;

  Logical_Operator_out9912_out1 <= Logical_Operator_out8888_out1 XOR Logical_Operator_out9144_out1;

  Logical_Operator_out9913_out1 <= Logical_Operator_out8889_out1 XOR Logical_Operator_out9145_out1;

  Logical_Operator_out9914_out1 <= Logical_Operator_out8890_out1 XOR Logical_Operator_out9146_out1;

  Logical_Operator_out9915_out1 <= Logical_Operator_out8891_out1 XOR Logical_Operator_out9147_out1;

  Logical_Operator_out9916_out1 <= Logical_Operator_out8892_out1 XOR Logical_Operator_out9148_out1;

  Logical_Operator_out9917_out1 <= Logical_Operator_out8893_out1 XOR Logical_Operator_out9149_out1;

  Logical_Operator_out9918_out1 <= Logical_Operator_out8894_out1 XOR Logical_Operator_out9150_out1;

  Logical_Operator_out9919_out1 <= Logical_Operator_out8895_out1 XOR Logical_Operator_out9151_out1;

  Logical_Operator_out9920_out1 <= Logical_Operator_out8896_out1 XOR Logical_Operator_out9152_out1;

  Logical_Operator_out9921_out1 <= Logical_Operator_out8897_out1 XOR Logical_Operator_out9153_out1;

  Logical_Operator_out9922_out1 <= Logical_Operator_out8898_out1 XOR Logical_Operator_out9154_out1;

  Logical_Operator_out9923_out1 <= Logical_Operator_out8899_out1 XOR Logical_Operator_out9155_out1;

  Logical_Operator_out9924_out1 <= Logical_Operator_out8900_out1 XOR Logical_Operator_out9156_out1;

  Logical_Operator_out9925_out1 <= Logical_Operator_out8901_out1 XOR Logical_Operator_out9157_out1;

  Logical_Operator_out9926_out1 <= Logical_Operator_out8902_out1 XOR Logical_Operator_out9158_out1;

  Logical_Operator_out9927_out1 <= Logical_Operator_out8903_out1 XOR Logical_Operator_out9159_out1;

  Logical_Operator_out9928_out1 <= Logical_Operator_out8904_out1 XOR Logical_Operator_out9160_out1;

  Logical_Operator_out9929_out1 <= Logical_Operator_out8905_out1 XOR Logical_Operator_out9161_out1;

  Logical_Operator_out9930_out1 <= Logical_Operator_out8906_out1 XOR Logical_Operator_out9162_out1;

  Logical_Operator_out9931_out1 <= Logical_Operator_out8907_out1 XOR Logical_Operator_out9163_out1;

  Logical_Operator_out9932_out1 <= Logical_Operator_out8908_out1 XOR Logical_Operator_out9164_out1;

  Logical_Operator_out9933_out1 <= Logical_Operator_out8909_out1 XOR Logical_Operator_out9165_out1;

  Logical_Operator_out9934_out1 <= Logical_Operator_out8910_out1 XOR Logical_Operator_out9166_out1;

  Logical_Operator_out9935_out1 <= Logical_Operator_out8911_out1 XOR Logical_Operator_out9167_out1;

  Logical_Operator_out9936_out1 <= Logical_Operator_out8912_out1 XOR Logical_Operator_out9168_out1;

  Logical_Operator_out9937_out1 <= Logical_Operator_out8913_out1 XOR Logical_Operator_out9169_out1;

  Logical_Operator_out9938_out1 <= Logical_Operator_out8914_out1 XOR Logical_Operator_out9170_out1;

  Logical_Operator_out9939_out1 <= Logical_Operator_out8915_out1 XOR Logical_Operator_out9171_out1;

  Logical_Operator_out9940_out1 <= Logical_Operator_out8916_out1 XOR Logical_Operator_out9172_out1;

  Logical_Operator_out9941_out1 <= Logical_Operator_out8917_out1 XOR Logical_Operator_out9173_out1;

  Logical_Operator_out9942_out1 <= Logical_Operator_out8918_out1 XOR Logical_Operator_out9174_out1;

  Logical_Operator_out9943_out1 <= Logical_Operator_out8919_out1 XOR Logical_Operator_out9175_out1;

  Logical_Operator_out9944_out1 <= Logical_Operator_out8920_out1 XOR Logical_Operator_out9176_out1;

  Logical_Operator_out9945_out1 <= Logical_Operator_out8921_out1 XOR Logical_Operator_out9177_out1;

  Logical_Operator_out9946_out1 <= Logical_Operator_out8922_out1 XOR Logical_Operator_out9178_out1;

  Logical_Operator_out9947_out1 <= Logical_Operator_out8923_out1 XOR Logical_Operator_out9179_out1;

  Logical_Operator_out9948_out1 <= Logical_Operator_out8924_out1 XOR Logical_Operator_out9180_out1;

  Logical_Operator_out9949_out1 <= Logical_Operator_out8925_out1 XOR Logical_Operator_out9181_out1;

  Logical_Operator_out9950_out1 <= Logical_Operator_out8926_out1 XOR Logical_Operator_out9182_out1;

  Logical_Operator_out9951_out1 <= Logical_Operator_out8927_out1 XOR Logical_Operator_out9183_out1;

  Logical_Operator_out9952_out1 <= Logical_Operator_out8928_out1 XOR Logical_Operator_out9184_out1;

  Logical_Operator_out9953_out1 <= Logical_Operator_out8929_out1 XOR Logical_Operator_out9185_out1;

  Logical_Operator_out9954_out1 <= Logical_Operator_out8930_out1 XOR Logical_Operator_out9186_out1;

  Logical_Operator_out9955_out1 <= Logical_Operator_out8931_out1 XOR Logical_Operator_out9187_out1;

  Logical_Operator_out9956_out1 <= Logical_Operator_out8932_out1 XOR Logical_Operator_out9188_out1;

  Logical_Operator_out9957_out1 <= Logical_Operator_out8933_out1 XOR Logical_Operator_out9189_out1;

  Logical_Operator_out9958_out1 <= Logical_Operator_out8934_out1 XOR Logical_Operator_out9190_out1;

  Logical_Operator_out9959_out1 <= Logical_Operator_out8935_out1 XOR Logical_Operator_out9191_out1;

  Logical_Operator_out9960_out1 <= Logical_Operator_out8936_out1 XOR Logical_Operator_out9192_out1;

  Logical_Operator_out9961_out1 <= Logical_Operator_out8937_out1 XOR Logical_Operator_out9193_out1;

  Logical_Operator_out9962_out1 <= Logical_Operator_out8938_out1 XOR Logical_Operator_out9194_out1;

  Logical_Operator_out9963_out1 <= Logical_Operator_out8939_out1 XOR Logical_Operator_out9195_out1;

  Logical_Operator_out9964_out1 <= Logical_Operator_out8940_out1 XOR Logical_Operator_out9196_out1;

  Logical_Operator_out9965_out1 <= Logical_Operator_out8941_out1 XOR Logical_Operator_out9197_out1;

  Logical_Operator_out9966_out1 <= Logical_Operator_out8942_out1 XOR Logical_Operator_out9198_out1;

  Logical_Operator_out9967_out1 <= Logical_Operator_out8943_out1 XOR Logical_Operator_out9199_out1;

  Logical_Operator_out9968_out1 <= Logical_Operator_out8944_out1 XOR Logical_Operator_out9200_out1;

  Logical_Operator_out9969_out1 <= Logical_Operator_out8945_out1 XOR Logical_Operator_out9201_out1;

  Logical_Operator_out9970_out1 <= Logical_Operator_out8946_out1 XOR Logical_Operator_out9202_out1;

  Logical_Operator_out9971_out1 <= Logical_Operator_out8947_out1 XOR Logical_Operator_out9203_out1;

  Logical_Operator_out9972_out1 <= Logical_Operator_out8948_out1 XOR Logical_Operator_out9204_out1;

  Logical_Operator_out9973_out1 <= Logical_Operator_out8949_out1 XOR Logical_Operator_out9205_out1;

  Logical_Operator_out9974_out1 <= Logical_Operator_out8950_out1 XOR Logical_Operator_out9206_out1;

  Logical_Operator_out9975_out1 <= Logical_Operator_out8951_out1 XOR Logical_Operator_out9207_out1;

  Logical_Operator_out9976_out1 <= Logical_Operator_out8952_out1 XOR Logical_Operator_out9208_out1;

  Logical_Operator_out9977_out1 <= Logical_Operator_out8953_out1 XOR Logical_Operator_out9209_out1;

  Logical_Operator_out9978_out1 <= Logical_Operator_out8954_out1 XOR Logical_Operator_out9210_out1;

  Logical_Operator_out9979_out1 <= Logical_Operator_out8955_out1 XOR Logical_Operator_out9211_out1;

  Logical_Operator_out9980_out1 <= Logical_Operator_out8956_out1 XOR Logical_Operator_out9212_out1;

  Logical_Operator_out9981_out1 <= Logical_Operator_out8957_out1 XOR Logical_Operator_out9213_out1;

  Logical_Operator_out9982_out1 <= Logical_Operator_out8958_out1 XOR Logical_Operator_out9214_out1;

  Logical_Operator_out9983_out1 <= Logical_Operator_out8959_out1 XOR Logical_Operator_out9215_out1;

  Logical_Operator_out9984_out1 <= Logical_Operator_out8960_out1 XOR Logical_Operator_out9216_out1;

  Logical_Operator_out9985_out1 <= Logical_Operator_out7809_out1 XOR Logical_Operator_out8065_out1;

  Logical_Operator_out9986_out1 <= Logical_Operator_out7810_out1 XOR Logical_Operator_out8066_out1;

  Logical_Operator_out9987_out1 <= Logical_Operator_out7811_out1 XOR Logical_Operator_out8067_out1;

  Logical_Operator_out9988_out1 <= Logical_Operator_out7812_out1 XOR Logical_Operator_out8068_out1;

  Logical_Operator_out9989_out1 <= Logical_Operator_out7813_out1 XOR Logical_Operator_out8069_out1;

  Logical_Operator_out9990_out1 <= Logical_Operator_out7814_out1 XOR Logical_Operator_out8070_out1;

  Logical_Operator_out9991_out1 <= Logical_Operator_out7815_out1 XOR Logical_Operator_out8071_out1;

  Logical_Operator_out9992_out1 <= Logical_Operator_out7816_out1 XOR Logical_Operator_out8072_out1;

  Logical_Operator_out9993_out1 <= Logical_Operator_out7817_out1 XOR Logical_Operator_out8073_out1;

  Logical_Operator_out9994_out1 <= Logical_Operator_out7818_out1 XOR Logical_Operator_out8074_out1;

  Logical_Operator_out9995_out1 <= Logical_Operator_out7819_out1 XOR Logical_Operator_out8075_out1;

  Logical_Operator_out9996_out1 <= Logical_Operator_out7820_out1 XOR Logical_Operator_out8076_out1;

  Logical_Operator_out9997_out1 <= Logical_Operator_out7821_out1 XOR Logical_Operator_out8077_out1;

  Logical_Operator_out9998_out1 <= Logical_Operator_out7822_out1 XOR Logical_Operator_out8078_out1;

  Logical_Operator_out9999_out1 <= Logical_Operator_out7823_out1 XOR Logical_Operator_out8079_out1;

  Logical_Operator_out10000_out1 <= Logical_Operator_out7824_out1 XOR Logical_Operator_out8080_out1;

  Logical_Operator_out10001_out1 <= Logical_Operator_out7825_out1 XOR Logical_Operator_out8081_out1;

  Logical_Operator_out10002_out1 <= Logical_Operator_out7826_out1 XOR Logical_Operator_out8082_out1;

  Logical_Operator_out10003_out1 <= Logical_Operator_out7827_out1 XOR Logical_Operator_out8083_out1;

  Logical_Operator_out10004_out1 <= Logical_Operator_out7828_out1 XOR Logical_Operator_out8084_out1;

  Logical_Operator_out10005_out1 <= Logical_Operator_out7829_out1 XOR Logical_Operator_out8085_out1;

  Logical_Operator_out10006_out1 <= Logical_Operator_out7830_out1 XOR Logical_Operator_out8086_out1;

  Logical_Operator_out10007_out1 <= Logical_Operator_out7831_out1 XOR Logical_Operator_out8087_out1;

  Logical_Operator_out10008_out1 <= Logical_Operator_out7832_out1 XOR Logical_Operator_out8088_out1;

  Logical_Operator_out10009_out1 <= Logical_Operator_out7833_out1 XOR Logical_Operator_out8089_out1;

  Logical_Operator_out10010_out1 <= Logical_Operator_out7834_out1 XOR Logical_Operator_out8090_out1;

  Logical_Operator_out10011_out1 <= Logical_Operator_out7835_out1 XOR Logical_Operator_out8091_out1;

  Logical_Operator_out10012_out1 <= Logical_Operator_out7836_out1 XOR Logical_Operator_out8092_out1;

  Logical_Operator_out10013_out1 <= Logical_Operator_out7837_out1 XOR Logical_Operator_out8093_out1;

  Logical_Operator_out10014_out1 <= Logical_Operator_out7838_out1 XOR Logical_Operator_out8094_out1;

  Logical_Operator_out10015_out1 <= Logical_Operator_out7839_out1 XOR Logical_Operator_out8095_out1;

  Logical_Operator_out10016_out1 <= Logical_Operator_out7840_out1 XOR Logical_Operator_out8096_out1;

  Logical_Operator_out10017_out1 <= Logical_Operator_out7841_out1 XOR Logical_Operator_out8097_out1;

  Logical_Operator_out10018_out1 <= Logical_Operator_out7842_out1 XOR Logical_Operator_out8098_out1;

  Logical_Operator_out10019_out1 <= Logical_Operator_out7843_out1 XOR Logical_Operator_out8099_out1;

  Logical_Operator_out10020_out1 <= Logical_Operator_out7844_out1 XOR Logical_Operator_out8100_out1;

  Logical_Operator_out10021_out1 <= Logical_Operator_out7845_out1 XOR Logical_Operator_out8101_out1;

  Logical_Operator_out10022_out1 <= Logical_Operator_out7846_out1 XOR Logical_Operator_out8102_out1;

  Logical_Operator_out10023_out1 <= Logical_Operator_out7847_out1 XOR Logical_Operator_out8103_out1;

  Logical_Operator_out10024_out1 <= Logical_Operator_out7848_out1 XOR Logical_Operator_out8104_out1;

  Logical_Operator_out10025_out1 <= Logical_Operator_out7849_out1 XOR Logical_Operator_out8105_out1;

  Logical_Operator_out10026_out1 <= Logical_Operator_out7850_out1 XOR Logical_Operator_out8106_out1;

  Logical_Operator_out10027_out1 <= Logical_Operator_out7851_out1 XOR Logical_Operator_out8107_out1;

  Logical_Operator_out10028_out1 <= Logical_Operator_out7852_out1 XOR Logical_Operator_out8108_out1;

  Logical_Operator_out10029_out1 <= Logical_Operator_out7853_out1 XOR Logical_Operator_out8109_out1;

  Logical_Operator_out10030_out1 <= Logical_Operator_out7854_out1 XOR Logical_Operator_out8110_out1;

  Logical_Operator_out10031_out1 <= Logical_Operator_out7855_out1 XOR Logical_Operator_out8111_out1;

  Logical_Operator_out10032_out1 <= Logical_Operator_out7856_out1 XOR Logical_Operator_out8112_out1;

  Logical_Operator_out10033_out1 <= Logical_Operator_out7857_out1 XOR Logical_Operator_out8113_out1;

  Logical_Operator_out10034_out1 <= Logical_Operator_out7858_out1 XOR Logical_Operator_out8114_out1;

  Logical_Operator_out10035_out1 <= Logical_Operator_out7859_out1 XOR Logical_Operator_out8115_out1;

  Logical_Operator_out10036_out1 <= Logical_Operator_out7860_out1 XOR Logical_Operator_out8116_out1;

  Logical_Operator_out10037_out1 <= Logical_Operator_out7861_out1 XOR Logical_Operator_out8117_out1;

  Logical_Operator_out10038_out1 <= Logical_Operator_out7862_out1 XOR Logical_Operator_out8118_out1;

  Logical_Operator_out10039_out1 <= Logical_Operator_out7863_out1 XOR Logical_Operator_out8119_out1;

  Logical_Operator_out10040_out1 <= Logical_Operator_out7864_out1 XOR Logical_Operator_out8120_out1;

  Logical_Operator_out10041_out1 <= Logical_Operator_out7865_out1 XOR Logical_Operator_out8121_out1;

  Logical_Operator_out10042_out1 <= Logical_Operator_out7866_out1 XOR Logical_Operator_out8122_out1;

  Logical_Operator_out10043_out1 <= Logical_Operator_out7867_out1 XOR Logical_Operator_out8123_out1;

  Logical_Operator_out10044_out1 <= Logical_Operator_out7868_out1 XOR Logical_Operator_out8124_out1;

  Logical_Operator_out10045_out1 <= Logical_Operator_out7869_out1 XOR Logical_Operator_out8125_out1;

  Logical_Operator_out10046_out1 <= Logical_Operator_out7870_out1 XOR Logical_Operator_out8126_out1;

  Logical_Operator_out10047_out1 <= Logical_Operator_out7871_out1 XOR Logical_Operator_out8127_out1;

  Logical_Operator_out10048_out1 <= Logical_Operator_out7872_out1 XOR Logical_Operator_out8128_out1;

  Logical_Operator_out10049_out1 <= Logical_Operator_out7873_out1 XOR Logical_Operator_out8129_out1;

  Logical_Operator_out10050_out1 <= Logical_Operator_out7874_out1 XOR Logical_Operator_out8130_out1;

  Logical_Operator_out10051_out1 <= Logical_Operator_out7875_out1 XOR Logical_Operator_out8131_out1;

  Logical_Operator_out10052_out1 <= Logical_Operator_out7876_out1 XOR Logical_Operator_out8132_out1;

  Logical_Operator_out10053_out1 <= Logical_Operator_out7877_out1 XOR Logical_Operator_out8133_out1;

  Logical_Operator_out10054_out1 <= Logical_Operator_out7878_out1 XOR Logical_Operator_out8134_out1;

  Logical_Operator_out10055_out1 <= Logical_Operator_out7879_out1 XOR Logical_Operator_out8135_out1;

  Logical_Operator_out10056_out1 <= Logical_Operator_out7880_out1 XOR Logical_Operator_out8136_out1;

  Logical_Operator_out10057_out1 <= Logical_Operator_out7881_out1 XOR Logical_Operator_out8137_out1;

  Logical_Operator_out10058_out1 <= Logical_Operator_out7882_out1 XOR Logical_Operator_out8138_out1;

  Logical_Operator_out10059_out1 <= Logical_Operator_out7883_out1 XOR Logical_Operator_out8139_out1;

  Logical_Operator_out10060_out1 <= Logical_Operator_out7884_out1 XOR Logical_Operator_out8140_out1;

  Logical_Operator_out10061_out1 <= Logical_Operator_out7885_out1 XOR Logical_Operator_out8141_out1;

  Logical_Operator_out10062_out1 <= Logical_Operator_out7886_out1 XOR Logical_Operator_out8142_out1;

  Logical_Operator_out10063_out1 <= Logical_Operator_out7887_out1 XOR Logical_Operator_out8143_out1;

  Logical_Operator_out10064_out1 <= Logical_Operator_out7888_out1 XOR Logical_Operator_out8144_out1;

  Logical_Operator_out10065_out1 <= Logical_Operator_out7889_out1 XOR Logical_Operator_out8145_out1;

  Logical_Operator_out10066_out1 <= Logical_Operator_out7890_out1 XOR Logical_Operator_out8146_out1;

  Logical_Operator_out10067_out1 <= Logical_Operator_out7891_out1 XOR Logical_Operator_out8147_out1;

  Logical_Operator_out10068_out1 <= Logical_Operator_out7892_out1 XOR Logical_Operator_out8148_out1;

  Logical_Operator_out10069_out1 <= Logical_Operator_out7893_out1 XOR Logical_Operator_out8149_out1;

  Logical_Operator_out10070_out1 <= Logical_Operator_out7894_out1 XOR Logical_Operator_out8150_out1;

  Logical_Operator_out10071_out1 <= Logical_Operator_out7895_out1 XOR Logical_Operator_out8151_out1;

  Logical_Operator_out10072_out1 <= Logical_Operator_out7896_out1 XOR Logical_Operator_out8152_out1;

  Logical_Operator_out10073_out1 <= Logical_Operator_out7897_out1 XOR Logical_Operator_out8153_out1;

  Logical_Operator_out10074_out1 <= Logical_Operator_out7898_out1 XOR Logical_Operator_out8154_out1;

  Logical_Operator_out10075_out1 <= Logical_Operator_out7899_out1 XOR Logical_Operator_out8155_out1;

  Logical_Operator_out10076_out1 <= Logical_Operator_out7900_out1 XOR Logical_Operator_out8156_out1;

  Logical_Operator_out10077_out1 <= Logical_Operator_out7901_out1 XOR Logical_Operator_out8157_out1;

  Logical_Operator_out10078_out1 <= Logical_Operator_out7902_out1 XOR Logical_Operator_out8158_out1;

  Logical_Operator_out10079_out1 <= Logical_Operator_out7903_out1 XOR Logical_Operator_out8159_out1;

  Logical_Operator_out10080_out1 <= Logical_Operator_out7904_out1 XOR Logical_Operator_out8160_out1;

  Logical_Operator_out10081_out1 <= Logical_Operator_out7905_out1 XOR Logical_Operator_out8161_out1;

  Logical_Operator_out10082_out1 <= Logical_Operator_out7906_out1 XOR Logical_Operator_out8162_out1;

  Logical_Operator_out10083_out1 <= Logical_Operator_out7907_out1 XOR Logical_Operator_out8163_out1;

  Logical_Operator_out10084_out1 <= Logical_Operator_out7908_out1 XOR Logical_Operator_out8164_out1;

  Logical_Operator_out10085_out1 <= Logical_Operator_out7909_out1 XOR Logical_Operator_out8165_out1;

  Logical_Operator_out10086_out1 <= Logical_Operator_out7910_out1 XOR Logical_Operator_out8166_out1;

  Logical_Operator_out10087_out1 <= Logical_Operator_out7911_out1 XOR Logical_Operator_out8167_out1;

  Logical_Operator_out10088_out1 <= Logical_Operator_out7912_out1 XOR Logical_Operator_out8168_out1;

  Logical_Operator_out10089_out1 <= Logical_Operator_out7913_out1 XOR Logical_Operator_out8169_out1;

  Logical_Operator_out10090_out1 <= Logical_Operator_out7914_out1 XOR Logical_Operator_out8170_out1;

  Logical_Operator_out10091_out1 <= Logical_Operator_out7915_out1 XOR Logical_Operator_out8171_out1;

  Logical_Operator_out10092_out1 <= Logical_Operator_out7916_out1 XOR Logical_Operator_out8172_out1;

  Logical_Operator_out10093_out1 <= Logical_Operator_out7917_out1 XOR Logical_Operator_out8173_out1;

  Logical_Operator_out10094_out1 <= Logical_Operator_out7918_out1 XOR Logical_Operator_out8174_out1;

  Logical_Operator_out10095_out1 <= Logical_Operator_out7919_out1 XOR Logical_Operator_out8175_out1;

  Logical_Operator_out10096_out1 <= Logical_Operator_out7920_out1 XOR Logical_Operator_out8176_out1;

  Logical_Operator_out10097_out1 <= Logical_Operator_out7921_out1 XOR Logical_Operator_out8177_out1;

  Logical_Operator_out10098_out1 <= Logical_Operator_out7922_out1 XOR Logical_Operator_out8178_out1;

  Logical_Operator_out10099_out1 <= Logical_Operator_out7923_out1 XOR Logical_Operator_out8179_out1;

  Logical_Operator_out10100_out1 <= Logical_Operator_out7924_out1 XOR Logical_Operator_out8180_out1;

  Logical_Operator_out10101_out1 <= Logical_Operator_out7925_out1 XOR Logical_Operator_out8181_out1;

  Logical_Operator_out10102_out1 <= Logical_Operator_out7926_out1 XOR Logical_Operator_out8182_out1;

  Logical_Operator_out10103_out1 <= Logical_Operator_out7927_out1 XOR Logical_Operator_out8183_out1;

  Logical_Operator_out10104_out1 <= Logical_Operator_out7928_out1 XOR Logical_Operator_out8184_out1;

  Logical_Operator_out10105_out1 <= Logical_Operator_out7929_out1 XOR Logical_Operator_out8185_out1;

  Logical_Operator_out10106_out1 <= Logical_Operator_out7930_out1 XOR Logical_Operator_out8186_out1;

  Logical_Operator_out10107_out1 <= Logical_Operator_out7931_out1 XOR Logical_Operator_out8187_out1;

  Logical_Operator_out10108_out1 <= Logical_Operator_out7932_out1 XOR Logical_Operator_out8188_out1;

  Logical_Operator_out10109_out1 <= Logical_Operator_out7933_out1 XOR Logical_Operator_out8189_out1;

  Logical_Operator_out10110_out1 <= Logical_Operator_out7934_out1 XOR Logical_Operator_out8190_out1;

  Logical_Operator_out10111_out1 <= Logical_Operator_out7935_out1 XOR Logical_Operator_out8191_out1;

  Logical_Operator_out10112_out1 <= Logical_Operator_out7936_out1 XOR Logical_Operator_out8192_out1;

  Logical_Operator_out10113_out1 <= Logical_Operator_out6849_out1 XOR Logical_Operator_out7105_out1;

  Logical_Operator_out10114_out1 <= Logical_Operator_out6850_out1 XOR Logical_Operator_out7106_out1;

  Logical_Operator_out10115_out1 <= Logical_Operator_out6851_out1 XOR Logical_Operator_out7107_out1;

  Logical_Operator_out10116_out1 <= Logical_Operator_out6852_out1 XOR Logical_Operator_out7108_out1;

  Logical_Operator_out10117_out1 <= Logical_Operator_out6853_out1 XOR Logical_Operator_out7109_out1;

  Logical_Operator_out10118_out1 <= Logical_Operator_out6854_out1 XOR Logical_Operator_out7110_out1;

  Logical_Operator_out10119_out1 <= Logical_Operator_out6855_out1 XOR Logical_Operator_out7111_out1;

  Logical_Operator_out10120_out1 <= Logical_Operator_out6856_out1 XOR Logical_Operator_out7112_out1;

  Logical_Operator_out10121_out1 <= Logical_Operator_out6857_out1 XOR Logical_Operator_out7113_out1;

  Logical_Operator_out10122_out1 <= Logical_Operator_out6858_out1 XOR Logical_Operator_out7114_out1;

  Logical_Operator_out10123_out1 <= Logical_Operator_out6859_out1 XOR Logical_Operator_out7115_out1;

  Logical_Operator_out10124_out1 <= Logical_Operator_out6860_out1 XOR Logical_Operator_out7116_out1;

  Logical_Operator_out10125_out1 <= Logical_Operator_out6861_out1 XOR Logical_Operator_out7117_out1;

  Logical_Operator_out10126_out1 <= Logical_Operator_out6862_out1 XOR Logical_Operator_out7118_out1;

  Logical_Operator_out10127_out1 <= Logical_Operator_out6863_out1 XOR Logical_Operator_out7119_out1;

  Logical_Operator_out10128_out1 <= Logical_Operator_out6864_out1 XOR Logical_Operator_out7120_out1;

  Logical_Operator_out10129_out1 <= Logical_Operator_out6865_out1 XOR Logical_Operator_out7121_out1;

  Logical_Operator_out10130_out1 <= Logical_Operator_out6866_out1 XOR Logical_Operator_out7122_out1;

  Logical_Operator_out10131_out1 <= Logical_Operator_out6867_out1 XOR Logical_Operator_out7123_out1;

  Logical_Operator_out10132_out1 <= Logical_Operator_out6868_out1 XOR Logical_Operator_out7124_out1;

  Logical_Operator_out10133_out1 <= Logical_Operator_out6869_out1 XOR Logical_Operator_out7125_out1;

  Logical_Operator_out10134_out1 <= Logical_Operator_out6870_out1 XOR Logical_Operator_out7126_out1;

  Logical_Operator_out10135_out1 <= Logical_Operator_out6871_out1 XOR Logical_Operator_out7127_out1;

  Logical_Operator_out10136_out1 <= Logical_Operator_out6872_out1 XOR Logical_Operator_out7128_out1;

  Logical_Operator_out10137_out1 <= Logical_Operator_out6873_out1 XOR Logical_Operator_out7129_out1;

  Logical_Operator_out10138_out1 <= Logical_Operator_out6874_out1 XOR Logical_Operator_out7130_out1;

  Logical_Operator_out10139_out1 <= Logical_Operator_out6875_out1 XOR Logical_Operator_out7131_out1;

  Logical_Operator_out10140_out1 <= Logical_Operator_out6876_out1 XOR Logical_Operator_out7132_out1;

  Logical_Operator_out10141_out1 <= Logical_Operator_out6877_out1 XOR Logical_Operator_out7133_out1;

  Logical_Operator_out10142_out1 <= Logical_Operator_out6878_out1 XOR Logical_Operator_out7134_out1;

  Logical_Operator_out10143_out1 <= Logical_Operator_out6879_out1 XOR Logical_Operator_out7135_out1;

  Logical_Operator_out10144_out1 <= Logical_Operator_out6880_out1 XOR Logical_Operator_out7136_out1;

  Logical_Operator_out10145_out1 <= Logical_Operator_out6881_out1 XOR Logical_Operator_out7137_out1;

  Logical_Operator_out10146_out1 <= Logical_Operator_out6882_out1 XOR Logical_Operator_out7138_out1;

  Logical_Operator_out10147_out1 <= Logical_Operator_out6883_out1 XOR Logical_Operator_out7139_out1;

  Logical_Operator_out10148_out1 <= Logical_Operator_out6884_out1 XOR Logical_Operator_out7140_out1;

  Logical_Operator_out10149_out1 <= Logical_Operator_out6885_out1 XOR Logical_Operator_out7141_out1;

  Logical_Operator_out10150_out1 <= Logical_Operator_out6886_out1 XOR Logical_Operator_out7142_out1;

  Logical_Operator_out10151_out1 <= Logical_Operator_out6887_out1 XOR Logical_Operator_out7143_out1;

  Logical_Operator_out10152_out1 <= Logical_Operator_out6888_out1 XOR Logical_Operator_out7144_out1;

  Logical_Operator_out10153_out1 <= Logical_Operator_out6889_out1 XOR Logical_Operator_out7145_out1;

  Logical_Operator_out10154_out1 <= Logical_Operator_out6890_out1 XOR Logical_Operator_out7146_out1;

  Logical_Operator_out10155_out1 <= Logical_Operator_out6891_out1 XOR Logical_Operator_out7147_out1;

  Logical_Operator_out10156_out1 <= Logical_Operator_out6892_out1 XOR Logical_Operator_out7148_out1;

  Logical_Operator_out10157_out1 <= Logical_Operator_out6893_out1 XOR Logical_Operator_out7149_out1;

  Logical_Operator_out10158_out1 <= Logical_Operator_out6894_out1 XOR Logical_Operator_out7150_out1;

  Logical_Operator_out10159_out1 <= Logical_Operator_out6895_out1 XOR Logical_Operator_out7151_out1;

  Logical_Operator_out10160_out1 <= Logical_Operator_out6896_out1 XOR Logical_Operator_out7152_out1;

  Logical_Operator_out10161_out1 <= Logical_Operator_out6897_out1 XOR Logical_Operator_out7153_out1;

  Logical_Operator_out10162_out1 <= Logical_Operator_out6898_out1 XOR Logical_Operator_out7154_out1;

  Logical_Operator_out10163_out1 <= Logical_Operator_out6899_out1 XOR Logical_Operator_out7155_out1;

  Logical_Operator_out10164_out1 <= Logical_Operator_out6900_out1 XOR Logical_Operator_out7156_out1;

  Logical_Operator_out10165_out1 <= Logical_Operator_out6901_out1 XOR Logical_Operator_out7157_out1;

  Logical_Operator_out10166_out1 <= Logical_Operator_out6902_out1 XOR Logical_Operator_out7158_out1;

  Logical_Operator_out10167_out1 <= Logical_Operator_out6903_out1 XOR Logical_Operator_out7159_out1;

  Logical_Operator_out10168_out1 <= Logical_Operator_out6904_out1 XOR Logical_Operator_out7160_out1;

  Logical_Operator_out10169_out1 <= Logical_Operator_out6905_out1 XOR Logical_Operator_out7161_out1;

  Logical_Operator_out10170_out1 <= Logical_Operator_out6906_out1 XOR Logical_Operator_out7162_out1;

  Logical_Operator_out10171_out1 <= Logical_Operator_out6907_out1 XOR Logical_Operator_out7163_out1;

  Logical_Operator_out10172_out1 <= Logical_Operator_out6908_out1 XOR Logical_Operator_out7164_out1;

  Logical_Operator_out10173_out1 <= Logical_Operator_out6909_out1 XOR Logical_Operator_out7165_out1;

  Logical_Operator_out10174_out1 <= Logical_Operator_out6910_out1 XOR Logical_Operator_out7166_out1;

  Logical_Operator_out10175_out1 <= Logical_Operator_out6911_out1 XOR Logical_Operator_out7167_out1;

  Logical_Operator_out10176_out1 <= Logical_Operator_out6912_out1 XOR Logical_Operator_out7168_out1;

  Logical_Operator_out10177_out1 <= Logical_Operator_out5857_out1 XOR Logical_Operator_out6113_out1;

  Logical_Operator_out10178_out1 <= Logical_Operator_out5858_out1 XOR Logical_Operator_out6114_out1;

  Logical_Operator_out10179_out1 <= Logical_Operator_out5859_out1 XOR Logical_Operator_out6115_out1;

  Logical_Operator_out10180_out1 <= Logical_Operator_out5860_out1 XOR Logical_Operator_out6116_out1;

  Logical_Operator_out10181_out1 <= Logical_Operator_out5861_out1 XOR Logical_Operator_out6117_out1;

  Logical_Operator_out10182_out1 <= Logical_Operator_out5862_out1 XOR Logical_Operator_out6118_out1;

  Logical_Operator_out10183_out1 <= Logical_Operator_out5863_out1 XOR Logical_Operator_out6119_out1;

  Logical_Operator_out10184_out1 <= Logical_Operator_out5864_out1 XOR Logical_Operator_out6120_out1;

  Logical_Operator_out10185_out1 <= Logical_Operator_out5865_out1 XOR Logical_Operator_out6121_out1;

  Logical_Operator_out10186_out1 <= Logical_Operator_out5866_out1 XOR Logical_Operator_out6122_out1;

  Logical_Operator_out10187_out1 <= Logical_Operator_out5867_out1 XOR Logical_Operator_out6123_out1;

  Logical_Operator_out10188_out1 <= Logical_Operator_out5868_out1 XOR Logical_Operator_out6124_out1;

  Logical_Operator_out10189_out1 <= Logical_Operator_out5869_out1 XOR Logical_Operator_out6125_out1;

  Logical_Operator_out10190_out1 <= Logical_Operator_out5870_out1 XOR Logical_Operator_out6126_out1;

  Logical_Operator_out10191_out1 <= Logical_Operator_out5871_out1 XOR Logical_Operator_out6127_out1;

  Logical_Operator_out10192_out1 <= Logical_Operator_out5872_out1 XOR Logical_Operator_out6128_out1;

  Logical_Operator_out10193_out1 <= Logical_Operator_out5873_out1 XOR Logical_Operator_out6129_out1;

  Logical_Operator_out10194_out1 <= Logical_Operator_out5874_out1 XOR Logical_Operator_out6130_out1;

  Logical_Operator_out10195_out1 <= Logical_Operator_out5875_out1 XOR Logical_Operator_out6131_out1;

  Logical_Operator_out10196_out1 <= Logical_Operator_out5876_out1 XOR Logical_Operator_out6132_out1;

  Logical_Operator_out10197_out1 <= Logical_Operator_out5877_out1 XOR Logical_Operator_out6133_out1;

  Logical_Operator_out10198_out1 <= Logical_Operator_out5878_out1 XOR Logical_Operator_out6134_out1;

  Logical_Operator_out10199_out1 <= Logical_Operator_out5879_out1 XOR Logical_Operator_out6135_out1;

  Logical_Operator_out10200_out1 <= Logical_Operator_out5880_out1 XOR Logical_Operator_out6136_out1;

  Logical_Operator_out10201_out1 <= Logical_Operator_out5881_out1 XOR Logical_Operator_out6137_out1;

  Logical_Operator_out10202_out1 <= Logical_Operator_out5882_out1 XOR Logical_Operator_out6138_out1;

  Logical_Operator_out10203_out1 <= Logical_Operator_out5883_out1 XOR Logical_Operator_out6139_out1;

  Logical_Operator_out10204_out1 <= Logical_Operator_out5884_out1 XOR Logical_Operator_out6140_out1;

  Logical_Operator_out10205_out1 <= Logical_Operator_out5885_out1 XOR Logical_Operator_out6141_out1;

  Logical_Operator_out10206_out1 <= Logical_Operator_out5886_out1 XOR Logical_Operator_out6142_out1;

  Logical_Operator_out10207_out1 <= Logical_Operator_out5887_out1 XOR Logical_Operator_out6143_out1;

  Logical_Operator_out10208_out1 <= Logical_Operator_out5888_out1 XOR Logical_Operator_out6144_out1;

  Logical_Operator_out10209_out1 <= Logical_Operator_out4849_out1 XOR Logical_Operator_out5105_out1;

  Logical_Operator_out10210_out1 <= Logical_Operator_out4850_out1 XOR Logical_Operator_out5106_out1;

  Logical_Operator_out10211_out1 <= Logical_Operator_out4851_out1 XOR Logical_Operator_out5107_out1;

  Logical_Operator_out10212_out1 <= Logical_Operator_out4852_out1 XOR Logical_Operator_out5108_out1;

  Logical_Operator_out10213_out1 <= Logical_Operator_out4853_out1 XOR Logical_Operator_out5109_out1;

  Logical_Operator_out10214_out1 <= Logical_Operator_out4854_out1 XOR Logical_Operator_out5110_out1;

  Logical_Operator_out10215_out1 <= Logical_Operator_out4855_out1 XOR Logical_Operator_out5111_out1;

  Logical_Operator_out10216_out1 <= Logical_Operator_out4856_out1 XOR Logical_Operator_out5112_out1;

  Logical_Operator_out10217_out1 <= Logical_Operator_out4857_out1 XOR Logical_Operator_out5113_out1;

  Logical_Operator_out10218_out1 <= Logical_Operator_out4858_out1 XOR Logical_Operator_out5114_out1;

  Logical_Operator_out10219_out1 <= Logical_Operator_out4859_out1 XOR Logical_Operator_out5115_out1;

  Logical_Operator_out10220_out1 <= Logical_Operator_out4860_out1 XOR Logical_Operator_out5116_out1;

  Logical_Operator_out10221_out1 <= Logical_Operator_out4861_out1 XOR Logical_Operator_out5117_out1;

  Logical_Operator_out10222_out1 <= Logical_Operator_out4862_out1 XOR Logical_Operator_out5118_out1;

  Logical_Operator_out10223_out1 <= Logical_Operator_out4863_out1 XOR Logical_Operator_out5119_out1;

  Logical_Operator_out10224_out1 <= Logical_Operator_out4864_out1 XOR Logical_Operator_out5120_out1;

  Logical_Operator_out10225_out1 <= Logical_Operator_out3833_out1 XOR Logical_Operator_out4089_out1;

  Logical_Operator_out10226_out1 <= Logical_Operator_out3834_out1 XOR Logical_Operator_out4090_out1;

  Logical_Operator_out10227_out1 <= Logical_Operator_out3835_out1 XOR Logical_Operator_out4091_out1;

  Logical_Operator_out10228_out1 <= Logical_Operator_out3836_out1 XOR Logical_Operator_out4092_out1;

  Logical_Operator_out10229_out1 <= Logical_Operator_out3837_out1 XOR Logical_Operator_out4093_out1;

  Logical_Operator_out10230_out1 <= Logical_Operator_out3838_out1 XOR Logical_Operator_out4094_out1;

  Logical_Operator_out10231_out1 <= Logical_Operator_out3839_out1 XOR Logical_Operator_out4095_out1;

  Logical_Operator_out10232_out1 <= Logical_Operator_out3840_out1 XOR Logical_Operator_out4096_out1;

  Logical_Operator_out10233_out1 <= Logical_Operator_out2813_out1 XOR Logical_Operator_out3069_out1;

  Logical_Operator_out10234_out1 <= Logical_Operator_out2814_out1 XOR Logical_Operator_out3070_out1;

  Logical_Operator_out10235_out1 <= Logical_Operator_out2815_out1 XOR Logical_Operator_out3071_out1;

  Logical_Operator_out10236_out1 <= Logical_Operator_out2816_out1 XOR Logical_Operator_out3072_out1;

  Logical_Operator_out10237_out1 <= Logical_Operator_out1791_out1 XOR Logical_Operator_out2047_out1;

  Logical_Operator_out10238_out1 <= Logical_Operator_out1792_out1 XOR Logical_Operator_out2048_out1;

  Logical_Operator_out10239_out1 <= Logical_Operator_out768_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out10240_out1 <= in1536 XOR in2048;

  Logical_Operator_out10241_out1 <= Logical_Operator_out9217_out1 XOR Logical_Operator_out9729_out1;

  Logical_Operator_out10242_out1 <= Logical_Operator_out9218_out1 XOR Logical_Operator_out9730_out1;

  Logical_Operator_out10243_out1 <= Logical_Operator_out9219_out1 XOR Logical_Operator_out9731_out1;

  Logical_Operator_out10244_out1 <= Logical_Operator_out9220_out1 XOR Logical_Operator_out9732_out1;

  Logical_Operator_out10245_out1 <= Logical_Operator_out9221_out1 XOR Logical_Operator_out9733_out1;

  Logical_Operator_out10246_out1 <= Logical_Operator_out9222_out1 XOR Logical_Operator_out9734_out1;

  Logical_Operator_out10247_out1 <= Logical_Operator_out9223_out1 XOR Logical_Operator_out9735_out1;

  Logical_Operator_out10248_out1 <= Logical_Operator_out9224_out1 XOR Logical_Operator_out9736_out1;

  Logical_Operator_out10249_out1 <= Logical_Operator_out9225_out1 XOR Logical_Operator_out9737_out1;

  Logical_Operator_out10250_out1 <= Logical_Operator_out9226_out1 XOR Logical_Operator_out9738_out1;

  Logical_Operator_out10251_out1 <= Logical_Operator_out9227_out1 XOR Logical_Operator_out9739_out1;

  Logical_Operator_out10252_out1 <= Logical_Operator_out9228_out1 XOR Logical_Operator_out9740_out1;

  Logical_Operator_out10253_out1 <= Logical_Operator_out9229_out1 XOR Logical_Operator_out9741_out1;

  Logical_Operator_out10254_out1 <= Logical_Operator_out9230_out1 XOR Logical_Operator_out9742_out1;

  Logical_Operator_out10255_out1 <= Logical_Operator_out9231_out1 XOR Logical_Operator_out9743_out1;

  Logical_Operator_out10256_out1 <= Logical_Operator_out9232_out1 XOR Logical_Operator_out9744_out1;

  Logical_Operator_out10257_out1 <= Logical_Operator_out9233_out1 XOR Logical_Operator_out9745_out1;

  Logical_Operator_out10258_out1 <= Logical_Operator_out9234_out1 XOR Logical_Operator_out9746_out1;

  Logical_Operator_out10259_out1 <= Logical_Operator_out9235_out1 XOR Logical_Operator_out9747_out1;

  Logical_Operator_out10260_out1 <= Logical_Operator_out9236_out1 XOR Logical_Operator_out9748_out1;

  Logical_Operator_out10261_out1 <= Logical_Operator_out9237_out1 XOR Logical_Operator_out9749_out1;

  Logical_Operator_out10262_out1 <= Logical_Operator_out9238_out1 XOR Logical_Operator_out9750_out1;

  Logical_Operator_out10263_out1 <= Logical_Operator_out9239_out1 XOR Logical_Operator_out9751_out1;

  Logical_Operator_out10264_out1 <= Logical_Operator_out9240_out1 XOR Logical_Operator_out9752_out1;

  Logical_Operator_out10265_out1 <= Logical_Operator_out9241_out1 XOR Logical_Operator_out9753_out1;

  Logical_Operator_out10266_out1 <= Logical_Operator_out9242_out1 XOR Logical_Operator_out9754_out1;

  Logical_Operator_out10267_out1 <= Logical_Operator_out9243_out1 XOR Logical_Operator_out9755_out1;

  Logical_Operator_out10268_out1 <= Logical_Operator_out9244_out1 XOR Logical_Operator_out9756_out1;

  Logical_Operator_out10269_out1 <= Logical_Operator_out9245_out1 XOR Logical_Operator_out9757_out1;

  Logical_Operator_out10270_out1 <= Logical_Operator_out9246_out1 XOR Logical_Operator_out9758_out1;

  Logical_Operator_out10271_out1 <= Logical_Operator_out9247_out1 XOR Logical_Operator_out9759_out1;

  Logical_Operator_out10272_out1 <= Logical_Operator_out9248_out1 XOR Logical_Operator_out9760_out1;

  Logical_Operator_out10273_out1 <= Logical_Operator_out9249_out1 XOR Logical_Operator_out9761_out1;

  Logical_Operator_out10274_out1 <= Logical_Operator_out9250_out1 XOR Logical_Operator_out9762_out1;

  Logical_Operator_out10275_out1 <= Logical_Operator_out9251_out1 XOR Logical_Operator_out9763_out1;

  Logical_Operator_out10276_out1 <= Logical_Operator_out9252_out1 XOR Logical_Operator_out9764_out1;

  Logical_Operator_out10277_out1 <= Logical_Operator_out9253_out1 XOR Logical_Operator_out9765_out1;

  Logical_Operator_out10278_out1 <= Logical_Operator_out9254_out1 XOR Logical_Operator_out9766_out1;

  Logical_Operator_out10279_out1 <= Logical_Operator_out9255_out1 XOR Logical_Operator_out9767_out1;

  Logical_Operator_out10280_out1 <= Logical_Operator_out9256_out1 XOR Logical_Operator_out9768_out1;

  Logical_Operator_out10281_out1 <= Logical_Operator_out9257_out1 XOR Logical_Operator_out9769_out1;

  Logical_Operator_out10282_out1 <= Logical_Operator_out9258_out1 XOR Logical_Operator_out9770_out1;

  Logical_Operator_out10283_out1 <= Logical_Operator_out9259_out1 XOR Logical_Operator_out9771_out1;

  Logical_Operator_out10284_out1 <= Logical_Operator_out9260_out1 XOR Logical_Operator_out9772_out1;

  Logical_Operator_out10285_out1 <= Logical_Operator_out9261_out1 XOR Logical_Operator_out9773_out1;

  Logical_Operator_out10286_out1 <= Logical_Operator_out9262_out1 XOR Logical_Operator_out9774_out1;

  Logical_Operator_out10287_out1 <= Logical_Operator_out9263_out1 XOR Logical_Operator_out9775_out1;

  Logical_Operator_out10288_out1 <= Logical_Operator_out9264_out1 XOR Logical_Operator_out9776_out1;

  Logical_Operator_out10289_out1 <= Logical_Operator_out9265_out1 XOR Logical_Operator_out9777_out1;

  Logical_Operator_out10290_out1 <= Logical_Operator_out9266_out1 XOR Logical_Operator_out9778_out1;

  Logical_Operator_out10291_out1 <= Logical_Operator_out9267_out1 XOR Logical_Operator_out9779_out1;

  Logical_Operator_out10292_out1 <= Logical_Operator_out9268_out1 XOR Logical_Operator_out9780_out1;

  Logical_Operator_out10293_out1 <= Logical_Operator_out9269_out1 XOR Logical_Operator_out9781_out1;

  Logical_Operator_out10294_out1 <= Logical_Operator_out9270_out1 XOR Logical_Operator_out9782_out1;

  Logical_Operator_out10295_out1 <= Logical_Operator_out9271_out1 XOR Logical_Operator_out9783_out1;

  Logical_Operator_out10296_out1 <= Logical_Operator_out9272_out1 XOR Logical_Operator_out9784_out1;

  Logical_Operator_out10297_out1 <= Logical_Operator_out9273_out1 XOR Logical_Operator_out9785_out1;

  Logical_Operator_out10298_out1 <= Logical_Operator_out9274_out1 XOR Logical_Operator_out9786_out1;

  Logical_Operator_out10299_out1 <= Logical_Operator_out9275_out1 XOR Logical_Operator_out9787_out1;

  Logical_Operator_out10300_out1 <= Logical_Operator_out9276_out1 XOR Logical_Operator_out9788_out1;

  Logical_Operator_out10301_out1 <= Logical_Operator_out9277_out1 XOR Logical_Operator_out9789_out1;

  Logical_Operator_out10302_out1 <= Logical_Operator_out9278_out1 XOR Logical_Operator_out9790_out1;

  Logical_Operator_out10303_out1 <= Logical_Operator_out9279_out1 XOR Logical_Operator_out9791_out1;

  Logical_Operator_out10304_out1 <= Logical_Operator_out9280_out1 XOR Logical_Operator_out9792_out1;

  Logical_Operator_out10305_out1 <= Logical_Operator_out9281_out1 XOR Logical_Operator_out9793_out1;

  Logical_Operator_out10306_out1 <= Logical_Operator_out9282_out1 XOR Logical_Operator_out9794_out1;

  Logical_Operator_out10307_out1 <= Logical_Operator_out9283_out1 XOR Logical_Operator_out9795_out1;

  Logical_Operator_out10308_out1 <= Logical_Operator_out9284_out1 XOR Logical_Operator_out9796_out1;

  Logical_Operator_out10309_out1 <= Logical_Operator_out9285_out1 XOR Logical_Operator_out9797_out1;

  Logical_Operator_out10310_out1 <= Logical_Operator_out9286_out1 XOR Logical_Operator_out9798_out1;

  Logical_Operator_out10311_out1 <= Logical_Operator_out9287_out1 XOR Logical_Operator_out9799_out1;

  Logical_Operator_out10312_out1 <= Logical_Operator_out9288_out1 XOR Logical_Operator_out9800_out1;

  Logical_Operator_out10313_out1 <= Logical_Operator_out9289_out1 XOR Logical_Operator_out9801_out1;

  Logical_Operator_out10314_out1 <= Logical_Operator_out9290_out1 XOR Logical_Operator_out9802_out1;

  Logical_Operator_out10315_out1 <= Logical_Operator_out9291_out1 XOR Logical_Operator_out9803_out1;

  Logical_Operator_out10316_out1 <= Logical_Operator_out9292_out1 XOR Logical_Operator_out9804_out1;

  Logical_Operator_out10317_out1 <= Logical_Operator_out9293_out1 XOR Logical_Operator_out9805_out1;

  Logical_Operator_out10318_out1 <= Logical_Operator_out9294_out1 XOR Logical_Operator_out9806_out1;

  Logical_Operator_out10319_out1 <= Logical_Operator_out9295_out1 XOR Logical_Operator_out9807_out1;

  Logical_Operator_out10320_out1 <= Logical_Operator_out9296_out1 XOR Logical_Operator_out9808_out1;

  Logical_Operator_out10321_out1 <= Logical_Operator_out9297_out1 XOR Logical_Operator_out9809_out1;

  Logical_Operator_out10322_out1 <= Logical_Operator_out9298_out1 XOR Logical_Operator_out9810_out1;

  Logical_Operator_out10323_out1 <= Logical_Operator_out9299_out1 XOR Logical_Operator_out9811_out1;

  Logical_Operator_out10324_out1 <= Logical_Operator_out9300_out1 XOR Logical_Operator_out9812_out1;

  Logical_Operator_out10325_out1 <= Logical_Operator_out9301_out1 XOR Logical_Operator_out9813_out1;

  Logical_Operator_out10326_out1 <= Logical_Operator_out9302_out1 XOR Logical_Operator_out9814_out1;

  Logical_Operator_out10327_out1 <= Logical_Operator_out9303_out1 XOR Logical_Operator_out9815_out1;

  Logical_Operator_out10328_out1 <= Logical_Operator_out9304_out1 XOR Logical_Operator_out9816_out1;

  Logical_Operator_out10329_out1 <= Logical_Operator_out9305_out1 XOR Logical_Operator_out9817_out1;

  Logical_Operator_out10330_out1 <= Logical_Operator_out9306_out1 XOR Logical_Operator_out9818_out1;

  Logical_Operator_out10331_out1 <= Logical_Operator_out9307_out1 XOR Logical_Operator_out9819_out1;

  Logical_Operator_out10332_out1 <= Logical_Operator_out9308_out1 XOR Logical_Operator_out9820_out1;

  Logical_Operator_out10333_out1 <= Logical_Operator_out9309_out1 XOR Logical_Operator_out9821_out1;

  Logical_Operator_out10334_out1 <= Logical_Operator_out9310_out1 XOR Logical_Operator_out9822_out1;

  Logical_Operator_out10335_out1 <= Logical_Operator_out9311_out1 XOR Logical_Operator_out9823_out1;

  Logical_Operator_out10336_out1 <= Logical_Operator_out9312_out1 XOR Logical_Operator_out9824_out1;

  Logical_Operator_out10337_out1 <= Logical_Operator_out9313_out1 XOR Logical_Operator_out9825_out1;

  Logical_Operator_out10338_out1 <= Logical_Operator_out9314_out1 XOR Logical_Operator_out9826_out1;

  Logical_Operator_out10339_out1 <= Logical_Operator_out9315_out1 XOR Logical_Operator_out9827_out1;

  Logical_Operator_out10340_out1 <= Logical_Operator_out9316_out1 XOR Logical_Operator_out9828_out1;

  Logical_Operator_out10341_out1 <= Logical_Operator_out9317_out1 XOR Logical_Operator_out9829_out1;

  Logical_Operator_out10342_out1 <= Logical_Operator_out9318_out1 XOR Logical_Operator_out9830_out1;

  Logical_Operator_out10343_out1 <= Logical_Operator_out9319_out1 XOR Logical_Operator_out9831_out1;

  Logical_Operator_out10344_out1 <= Logical_Operator_out9320_out1 XOR Logical_Operator_out9832_out1;

  Logical_Operator_out10345_out1 <= Logical_Operator_out9321_out1 XOR Logical_Operator_out9833_out1;

  Logical_Operator_out10346_out1 <= Logical_Operator_out9322_out1 XOR Logical_Operator_out9834_out1;

  Logical_Operator_out10347_out1 <= Logical_Operator_out9323_out1 XOR Logical_Operator_out9835_out1;

  Logical_Operator_out10348_out1 <= Logical_Operator_out9324_out1 XOR Logical_Operator_out9836_out1;

  Logical_Operator_out10349_out1 <= Logical_Operator_out9325_out1 XOR Logical_Operator_out9837_out1;

  Logical_Operator_out10350_out1 <= Logical_Operator_out9326_out1 XOR Logical_Operator_out9838_out1;

  Logical_Operator_out10351_out1 <= Logical_Operator_out9327_out1 XOR Logical_Operator_out9839_out1;

  Logical_Operator_out10352_out1 <= Logical_Operator_out9328_out1 XOR Logical_Operator_out9840_out1;

  Logical_Operator_out10353_out1 <= Logical_Operator_out9329_out1 XOR Logical_Operator_out9841_out1;

  Logical_Operator_out10354_out1 <= Logical_Operator_out9330_out1 XOR Logical_Operator_out9842_out1;

  Logical_Operator_out10355_out1 <= Logical_Operator_out9331_out1 XOR Logical_Operator_out9843_out1;

  Logical_Operator_out10356_out1 <= Logical_Operator_out9332_out1 XOR Logical_Operator_out9844_out1;

  Logical_Operator_out10357_out1 <= Logical_Operator_out9333_out1 XOR Logical_Operator_out9845_out1;

  Logical_Operator_out10358_out1 <= Logical_Operator_out9334_out1 XOR Logical_Operator_out9846_out1;

  Logical_Operator_out10359_out1 <= Logical_Operator_out9335_out1 XOR Logical_Operator_out9847_out1;

  Logical_Operator_out10360_out1 <= Logical_Operator_out9336_out1 XOR Logical_Operator_out9848_out1;

  Logical_Operator_out10361_out1 <= Logical_Operator_out9337_out1 XOR Logical_Operator_out9849_out1;

  Logical_Operator_out10362_out1 <= Logical_Operator_out9338_out1 XOR Logical_Operator_out9850_out1;

  Logical_Operator_out10363_out1 <= Logical_Operator_out9339_out1 XOR Logical_Operator_out9851_out1;

  Logical_Operator_out10364_out1 <= Logical_Operator_out9340_out1 XOR Logical_Operator_out9852_out1;

  Logical_Operator_out10365_out1 <= Logical_Operator_out9341_out1 XOR Logical_Operator_out9853_out1;

  Logical_Operator_out10366_out1 <= Logical_Operator_out9342_out1 XOR Logical_Operator_out9854_out1;

  Logical_Operator_out10367_out1 <= Logical_Operator_out9343_out1 XOR Logical_Operator_out9855_out1;

  Logical_Operator_out10368_out1 <= Logical_Operator_out9344_out1 XOR Logical_Operator_out9856_out1;

  Logical_Operator_out10369_out1 <= Logical_Operator_out9345_out1 XOR Logical_Operator_out9857_out1;

  Logical_Operator_out10370_out1 <= Logical_Operator_out9346_out1 XOR Logical_Operator_out9858_out1;

  Logical_Operator_out10371_out1 <= Logical_Operator_out9347_out1 XOR Logical_Operator_out9859_out1;

  Logical_Operator_out10372_out1 <= Logical_Operator_out9348_out1 XOR Logical_Operator_out9860_out1;

  Logical_Operator_out10373_out1 <= Logical_Operator_out9349_out1 XOR Logical_Operator_out9861_out1;

  Logical_Operator_out10374_out1 <= Logical_Operator_out9350_out1 XOR Logical_Operator_out9862_out1;

  Logical_Operator_out10375_out1 <= Logical_Operator_out9351_out1 XOR Logical_Operator_out9863_out1;

  Logical_Operator_out10376_out1 <= Logical_Operator_out9352_out1 XOR Logical_Operator_out9864_out1;

  Logical_Operator_out10377_out1 <= Logical_Operator_out9353_out1 XOR Logical_Operator_out9865_out1;

  Logical_Operator_out10378_out1 <= Logical_Operator_out9354_out1 XOR Logical_Operator_out9866_out1;

  Logical_Operator_out10379_out1 <= Logical_Operator_out9355_out1 XOR Logical_Operator_out9867_out1;

  Logical_Operator_out10380_out1 <= Logical_Operator_out9356_out1 XOR Logical_Operator_out9868_out1;

  Logical_Operator_out10381_out1 <= Logical_Operator_out9357_out1 XOR Logical_Operator_out9869_out1;

  Logical_Operator_out10382_out1 <= Logical_Operator_out9358_out1 XOR Logical_Operator_out9870_out1;

  Logical_Operator_out10383_out1 <= Logical_Operator_out9359_out1 XOR Logical_Operator_out9871_out1;

  Logical_Operator_out10384_out1 <= Logical_Operator_out9360_out1 XOR Logical_Operator_out9872_out1;

  Logical_Operator_out10385_out1 <= Logical_Operator_out9361_out1 XOR Logical_Operator_out9873_out1;

  Logical_Operator_out10386_out1 <= Logical_Operator_out9362_out1 XOR Logical_Operator_out9874_out1;

  Logical_Operator_out10387_out1 <= Logical_Operator_out9363_out1 XOR Logical_Operator_out9875_out1;

  Logical_Operator_out10388_out1 <= Logical_Operator_out9364_out1 XOR Logical_Operator_out9876_out1;

  Logical_Operator_out10389_out1 <= Logical_Operator_out9365_out1 XOR Logical_Operator_out9877_out1;

  Logical_Operator_out10390_out1 <= Logical_Operator_out9366_out1 XOR Logical_Operator_out9878_out1;

  Logical_Operator_out10391_out1 <= Logical_Operator_out9367_out1 XOR Logical_Operator_out9879_out1;

  Logical_Operator_out10392_out1 <= Logical_Operator_out9368_out1 XOR Logical_Operator_out9880_out1;

  Logical_Operator_out10393_out1 <= Logical_Operator_out9369_out1 XOR Logical_Operator_out9881_out1;

  Logical_Operator_out10394_out1 <= Logical_Operator_out9370_out1 XOR Logical_Operator_out9882_out1;

  Logical_Operator_out10395_out1 <= Logical_Operator_out9371_out1 XOR Logical_Operator_out9883_out1;

  Logical_Operator_out10396_out1 <= Logical_Operator_out9372_out1 XOR Logical_Operator_out9884_out1;

  Logical_Operator_out10397_out1 <= Logical_Operator_out9373_out1 XOR Logical_Operator_out9885_out1;

  Logical_Operator_out10398_out1 <= Logical_Operator_out9374_out1 XOR Logical_Operator_out9886_out1;

  Logical_Operator_out10399_out1 <= Logical_Operator_out9375_out1 XOR Logical_Operator_out9887_out1;

  Logical_Operator_out10400_out1 <= Logical_Operator_out9376_out1 XOR Logical_Operator_out9888_out1;

  Logical_Operator_out10401_out1 <= Logical_Operator_out9377_out1 XOR Logical_Operator_out9889_out1;

  Logical_Operator_out10402_out1 <= Logical_Operator_out9378_out1 XOR Logical_Operator_out9890_out1;

  Logical_Operator_out10403_out1 <= Logical_Operator_out9379_out1 XOR Logical_Operator_out9891_out1;

  Logical_Operator_out10404_out1 <= Logical_Operator_out9380_out1 XOR Logical_Operator_out9892_out1;

  Logical_Operator_out10405_out1 <= Logical_Operator_out9381_out1 XOR Logical_Operator_out9893_out1;

  Logical_Operator_out10406_out1 <= Logical_Operator_out9382_out1 XOR Logical_Operator_out9894_out1;

  Logical_Operator_out10407_out1 <= Logical_Operator_out9383_out1 XOR Logical_Operator_out9895_out1;

  Logical_Operator_out10408_out1 <= Logical_Operator_out9384_out1 XOR Logical_Operator_out9896_out1;

  Logical_Operator_out10409_out1 <= Logical_Operator_out9385_out1 XOR Logical_Operator_out9897_out1;

  Logical_Operator_out10410_out1 <= Logical_Operator_out9386_out1 XOR Logical_Operator_out9898_out1;

  Logical_Operator_out10411_out1 <= Logical_Operator_out9387_out1 XOR Logical_Operator_out9899_out1;

  Logical_Operator_out10412_out1 <= Logical_Operator_out9388_out1 XOR Logical_Operator_out9900_out1;

  Logical_Operator_out10413_out1 <= Logical_Operator_out9389_out1 XOR Logical_Operator_out9901_out1;

  Logical_Operator_out10414_out1 <= Logical_Operator_out9390_out1 XOR Logical_Operator_out9902_out1;

  Logical_Operator_out10415_out1 <= Logical_Operator_out9391_out1 XOR Logical_Operator_out9903_out1;

  Logical_Operator_out10416_out1 <= Logical_Operator_out9392_out1 XOR Logical_Operator_out9904_out1;

  Logical_Operator_out10417_out1 <= Logical_Operator_out9393_out1 XOR Logical_Operator_out9905_out1;

  Logical_Operator_out10418_out1 <= Logical_Operator_out9394_out1 XOR Logical_Operator_out9906_out1;

  Logical_Operator_out10419_out1 <= Logical_Operator_out9395_out1 XOR Logical_Operator_out9907_out1;

  Logical_Operator_out10420_out1 <= Logical_Operator_out9396_out1 XOR Logical_Operator_out9908_out1;

  Logical_Operator_out10421_out1 <= Logical_Operator_out9397_out1 XOR Logical_Operator_out9909_out1;

  Logical_Operator_out10422_out1 <= Logical_Operator_out9398_out1 XOR Logical_Operator_out9910_out1;

  Logical_Operator_out10423_out1 <= Logical_Operator_out9399_out1 XOR Logical_Operator_out9911_out1;

  Logical_Operator_out10424_out1 <= Logical_Operator_out9400_out1 XOR Logical_Operator_out9912_out1;

  Logical_Operator_out10425_out1 <= Logical_Operator_out9401_out1 XOR Logical_Operator_out9913_out1;

  Logical_Operator_out10426_out1 <= Logical_Operator_out9402_out1 XOR Logical_Operator_out9914_out1;

  Logical_Operator_out10427_out1 <= Logical_Operator_out9403_out1 XOR Logical_Operator_out9915_out1;

  Logical_Operator_out10428_out1 <= Logical_Operator_out9404_out1 XOR Logical_Operator_out9916_out1;

  Logical_Operator_out10429_out1 <= Logical_Operator_out9405_out1 XOR Logical_Operator_out9917_out1;

  Logical_Operator_out10430_out1 <= Logical_Operator_out9406_out1 XOR Logical_Operator_out9918_out1;

  Logical_Operator_out10431_out1 <= Logical_Operator_out9407_out1 XOR Logical_Operator_out9919_out1;

  Logical_Operator_out10432_out1 <= Logical_Operator_out9408_out1 XOR Logical_Operator_out9920_out1;

  Logical_Operator_out10433_out1 <= Logical_Operator_out9409_out1 XOR Logical_Operator_out9921_out1;

  Logical_Operator_out10434_out1 <= Logical_Operator_out9410_out1 XOR Logical_Operator_out9922_out1;

  Logical_Operator_out10435_out1 <= Logical_Operator_out9411_out1 XOR Logical_Operator_out9923_out1;

  Logical_Operator_out10436_out1 <= Logical_Operator_out9412_out1 XOR Logical_Operator_out9924_out1;

  Logical_Operator_out10437_out1 <= Logical_Operator_out9413_out1 XOR Logical_Operator_out9925_out1;

  Logical_Operator_out10438_out1 <= Logical_Operator_out9414_out1 XOR Logical_Operator_out9926_out1;

  Logical_Operator_out10439_out1 <= Logical_Operator_out9415_out1 XOR Logical_Operator_out9927_out1;

  Logical_Operator_out10440_out1 <= Logical_Operator_out9416_out1 XOR Logical_Operator_out9928_out1;

  Logical_Operator_out10441_out1 <= Logical_Operator_out9417_out1 XOR Logical_Operator_out9929_out1;

  Logical_Operator_out10442_out1 <= Logical_Operator_out9418_out1 XOR Logical_Operator_out9930_out1;

  Logical_Operator_out10443_out1 <= Logical_Operator_out9419_out1 XOR Logical_Operator_out9931_out1;

  Logical_Operator_out10444_out1 <= Logical_Operator_out9420_out1 XOR Logical_Operator_out9932_out1;

  Logical_Operator_out10445_out1 <= Logical_Operator_out9421_out1 XOR Logical_Operator_out9933_out1;

  Logical_Operator_out10446_out1 <= Logical_Operator_out9422_out1 XOR Logical_Operator_out9934_out1;

  Logical_Operator_out10447_out1 <= Logical_Operator_out9423_out1 XOR Logical_Operator_out9935_out1;

  Logical_Operator_out10448_out1 <= Logical_Operator_out9424_out1 XOR Logical_Operator_out9936_out1;

  Logical_Operator_out10449_out1 <= Logical_Operator_out9425_out1 XOR Logical_Operator_out9937_out1;

  Logical_Operator_out10450_out1 <= Logical_Operator_out9426_out1 XOR Logical_Operator_out9938_out1;

  Logical_Operator_out10451_out1 <= Logical_Operator_out9427_out1 XOR Logical_Operator_out9939_out1;

  Logical_Operator_out10452_out1 <= Logical_Operator_out9428_out1 XOR Logical_Operator_out9940_out1;

  Logical_Operator_out10453_out1 <= Logical_Operator_out9429_out1 XOR Logical_Operator_out9941_out1;

  Logical_Operator_out10454_out1 <= Logical_Operator_out9430_out1 XOR Logical_Operator_out9942_out1;

  Logical_Operator_out10455_out1 <= Logical_Operator_out9431_out1 XOR Logical_Operator_out9943_out1;

  Logical_Operator_out10456_out1 <= Logical_Operator_out9432_out1 XOR Logical_Operator_out9944_out1;

  Logical_Operator_out10457_out1 <= Logical_Operator_out9433_out1 XOR Logical_Operator_out9945_out1;

  Logical_Operator_out10458_out1 <= Logical_Operator_out9434_out1 XOR Logical_Operator_out9946_out1;

  Logical_Operator_out10459_out1 <= Logical_Operator_out9435_out1 XOR Logical_Operator_out9947_out1;

  Logical_Operator_out10460_out1 <= Logical_Operator_out9436_out1 XOR Logical_Operator_out9948_out1;

  Logical_Operator_out10461_out1 <= Logical_Operator_out9437_out1 XOR Logical_Operator_out9949_out1;

  Logical_Operator_out10462_out1 <= Logical_Operator_out9438_out1 XOR Logical_Operator_out9950_out1;

  Logical_Operator_out10463_out1 <= Logical_Operator_out9439_out1 XOR Logical_Operator_out9951_out1;

  Logical_Operator_out10464_out1 <= Logical_Operator_out9440_out1 XOR Logical_Operator_out9952_out1;

  Logical_Operator_out10465_out1 <= Logical_Operator_out9441_out1 XOR Logical_Operator_out9953_out1;

  Logical_Operator_out10466_out1 <= Logical_Operator_out9442_out1 XOR Logical_Operator_out9954_out1;

  Logical_Operator_out10467_out1 <= Logical_Operator_out9443_out1 XOR Logical_Operator_out9955_out1;

  Logical_Operator_out10468_out1 <= Logical_Operator_out9444_out1 XOR Logical_Operator_out9956_out1;

  Logical_Operator_out10469_out1 <= Logical_Operator_out9445_out1 XOR Logical_Operator_out9957_out1;

  Logical_Operator_out10470_out1 <= Logical_Operator_out9446_out1 XOR Logical_Operator_out9958_out1;

  Logical_Operator_out10471_out1 <= Logical_Operator_out9447_out1 XOR Logical_Operator_out9959_out1;

  Logical_Operator_out10472_out1 <= Logical_Operator_out9448_out1 XOR Logical_Operator_out9960_out1;

  Logical_Operator_out10473_out1 <= Logical_Operator_out9449_out1 XOR Logical_Operator_out9961_out1;

  Logical_Operator_out10474_out1 <= Logical_Operator_out9450_out1 XOR Logical_Operator_out9962_out1;

  Logical_Operator_out10475_out1 <= Logical_Operator_out9451_out1 XOR Logical_Operator_out9963_out1;

  Logical_Operator_out10476_out1 <= Logical_Operator_out9452_out1 XOR Logical_Operator_out9964_out1;

  Logical_Operator_out10477_out1 <= Logical_Operator_out9453_out1 XOR Logical_Operator_out9965_out1;

  Logical_Operator_out10478_out1 <= Logical_Operator_out9454_out1 XOR Logical_Operator_out9966_out1;

  Logical_Operator_out10479_out1 <= Logical_Operator_out9455_out1 XOR Logical_Operator_out9967_out1;

  Logical_Operator_out10480_out1 <= Logical_Operator_out9456_out1 XOR Logical_Operator_out9968_out1;

  Logical_Operator_out10481_out1 <= Logical_Operator_out9457_out1 XOR Logical_Operator_out9969_out1;

  Logical_Operator_out10482_out1 <= Logical_Operator_out9458_out1 XOR Logical_Operator_out9970_out1;

  Logical_Operator_out10483_out1 <= Logical_Operator_out9459_out1 XOR Logical_Operator_out9971_out1;

  Logical_Operator_out10484_out1 <= Logical_Operator_out9460_out1 XOR Logical_Operator_out9972_out1;

  Logical_Operator_out10485_out1 <= Logical_Operator_out9461_out1 XOR Logical_Operator_out9973_out1;

  Logical_Operator_out10486_out1 <= Logical_Operator_out9462_out1 XOR Logical_Operator_out9974_out1;

  Logical_Operator_out10487_out1 <= Logical_Operator_out9463_out1 XOR Logical_Operator_out9975_out1;

  Logical_Operator_out10488_out1 <= Logical_Operator_out9464_out1 XOR Logical_Operator_out9976_out1;

  Logical_Operator_out10489_out1 <= Logical_Operator_out9465_out1 XOR Logical_Operator_out9977_out1;

  Logical_Operator_out10490_out1 <= Logical_Operator_out9466_out1 XOR Logical_Operator_out9978_out1;

  Logical_Operator_out10491_out1 <= Logical_Operator_out9467_out1 XOR Logical_Operator_out9979_out1;

  Logical_Operator_out10492_out1 <= Logical_Operator_out9468_out1 XOR Logical_Operator_out9980_out1;

  Logical_Operator_out10493_out1 <= Logical_Operator_out9469_out1 XOR Logical_Operator_out9981_out1;

  Logical_Operator_out10494_out1 <= Logical_Operator_out9470_out1 XOR Logical_Operator_out9982_out1;

  Logical_Operator_out10495_out1 <= Logical_Operator_out9471_out1 XOR Logical_Operator_out9983_out1;

  Logical_Operator_out10496_out1 <= Logical_Operator_out9472_out1 XOR Logical_Operator_out9984_out1;

  Logical_Operator_out10497_out1 <= Logical_Operator_out9473_out1 XOR Logical_Operator_out9985_out1;

  Logical_Operator_out10498_out1 <= Logical_Operator_out9474_out1 XOR Logical_Operator_out9986_out1;

  Logical_Operator_out10499_out1 <= Logical_Operator_out9475_out1 XOR Logical_Operator_out9987_out1;

  Logical_Operator_out10500_out1 <= Logical_Operator_out9476_out1 XOR Logical_Operator_out9988_out1;

  Logical_Operator_out10501_out1 <= Logical_Operator_out9477_out1 XOR Logical_Operator_out9989_out1;

  Logical_Operator_out10502_out1 <= Logical_Operator_out9478_out1 XOR Logical_Operator_out9990_out1;

  Logical_Operator_out10503_out1 <= Logical_Operator_out9479_out1 XOR Logical_Operator_out9991_out1;

  Logical_Operator_out10504_out1 <= Logical_Operator_out9480_out1 XOR Logical_Operator_out9992_out1;

  Logical_Operator_out10505_out1 <= Logical_Operator_out9481_out1 XOR Logical_Operator_out9993_out1;

  Logical_Operator_out10506_out1 <= Logical_Operator_out9482_out1 XOR Logical_Operator_out9994_out1;

  Logical_Operator_out10507_out1 <= Logical_Operator_out9483_out1 XOR Logical_Operator_out9995_out1;

  Logical_Operator_out10508_out1 <= Logical_Operator_out9484_out1 XOR Logical_Operator_out9996_out1;

  Logical_Operator_out10509_out1 <= Logical_Operator_out9485_out1 XOR Logical_Operator_out9997_out1;

  Logical_Operator_out10510_out1 <= Logical_Operator_out9486_out1 XOR Logical_Operator_out9998_out1;

  Logical_Operator_out10511_out1 <= Logical_Operator_out9487_out1 XOR Logical_Operator_out9999_out1;

  Logical_Operator_out10512_out1 <= Logical_Operator_out9488_out1 XOR Logical_Operator_out10000_out1;

  Logical_Operator_out10513_out1 <= Logical_Operator_out9489_out1 XOR Logical_Operator_out10001_out1;

  Logical_Operator_out10514_out1 <= Logical_Operator_out9490_out1 XOR Logical_Operator_out10002_out1;

  Logical_Operator_out10515_out1 <= Logical_Operator_out9491_out1 XOR Logical_Operator_out10003_out1;

  Logical_Operator_out10516_out1 <= Logical_Operator_out9492_out1 XOR Logical_Operator_out10004_out1;

  Logical_Operator_out10517_out1 <= Logical_Operator_out9493_out1 XOR Logical_Operator_out10005_out1;

  Logical_Operator_out10518_out1 <= Logical_Operator_out9494_out1 XOR Logical_Operator_out10006_out1;

  Logical_Operator_out10519_out1 <= Logical_Operator_out9495_out1 XOR Logical_Operator_out10007_out1;

  Logical_Operator_out10520_out1 <= Logical_Operator_out9496_out1 XOR Logical_Operator_out10008_out1;

  Logical_Operator_out10521_out1 <= Logical_Operator_out9497_out1 XOR Logical_Operator_out10009_out1;

  Logical_Operator_out10522_out1 <= Logical_Operator_out9498_out1 XOR Logical_Operator_out10010_out1;

  Logical_Operator_out10523_out1 <= Logical_Operator_out9499_out1 XOR Logical_Operator_out10011_out1;

  Logical_Operator_out10524_out1 <= Logical_Operator_out9500_out1 XOR Logical_Operator_out10012_out1;

  Logical_Operator_out10525_out1 <= Logical_Operator_out9501_out1 XOR Logical_Operator_out10013_out1;

  Logical_Operator_out10526_out1 <= Logical_Operator_out9502_out1 XOR Logical_Operator_out10014_out1;

  Logical_Operator_out10527_out1 <= Logical_Operator_out9503_out1 XOR Logical_Operator_out10015_out1;

  Logical_Operator_out10528_out1 <= Logical_Operator_out9504_out1 XOR Logical_Operator_out10016_out1;

  Logical_Operator_out10529_out1 <= Logical_Operator_out9505_out1 XOR Logical_Operator_out10017_out1;

  Logical_Operator_out10530_out1 <= Logical_Operator_out9506_out1 XOR Logical_Operator_out10018_out1;

  Logical_Operator_out10531_out1 <= Logical_Operator_out9507_out1 XOR Logical_Operator_out10019_out1;

  Logical_Operator_out10532_out1 <= Logical_Operator_out9508_out1 XOR Logical_Operator_out10020_out1;

  Logical_Operator_out10533_out1 <= Logical_Operator_out9509_out1 XOR Logical_Operator_out10021_out1;

  Logical_Operator_out10534_out1 <= Logical_Operator_out9510_out1 XOR Logical_Operator_out10022_out1;

  Logical_Operator_out10535_out1 <= Logical_Operator_out9511_out1 XOR Logical_Operator_out10023_out1;

  Logical_Operator_out10536_out1 <= Logical_Operator_out9512_out1 XOR Logical_Operator_out10024_out1;

  Logical_Operator_out10537_out1 <= Logical_Operator_out9513_out1 XOR Logical_Operator_out10025_out1;

  Logical_Operator_out10538_out1 <= Logical_Operator_out9514_out1 XOR Logical_Operator_out10026_out1;

  Logical_Operator_out10539_out1 <= Logical_Operator_out9515_out1 XOR Logical_Operator_out10027_out1;

  Logical_Operator_out10540_out1 <= Logical_Operator_out9516_out1 XOR Logical_Operator_out10028_out1;

  Logical_Operator_out10541_out1 <= Logical_Operator_out9517_out1 XOR Logical_Operator_out10029_out1;

  Logical_Operator_out10542_out1 <= Logical_Operator_out9518_out1 XOR Logical_Operator_out10030_out1;

  Logical_Operator_out10543_out1 <= Logical_Operator_out9519_out1 XOR Logical_Operator_out10031_out1;

  Logical_Operator_out10544_out1 <= Logical_Operator_out9520_out1 XOR Logical_Operator_out10032_out1;

  Logical_Operator_out10545_out1 <= Logical_Operator_out9521_out1 XOR Logical_Operator_out10033_out1;

  Logical_Operator_out10546_out1 <= Logical_Operator_out9522_out1 XOR Logical_Operator_out10034_out1;

  Logical_Operator_out10547_out1 <= Logical_Operator_out9523_out1 XOR Logical_Operator_out10035_out1;

  Logical_Operator_out10548_out1 <= Logical_Operator_out9524_out1 XOR Logical_Operator_out10036_out1;

  Logical_Operator_out10549_out1 <= Logical_Operator_out9525_out1 XOR Logical_Operator_out10037_out1;

  Logical_Operator_out10550_out1 <= Logical_Operator_out9526_out1 XOR Logical_Operator_out10038_out1;

  Logical_Operator_out10551_out1 <= Logical_Operator_out9527_out1 XOR Logical_Operator_out10039_out1;

  Logical_Operator_out10552_out1 <= Logical_Operator_out9528_out1 XOR Logical_Operator_out10040_out1;

  Logical_Operator_out10553_out1 <= Logical_Operator_out9529_out1 XOR Logical_Operator_out10041_out1;

  Logical_Operator_out10554_out1 <= Logical_Operator_out9530_out1 XOR Logical_Operator_out10042_out1;

  Logical_Operator_out10555_out1 <= Logical_Operator_out9531_out1 XOR Logical_Operator_out10043_out1;

  Logical_Operator_out10556_out1 <= Logical_Operator_out9532_out1 XOR Logical_Operator_out10044_out1;

  Logical_Operator_out10557_out1 <= Logical_Operator_out9533_out1 XOR Logical_Operator_out10045_out1;

  Logical_Operator_out10558_out1 <= Logical_Operator_out9534_out1 XOR Logical_Operator_out10046_out1;

  Logical_Operator_out10559_out1 <= Logical_Operator_out9535_out1 XOR Logical_Operator_out10047_out1;

  Logical_Operator_out10560_out1 <= Logical_Operator_out9536_out1 XOR Logical_Operator_out10048_out1;

  Logical_Operator_out10561_out1 <= Logical_Operator_out9537_out1 XOR Logical_Operator_out10049_out1;

  Logical_Operator_out10562_out1 <= Logical_Operator_out9538_out1 XOR Logical_Operator_out10050_out1;

  Logical_Operator_out10563_out1 <= Logical_Operator_out9539_out1 XOR Logical_Operator_out10051_out1;

  Logical_Operator_out10564_out1 <= Logical_Operator_out9540_out1 XOR Logical_Operator_out10052_out1;

  Logical_Operator_out10565_out1 <= Logical_Operator_out9541_out1 XOR Logical_Operator_out10053_out1;

  Logical_Operator_out10566_out1 <= Logical_Operator_out9542_out1 XOR Logical_Operator_out10054_out1;

  Logical_Operator_out10567_out1 <= Logical_Operator_out9543_out1 XOR Logical_Operator_out10055_out1;

  Logical_Operator_out10568_out1 <= Logical_Operator_out9544_out1 XOR Logical_Operator_out10056_out1;

  Logical_Operator_out10569_out1 <= Logical_Operator_out9545_out1 XOR Logical_Operator_out10057_out1;

  Logical_Operator_out10570_out1 <= Logical_Operator_out9546_out1 XOR Logical_Operator_out10058_out1;

  Logical_Operator_out10571_out1 <= Logical_Operator_out9547_out1 XOR Logical_Operator_out10059_out1;

  Logical_Operator_out10572_out1 <= Logical_Operator_out9548_out1 XOR Logical_Operator_out10060_out1;

  Logical_Operator_out10573_out1 <= Logical_Operator_out9549_out1 XOR Logical_Operator_out10061_out1;

  Logical_Operator_out10574_out1 <= Logical_Operator_out9550_out1 XOR Logical_Operator_out10062_out1;

  Logical_Operator_out10575_out1 <= Logical_Operator_out9551_out1 XOR Logical_Operator_out10063_out1;

  Logical_Operator_out10576_out1 <= Logical_Operator_out9552_out1 XOR Logical_Operator_out10064_out1;

  Logical_Operator_out10577_out1 <= Logical_Operator_out9553_out1 XOR Logical_Operator_out10065_out1;

  Logical_Operator_out10578_out1 <= Logical_Operator_out9554_out1 XOR Logical_Operator_out10066_out1;

  Logical_Operator_out10579_out1 <= Logical_Operator_out9555_out1 XOR Logical_Operator_out10067_out1;

  Logical_Operator_out10580_out1 <= Logical_Operator_out9556_out1 XOR Logical_Operator_out10068_out1;

  Logical_Operator_out10581_out1 <= Logical_Operator_out9557_out1 XOR Logical_Operator_out10069_out1;

  Logical_Operator_out10582_out1 <= Logical_Operator_out9558_out1 XOR Logical_Operator_out10070_out1;

  Logical_Operator_out10583_out1 <= Logical_Operator_out9559_out1 XOR Logical_Operator_out10071_out1;

  Logical_Operator_out10584_out1 <= Logical_Operator_out9560_out1 XOR Logical_Operator_out10072_out1;

  Logical_Operator_out10585_out1 <= Logical_Operator_out9561_out1 XOR Logical_Operator_out10073_out1;

  Logical_Operator_out10586_out1 <= Logical_Operator_out9562_out1 XOR Logical_Operator_out10074_out1;

  Logical_Operator_out10587_out1 <= Logical_Operator_out9563_out1 XOR Logical_Operator_out10075_out1;

  Logical_Operator_out10588_out1 <= Logical_Operator_out9564_out1 XOR Logical_Operator_out10076_out1;

  Logical_Operator_out10589_out1 <= Logical_Operator_out9565_out1 XOR Logical_Operator_out10077_out1;

  Logical_Operator_out10590_out1 <= Logical_Operator_out9566_out1 XOR Logical_Operator_out10078_out1;

  Logical_Operator_out10591_out1 <= Logical_Operator_out9567_out1 XOR Logical_Operator_out10079_out1;

  Logical_Operator_out10592_out1 <= Logical_Operator_out9568_out1 XOR Logical_Operator_out10080_out1;

  Logical_Operator_out10593_out1 <= Logical_Operator_out9569_out1 XOR Logical_Operator_out10081_out1;

  Logical_Operator_out10594_out1 <= Logical_Operator_out9570_out1 XOR Logical_Operator_out10082_out1;

  Logical_Operator_out10595_out1 <= Logical_Operator_out9571_out1 XOR Logical_Operator_out10083_out1;

  Logical_Operator_out10596_out1 <= Logical_Operator_out9572_out1 XOR Logical_Operator_out10084_out1;

  Logical_Operator_out10597_out1 <= Logical_Operator_out9573_out1 XOR Logical_Operator_out10085_out1;

  Logical_Operator_out10598_out1 <= Logical_Operator_out9574_out1 XOR Logical_Operator_out10086_out1;

  Logical_Operator_out10599_out1 <= Logical_Operator_out9575_out1 XOR Logical_Operator_out10087_out1;

  Logical_Operator_out10600_out1 <= Logical_Operator_out9576_out1 XOR Logical_Operator_out10088_out1;

  Logical_Operator_out10601_out1 <= Logical_Operator_out9577_out1 XOR Logical_Operator_out10089_out1;

  Logical_Operator_out10602_out1 <= Logical_Operator_out9578_out1 XOR Logical_Operator_out10090_out1;

  Logical_Operator_out10603_out1 <= Logical_Operator_out9579_out1 XOR Logical_Operator_out10091_out1;

  Logical_Operator_out10604_out1 <= Logical_Operator_out9580_out1 XOR Logical_Operator_out10092_out1;

  Logical_Operator_out10605_out1 <= Logical_Operator_out9581_out1 XOR Logical_Operator_out10093_out1;

  Logical_Operator_out10606_out1 <= Logical_Operator_out9582_out1 XOR Logical_Operator_out10094_out1;

  Logical_Operator_out10607_out1 <= Logical_Operator_out9583_out1 XOR Logical_Operator_out10095_out1;

  Logical_Operator_out10608_out1 <= Logical_Operator_out9584_out1 XOR Logical_Operator_out10096_out1;

  Logical_Operator_out10609_out1 <= Logical_Operator_out9585_out1 XOR Logical_Operator_out10097_out1;

  Logical_Operator_out10610_out1 <= Logical_Operator_out9586_out1 XOR Logical_Operator_out10098_out1;

  Logical_Operator_out10611_out1 <= Logical_Operator_out9587_out1 XOR Logical_Operator_out10099_out1;

  Logical_Operator_out10612_out1 <= Logical_Operator_out9588_out1 XOR Logical_Operator_out10100_out1;

  Logical_Operator_out10613_out1 <= Logical_Operator_out9589_out1 XOR Logical_Operator_out10101_out1;

  Logical_Operator_out10614_out1 <= Logical_Operator_out9590_out1 XOR Logical_Operator_out10102_out1;

  Logical_Operator_out10615_out1 <= Logical_Operator_out9591_out1 XOR Logical_Operator_out10103_out1;

  Logical_Operator_out10616_out1 <= Logical_Operator_out9592_out1 XOR Logical_Operator_out10104_out1;

  Logical_Operator_out10617_out1 <= Logical_Operator_out9593_out1 XOR Logical_Operator_out10105_out1;

  Logical_Operator_out10618_out1 <= Logical_Operator_out9594_out1 XOR Logical_Operator_out10106_out1;

  Logical_Operator_out10619_out1 <= Logical_Operator_out9595_out1 XOR Logical_Operator_out10107_out1;

  Logical_Operator_out10620_out1 <= Logical_Operator_out9596_out1 XOR Logical_Operator_out10108_out1;

  Logical_Operator_out10621_out1 <= Logical_Operator_out9597_out1 XOR Logical_Operator_out10109_out1;

  Logical_Operator_out10622_out1 <= Logical_Operator_out9598_out1 XOR Logical_Operator_out10110_out1;

  Logical_Operator_out10623_out1 <= Logical_Operator_out9599_out1 XOR Logical_Operator_out10111_out1;

  Logical_Operator_out10624_out1 <= Logical_Operator_out9600_out1 XOR Logical_Operator_out10112_out1;

  Logical_Operator_out10625_out1 <= Logical_Operator_out9601_out1 XOR Logical_Operator_out10113_out1;

  Logical_Operator_out10626_out1 <= Logical_Operator_out9602_out1 XOR Logical_Operator_out10114_out1;

  Logical_Operator_out10627_out1 <= Logical_Operator_out9603_out1 XOR Logical_Operator_out10115_out1;

  Logical_Operator_out10628_out1 <= Logical_Operator_out9604_out1 XOR Logical_Operator_out10116_out1;

  Logical_Operator_out10629_out1 <= Logical_Operator_out9605_out1 XOR Logical_Operator_out10117_out1;

  Logical_Operator_out10630_out1 <= Logical_Operator_out9606_out1 XOR Logical_Operator_out10118_out1;

  Logical_Operator_out10631_out1 <= Logical_Operator_out9607_out1 XOR Logical_Operator_out10119_out1;

  Logical_Operator_out10632_out1 <= Logical_Operator_out9608_out1 XOR Logical_Operator_out10120_out1;

  Logical_Operator_out10633_out1 <= Logical_Operator_out9609_out1 XOR Logical_Operator_out10121_out1;

  Logical_Operator_out10634_out1 <= Logical_Operator_out9610_out1 XOR Logical_Operator_out10122_out1;

  Logical_Operator_out10635_out1 <= Logical_Operator_out9611_out1 XOR Logical_Operator_out10123_out1;

  Logical_Operator_out10636_out1 <= Logical_Operator_out9612_out1 XOR Logical_Operator_out10124_out1;

  Logical_Operator_out10637_out1 <= Logical_Operator_out9613_out1 XOR Logical_Operator_out10125_out1;

  Logical_Operator_out10638_out1 <= Logical_Operator_out9614_out1 XOR Logical_Operator_out10126_out1;

  Logical_Operator_out10639_out1 <= Logical_Operator_out9615_out1 XOR Logical_Operator_out10127_out1;

  Logical_Operator_out10640_out1 <= Logical_Operator_out9616_out1 XOR Logical_Operator_out10128_out1;

  Logical_Operator_out10641_out1 <= Logical_Operator_out9617_out1 XOR Logical_Operator_out10129_out1;

  Logical_Operator_out10642_out1 <= Logical_Operator_out9618_out1 XOR Logical_Operator_out10130_out1;

  Logical_Operator_out10643_out1 <= Logical_Operator_out9619_out1 XOR Logical_Operator_out10131_out1;

  Logical_Operator_out10644_out1 <= Logical_Operator_out9620_out1 XOR Logical_Operator_out10132_out1;

  Logical_Operator_out10645_out1 <= Logical_Operator_out9621_out1 XOR Logical_Operator_out10133_out1;

  Logical_Operator_out10646_out1 <= Logical_Operator_out9622_out1 XOR Logical_Operator_out10134_out1;

  Logical_Operator_out10647_out1 <= Logical_Operator_out9623_out1 XOR Logical_Operator_out10135_out1;

  Logical_Operator_out10648_out1 <= Logical_Operator_out9624_out1 XOR Logical_Operator_out10136_out1;

  Logical_Operator_out10649_out1 <= Logical_Operator_out9625_out1 XOR Logical_Operator_out10137_out1;

  Logical_Operator_out10650_out1 <= Logical_Operator_out9626_out1 XOR Logical_Operator_out10138_out1;

  Logical_Operator_out10651_out1 <= Logical_Operator_out9627_out1 XOR Logical_Operator_out10139_out1;

  Logical_Operator_out10652_out1 <= Logical_Operator_out9628_out1 XOR Logical_Operator_out10140_out1;

  Logical_Operator_out10653_out1 <= Logical_Operator_out9629_out1 XOR Logical_Operator_out10141_out1;

  Logical_Operator_out10654_out1 <= Logical_Operator_out9630_out1 XOR Logical_Operator_out10142_out1;

  Logical_Operator_out10655_out1 <= Logical_Operator_out9631_out1 XOR Logical_Operator_out10143_out1;

  Logical_Operator_out10656_out1 <= Logical_Operator_out9632_out1 XOR Logical_Operator_out10144_out1;

  Logical_Operator_out10657_out1 <= Logical_Operator_out9633_out1 XOR Logical_Operator_out10145_out1;

  Logical_Operator_out10658_out1 <= Logical_Operator_out9634_out1 XOR Logical_Operator_out10146_out1;

  Logical_Operator_out10659_out1 <= Logical_Operator_out9635_out1 XOR Logical_Operator_out10147_out1;

  Logical_Operator_out10660_out1 <= Logical_Operator_out9636_out1 XOR Logical_Operator_out10148_out1;

  Logical_Operator_out10661_out1 <= Logical_Operator_out9637_out1 XOR Logical_Operator_out10149_out1;

  Logical_Operator_out10662_out1 <= Logical_Operator_out9638_out1 XOR Logical_Operator_out10150_out1;

  Logical_Operator_out10663_out1 <= Logical_Operator_out9639_out1 XOR Logical_Operator_out10151_out1;

  Logical_Operator_out10664_out1 <= Logical_Operator_out9640_out1 XOR Logical_Operator_out10152_out1;

  Logical_Operator_out10665_out1 <= Logical_Operator_out9641_out1 XOR Logical_Operator_out10153_out1;

  Logical_Operator_out10666_out1 <= Logical_Operator_out9642_out1 XOR Logical_Operator_out10154_out1;

  Logical_Operator_out10667_out1 <= Logical_Operator_out9643_out1 XOR Logical_Operator_out10155_out1;

  Logical_Operator_out10668_out1 <= Logical_Operator_out9644_out1 XOR Logical_Operator_out10156_out1;

  Logical_Operator_out10669_out1 <= Logical_Operator_out9645_out1 XOR Logical_Operator_out10157_out1;

  Logical_Operator_out10670_out1 <= Logical_Operator_out9646_out1 XOR Logical_Operator_out10158_out1;

  Logical_Operator_out10671_out1 <= Logical_Operator_out9647_out1 XOR Logical_Operator_out10159_out1;

  Logical_Operator_out10672_out1 <= Logical_Operator_out9648_out1 XOR Logical_Operator_out10160_out1;

  Logical_Operator_out10673_out1 <= Logical_Operator_out9649_out1 XOR Logical_Operator_out10161_out1;

  Logical_Operator_out10674_out1 <= Logical_Operator_out9650_out1 XOR Logical_Operator_out10162_out1;

  Logical_Operator_out10675_out1 <= Logical_Operator_out9651_out1 XOR Logical_Operator_out10163_out1;

  Logical_Operator_out10676_out1 <= Logical_Operator_out9652_out1 XOR Logical_Operator_out10164_out1;

  Logical_Operator_out10677_out1 <= Logical_Operator_out9653_out1 XOR Logical_Operator_out10165_out1;

  Logical_Operator_out10678_out1 <= Logical_Operator_out9654_out1 XOR Logical_Operator_out10166_out1;

  Logical_Operator_out10679_out1 <= Logical_Operator_out9655_out1 XOR Logical_Operator_out10167_out1;

  Logical_Operator_out10680_out1 <= Logical_Operator_out9656_out1 XOR Logical_Operator_out10168_out1;

  Logical_Operator_out10681_out1 <= Logical_Operator_out9657_out1 XOR Logical_Operator_out10169_out1;

  Logical_Operator_out10682_out1 <= Logical_Operator_out9658_out1 XOR Logical_Operator_out10170_out1;

  Logical_Operator_out10683_out1 <= Logical_Operator_out9659_out1 XOR Logical_Operator_out10171_out1;

  Logical_Operator_out10684_out1 <= Logical_Operator_out9660_out1 XOR Logical_Operator_out10172_out1;

  Logical_Operator_out10685_out1 <= Logical_Operator_out9661_out1 XOR Logical_Operator_out10173_out1;

  Logical_Operator_out10686_out1 <= Logical_Operator_out9662_out1 XOR Logical_Operator_out10174_out1;

  Logical_Operator_out10687_out1 <= Logical_Operator_out9663_out1 XOR Logical_Operator_out10175_out1;

  Logical_Operator_out10688_out1 <= Logical_Operator_out9664_out1 XOR Logical_Operator_out10176_out1;

  Logical_Operator_out10689_out1 <= Logical_Operator_out9665_out1 XOR Logical_Operator_out10177_out1;

  Logical_Operator_out10690_out1 <= Logical_Operator_out9666_out1 XOR Logical_Operator_out10178_out1;

  Logical_Operator_out10691_out1 <= Logical_Operator_out9667_out1 XOR Logical_Operator_out10179_out1;

  Logical_Operator_out10692_out1 <= Logical_Operator_out9668_out1 XOR Logical_Operator_out10180_out1;

  Logical_Operator_out10693_out1 <= Logical_Operator_out9669_out1 XOR Logical_Operator_out10181_out1;

  Logical_Operator_out10694_out1 <= Logical_Operator_out9670_out1 XOR Logical_Operator_out10182_out1;

  Logical_Operator_out10695_out1 <= Logical_Operator_out9671_out1 XOR Logical_Operator_out10183_out1;

  Logical_Operator_out10696_out1 <= Logical_Operator_out9672_out1 XOR Logical_Operator_out10184_out1;

  Logical_Operator_out10697_out1 <= Logical_Operator_out9673_out1 XOR Logical_Operator_out10185_out1;

  Logical_Operator_out10698_out1 <= Logical_Operator_out9674_out1 XOR Logical_Operator_out10186_out1;

  Logical_Operator_out10699_out1 <= Logical_Operator_out9675_out1 XOR Logical_Operator_out10187_out1;

  Logical_Operator_out10700_out1 <= Logical_Operator_out9676_out1 XOR Logical_Operator_out10188_out1;

  Logical_Operator_out10701_out1 <= Logical_Operator_out9677_out1 XOR Logical_Operator_out10189_out1;

  Logical_Operator_out10702_out1 <= Logical_Operator_out9678_out1 XOR Logical_Operator_out10190_out1;

  Logical_Operator_out10703_out1 <= Logical_Operator_out9679_out1 XOR Logical_Operator_out10191_out1;

  Logical_Operator_out10704_out1 <= Logical_Operator_out9680_out1 XOR Logical_Operator_out10192_out1;

  Logical_Operator_out10705_out1 <= Logical_Operator_out9681_out1 XOR Logical_Operator_out10193_out1;

  Logical_Operator_out10706_out1 <= Logical_Operator_out9682_out1 XOR Logical_Operator_out10194_out1;

  Logical_Operator_out10707_out1 <= Logical_Operator_out9683_out1 XOR Logical_Operator_out10195_out1;

  Logical_Operator_out10708_out1 <= Logical_Operator_out9684_out1 XOR Logical_Operator_out10196_out1;

  Logical_Operator_out10709_out1 <= Logical_Operator_out9685_out1 XOR Logical_Operator_out10197_out1;

  Logical_Operator_out10710_out1 <= Logical_Operator_out9686_out1 XOR Logical_Operator_out10198_out1;

  Logical_Operator_out10711_out1 <= Logical_Operator_out9687_out1 XOR Logical_Operator_out10199_out1;

  Logical_Operator_out10712_out1 <= Logical_Operator_out9688_out1 XOR Logical_Operator_out10200_out1;

  Logical_Operator_out10713_out1 <= Logical_Operator_out9689_out1 XOR Logical_Operator_out10201_out1;

  Logical_Operator_out10714_out1 <= Logical_Operator_out9690_out1 XOR Logical_Operator_out10202_out1;

  Logical_Operator_out10715_out1 <= Logical_Operator_out9691_out1 XOR Logical_Operator_out10203_out1;

  Logical_Operator_out10716_out1 <= Logical_Operator_out9692_out1 XOR Logical_Operator_out10204_out1;

  Logical_Operator_out10717_out1 <= Logical_Operator_out9693_out1 XOR Logical_Operator_out10205_out1;

  Logical_Operator_out10718_out1 <= Logical_Operator_out9694_out1 XOR Logical_Operator_out10206_out1;

  Logical_Operator_out10719_out1 <= Logical_Operator_out9695_out1 XOR Logical_Operator_out10207_out1;

  Logical_Operator_out10720_out1 <= Logical_Operator_out9696_out1 XOR Logical_Operator_out10208_out1;

  Logical_Operator_out10721_out1 <= Logical_Operator_out9697_out1 XOR Logical_Operator_out10209_out1;

  Logical_Operator_out10722_out1 <= Logical_Operator_out9698_out1 XOR Logical_Operator_out10210_out1;

  Logical_Operator_out10723_out1 <= Logical_Operator_out9699_out1 XOR Logical_Operator_out10211_out1;

  Logical_Operator_out10724_out1 <= Logical_Operator_out9700_out1 XOR Logical_Operator_out10212_out1;

  Logical_Operator_out10725_out1 <= Logical_Operator_out9701_out1 XOR Logical_Operator_out10213_out1;

  Logical_Operator_out10726_out1 <= Logical_Operator_out9702_out1 XOR Logical_Operator_out10214_out1;

  Logical_Operator_out10727_out1 <= Logical_Operator_out9703_out1 XOR Logical_Operator_out10215_out1;

  Logical_Operator_out10728_out1 <= Logical_Operator_out9704_out1 XOR Logical_Operator_out10216_out1;

  Logical_Operator_out10729_out1 <= Logical_Operator_out9705_out1 XOR Logical_Operator_out10217_out1;

  Logical_Operator_out10730_out1 <= Logical_Operator_out9706_out1 XOR Logical_Operator_out10218_out1;

  Logical_Operator_out10731_out1 <= Logical_Operator_out9707_out1 XOR Logical_Operator_out10219_out1;

  Logical_Operator_out10732_out1 <= Logical_Operator_out9708_out1 XOR Logical_Operator_out10220_out1;

  Logical_Operator_out10733_out1 <= Logical_Operator_out9709_out1 XOR Logical_Operator_out10221_out1;

  Logical_Operator_out10734_out1 <= Logical_Operator_out9710_out1 XOR Logical_Operator_out10222_out1;

  Logical_Operator_out10735_out1 <= Logical_Operator_out9711_out1 XOR Logical_Operator_out10223_out1;

  Logical_Operator_out10736_out1 <= Logical_Operator_out9712_out1 XOR Logical_Operator_out10224_out1;

  Logical_Operator_out10737_out1 <= Logical_Operator_out9713_out1 XOR Logical_Operator_out10225_out1;

  Logical_Operator_out10738_out1 <= Logical_Operator_out9714_out1 XOR Logical_Operator_out10226_out1;

  Logical_Operator_out10739_out1 <= Logical_Operator_out9715_out1 XOR Logical_Operator_out10227_out1;

  Logical_Operator_out10740_out1 <= Logical_Operator_out9716_out1 XOR Logical_Operator_out10228_out1;

  Logical_Operator_out10741_out1 <= Logical_Operator_out9717_out1 XOR Logical_Operator_out10229_out1;

  Logical_Operator_out10742_out1 <= Logical_Operator_out9718_out1 XOR Logical_Operator_out10230_out1;

  Logical_Operator_out10743_out1 <= Logical_Operator_out9719_out1 XOR Logical_Operator_out10231_out1;

  Logical_Operator_out10744_out1 <= Logical_Operator_out9720_out1 XOR Logical_Operator_out10232_out1;

  Logical_Operator_out10745_out1 <= Logical_Operator_out9721_out1 XOR Logical_Operator_out10233_out1;

  Logical_Operator_out10746_out1 <= Logical_Operator_out9722_out1 XOR Logical_Operator_out10234_out1;

  Logical_Operator_out10747_out1 <= Logical_Operator_out9723_out1 XOR Logical_Operator_out10235_out1;

  Logical_Operator_out10748_out1 <= Logical_Operator_out9724_out1 XOR Logical_Operator_out10236_out1;

  Logical_Operator_out10749_out1 <= Logical_Operator_out9725_out1 XOR Logical_Operator_out10237_out1;

  Logical_Operator_out10750_out1 <= Logical_Operator_out9726_out1 XOR Logical_Operator_out10238_out1;

  Logical_Operator_out10751_out1 <= Logical_Operator_out9727_out1 XOR Logical_Operator_out10239_out1;

  Logical_Operator_out10752_out1 <= Logical_Operator_out9728_out1 XOR Logical_Operator_out10240_out1;

  Logical_Operator_out10753_out1 <= Logical_Operator_out8449_out1 XOR Logical_Operator_out8961_out1;

  Logical_Operator_out10754_out1 <= Logical_Operator_out8450_out1 XOR Logical_Operator_out8962_out1;

  Logical_Operator_out10755_out1 <= Logical_Operator_out8451_out1 XOR Logical_Operator_out8963_out1;

  Logical_Operator_out10756_out1 <= Logical_Operator_out8452_out1 XOR Logical_Operator_out8964_out1;

  Logical_Operator_out10757_out1 <= Logical_Operator_out8453_out1 XOR Logical_Operator_out8965_out1;

  Logical_Operator_out10758_out1 <= Logical_Operator_out8454_out1 XOR Logical_Operator_out8966_out1;

  Logical_Operator_out10759_out1 <= Logical_Operator_out8455_out1 XOR Logical_Operator_out8967_out1;

  Logical_Operator_out10760_out1 <= Logical_Operator_out8456_out1 XOR Logical_Operator_out8968_out1;

  Logical_Operator_out10761_out1 <= Logical_Operator_out8457_out1 XOR Logical_Operator_out8969_out1;

  Logical_Operator_out10762_out1 <= Logical_Operator_out8458_out1 XOR Logical_Operator_out8970_out1;

  Logical_Operator_out10763_out1 <= Logical_Operator_out8459_out1 XOR Logical_Operator_out8971_out1;

  Logical_Operator_out10764_out1 <= Logical_Operator_out8460_out1 XOR Logical_Operator_out8972_out1;

  Logical_Operator_out10765_out1 <= Logical_Operator_out8461_out1 XOR Logical_Operator_out8973_out1;

  Logical_Operator_out10766_out1 <= Logical_Operator_out8462_out1 XOR Logical_Operator_out8974_out1;

  Logical_Operator_out10767_out1 <= Logical_Operator_out8463_out1 XOR Logical_Operator_out8975_out1;

  Logical_Operator_out10768_out1 <= Logical_Operator_out8464_out1 XOR Logical_Operator_out8976_out1;

  Logical_Operator_out10769_out1 <= Logical_Operator_out8465_out1 XOR Logical_Operator_out8977_out1;

  Logical_Operator_out10770_out1 <= Logical_Operator_out8466_out1 XOR Logical_Operator_out8978_out1;

  Logical_Operator_out10771_out1 <= Logical_Operator_out8467_out1 XOR Logical_Operator_out8979_out1;

  Logical_Operator_out10772_out1 <= Logical_Operator_out8468_out1 XOR Logical_Operator_out8980_out1;

  Logical_Operator_out10773_out1 <= Logical_Operator_out8469_out1 XOR Logical_Operator_out8981_out1;

  Logical_Operator_out10774_out1 <= Logical_Operator_out8470_out1 XOR Logical_Operator_out8982_out1;

  Logical_Operator_out10775_out1 <= Logical_Operator_out8471_out1 XOR Logical_Operator_out8983_out1;

  Logical_Operator_out10776_out1 <= Logical_Operator_out8472_out1 XOR Logical_Operator_out8984_out1;

  Logical_Operator_out10777_out1 <= Logical_Operator_out8473_out1 XOR Logical_Operator_out8985_out1;

  Logical_Operator_out10778_out1 <= Logical_Operator_out8474_out1 XOR Logical_Operator_out8986_out1;

  Logical_Operator_out10779_out1 <= Logical_Operator_out8475_out1 XOR Logical_Operator_out8987_out1;

  Logical_Operator_out10780_out1 <= Logical_Operator_out8476_out1 XOR Logical_Operator_out8988_out1;

  Logical_Operator_out10781_out1 <= Logical_Operator_out8477_out1 XOR Logical_Operator_out8989_out1;

  Logical_Operator_out10782_out1 <= Logical_Operator_out8478_out1 XOR Logical_Operator_out8990_out1;

  Logical_Operator_out10783_out1 <= Logical_Operator_out8479_out1 XOR Logical_Operator_out8991_out1;

  Logical_Operator_out10784_out1 <= Logical_Operator_out8480_out1 XOR Logical_Operator_out8992_out1;

  Logical_Operator_out10785_out1 <= Logical_Operator_out8481_out1 XOR Logical_Operator_out8993_out1;

  Logical_Operator_out10786_out1 <= Logical_Operator_out8482_out1 XOR Logical_Operator_out8994_out1;

  Logical_Operator_out10787_out1 <= Logical_Operator_out8483_out1 XOR Logical_Operator_out8995_out1;

  Logical_Operator_out10788_out1 <= Logical_Operator_out8484_out1 XOR Logical_Operator_out8996_out1;

  Logical_Operator_out10789_out1 <= Logical_Operator_out8485_out1 XOR Logical_Operator_out8997_out1;

  Logical_Operator_out10790_out1 <= Logical_Operator_out8486_out1 XOR Logical_Operator_out8998_out1;

  Logical_Operator_out10791_out1 <= Logical_Operator_out8487_out1 XOR Logical_Operator_out8999_out1;

  Logical_Operator_out10792_out1 <= Logical_Operator_out8488_out1 XOR Logical_Operator_out9000_out1;

  Logical_Operator_out10793_out1 <= Logical_Operator_out8489_out1 XOR Logical_Operator_out9001_out1;

  Logical_Operator_out10794_out1 <= Logical_Operator_out8490_out1 XOR Logical_Operator_out9002_out1;

  Logical_Operator_out10795_out1 <= Logical_Operator_out8491_out1 XOR Logical_Operator_out9003_out1;

  Logical_Operator_out10796_out1 <= Logical_Operator_out8492_out1 XOR Logical_Operator_out9004_out1;

  Logical_Operator_out10797_out1 <= Logical_Operator_out8493_out1 XOR Logical_Operator_out9005_out1;

  Logical_Operator_out10798_out1 <= Logical_Operator_out8494_out1 XOR Logical_Operator_out9006_out1;

  Logical_Operator_out10799_out1 <= Logical_Operator_out8495_out1 XOR Logical_Operator_out9007_out1;

  Logical_Operator_out10800_out1 <= Logical_Operator_out8496_out1 XOR Logical_Operator_out9008_out1;

  Logical_Operator_out10801_out1 <= Logical_Operator_out8497_out1 XOR Logical_Operator_out9009_out1;

  Logical_Operator_out10802_out1 <= Logical_Operator_out8498_out1 XOR Logical_Operator_out9010_out1;

  Logical_Operator_out10803_out1 <= Logical_Operator_out8499_out1 XOR Logical_Operator_out9011_out1;

  Logical_Operator_out10804_out1 <= Logical_Operator_out8500_out1 XOR Logical_Operator_out9012_out1;

  Logical_Operator_out10805_out1 <= Logical_Operator_out8501_out1 XOR Logical_Operator_out9013_out1;

  Logical_Operator_out10806_out1 <= Logical_Operator_out8502_out1 XOR Logical_Operator_out9014_out1;

  Logical_Operator_out10807_out1 <= Logical_Operator_out8503_out1 XOR Logical_Operator_out9015_out1;

  Logical_Operator_out10808_out1 <= Logical_Operator_out8504_out1 XOR Logical_Operator_out9016_out1;

  Logical_Operator_out10809_out1 <= Logical_Operator_out8505_out1 XOR Logical_Operator_out9017_out1;

  Logical_Operator_out10810_out1 <= Logical_Operator_out8506_out1 XOR Logical_Operator_out9018_out1;

  Logical_Operator_out10811_out1 <= Logical_Operator_out8507_out1 XOR Logical_Operator_out9019_out1;

  Logical_Operator_out10812_out1 <= Logical_Operator_out8508_out1 XOR Logical_Operator_out9020_out1;

  Logical_Operator_out10813_out1 <= Logical_Operator_out8509_out1 XOR Logical_Operator_out9021_out1;

  Logical_Operator_out10814_out1 <= Logical_Operator_out8510_out1 XOR Logical_Operator_out9022_out1;

  Logical_Operator_out10815_out1 <= Logical_Operator_out8511_out1 XOR Logical_Operator_out9023_out1;

  Logical_Operator_out10816_out1 <= Logical_Operator_out8512_out1 XOR Logical_Operator_out9024_out1;

  Logical_Operator_out10817_out1 <= Logical_Operator_out8513_out1 XOR Logical_Operator_out9025_out1;

  Logical_Operator_out10818_out1 <= Logical_Operator_out8514_out1 XOR Logical_Operator_out9026_out1;

  Logical_Operator_out10819_out1 <= Logical_Operator_out8515_out1 XOR Logical_Operator_out9027_out1;

  Logical_Operator_out10820_out1 <= Logical_Operator_out8516_out1 XOR Logical_Operator_out9028_out1;

  Logical_Operator_out10821_out1 <= Logical_Operator_out8517_out1 XOR Logical_Operator_out9029_out1;

  Logical_Operator_out10822_out1 <= Logical_Operator_out8518_out1 XOR Logical_Operator_out9030_out1;

  Logical_Operator_out10823_out1 <= Logical_Operator_out8519_out1 XOR Logical_Operator_out9031_out1;

  Logical_Operator_out10824_out1 <= Logical_Operator_out8520_out1 XOR Logical_Operator_out9032_out1;

  Logical_Operator_out10825_out1 <= Logical_Operator_out8521_out1 XOR Logical_Operator_out9033_out1;

  Logical_Operator_out10826_out1 <= Logical_Operator_out8522_out1 XOR Logical_Operator_out9034_out1;

  Logical_Operator_out10827_out1 <= Logical_Operator_out8523_out1 XOR Logical_Operator_out9035_out1;

  Logical_Operator_out10828_out1 <= Logical_Operator_out8524_out1 XOR Logical_Operator_out9036_out1;

  Logical_Operator_out10829_out1 <= Logical_Operator_out8525_out1 XOR Logical_Operator_out9037_out1;

  Logical_Operator_out10830_out1 <= Logical_Operator_out8526_out1 XOR Logical_Operator_out9038_out1;

  Logical_Operator_out10831_out1 <= Logical_Operator_out8527_out1 XOR Logical_Operator_out9039_out1;

  Logical_Operator_out10832_out1 <= Logical_Operator_out8528_out1 XOR Logical_Operator_out9040_out1;

  Logical_Operator_out10833_out1 <= Logical_Operator_out8529_out1 XOR Logical_Operator_out9041_out1;

  Logical_Operator_out10834_out1 <= Logical_Operator_out8530_out1 XOR Logical_Operator_out9042_out1;

  Logical_Operator_out10835_out1 <= Logical_Operator_out8531_out1 XOR Logical_Operator_out9043_out1;

  Logical_Operator_out10836_out1 <= Logical_Operator_out8532_out1 XOR Logical_Operator_out9044_out1;

  Logical_Operator_out10837_out1 <= Logical_Operator_out8533_out1 XOR Logical_Operator_out9045_out1;

  Logical_Operator_out10838_out1 <= Logical_Operator_out8534_out1 XOR Logical_Operator_out9046_out1;

  Logical_Operator_out10839_out1 <= Logical_Operator_out8535_out1 XOR Logical_Operator_out9047_out1;

  Logical_Operator_out10840_out1 <= Logical_Operator_out8536_out1 XOR Logical_Operator_out9048_out1;

  Logical_Operator_out10841_out1 <= Logical_Operator_out8537_out1 XOR Logical_Operator_out9049_out1;

  Logical_Operator_out10842_out1 <= Logical_Operator_out8538_out1 XOR Logical_Operator_out9050_out1;

  Logical_Operator_out10843_out1 <= Logical_Operator_out8539_out1 XOR Logical_Operator_out9051_out1;

  Logical_Operator_out10844_out1 <= Logical_Operator_out8540_out1 XOR Logical_Operator_out9052_out1;

  Logical_Operator_out10845_out1 <= Logical_Operator_out8541_out1 XOR Logical_Operator_out9053_out1;

  Logical_Operator_out10846_out1 <= Logical_Operator_out8542_out1 XOR Logical_Operator_out9054_out1;

  Logical_Operator_out10847_out1 <= Logical_Operator_out8543_out1 XOR Logical_Operator_out9055_out1;

  Logical_Operator_out10848_out1 <= Logical_Operator_out8544_out1 XOR Logical_Operator_out9056_out1;

  Logical_Operator_out10849_out1 <= Logical_Operator_out8545_out1 XOR Logical_Operator_out9057_out1;

  Logical_Operator_out10850_out1 <= Logical_Operator_out8546_out1 XOR Logical_Operator_out9058_out1;

  Logical_Operator_out10851_out1 <= Logical_Operator_out8547_out1 XOR Logical_Operator_out9059_out1;

  Logical_Operator_out10852_out1 <= Logical_Operator_out8548_out1 XOR Logical_Operator_out9060_out1;

  Logical_Operator_out10853_out1 <= Logical_Operator_out8549_out1 XOR Logical_Operator_out9061_out1;

  Logical_Operator_out10854_out1 <= Logical_Operator_out8550_out1 XOR Logical_Operator_out9062_out1;

  Logical_Operator_out10855_out1 <= Logical_Operator_out8551_out1 XOR Logical_Operator_out9063_out1;

  Logical_Operator_out10856_out1 <= Logical_Operator_out8552_out1 XOR Logical_Operator_out9064_out1;

  Logical_Operator_out10857_out1 <= Logical_Operator_out8553_out1 XOR Logical_Operator_out9065_out1;

  Logical_Operator_out10858_out1 <= Logical_Operator_out8554_out1 XOR Logical_Operator_out9066_out1;

  Logical_Operator_out10859_out1 <= Logical_Operator_out8555_out1 XOR Logical_Operator_out9067_out1;

  Logical_Operator_out10860_out1 <= Logical_Operator_out8556_out1 XOR Logical_Operator_out9068_out1;

  Logical_Operator_out10861_out1 <= Logical_Operator_out8557_out1 XOR Logical_Operator_out9069_out1;

  Logical_Operator_out10862_out1 <= Logical_Operator_out8558_out1 XOR Logical_Operator_out9070_out1;

  Logical_Operator_out10863_out1 <= Logical_Operator_out8559_out1 XOR Logical_Operator_out9071_out1;

  Logical_Operator_out10864_out1 <= Logical_Operator_out8560_out1 XOR Logical_Operator_out9072_out1;

  Logical_Operator_out10865_out1 <= Logical_Operator_out8561_out1 XOR Logical_Operator_out9073_out1;

  Logical_Operator_out10866_out1 <= Logical_Operator_out8562_out1 XOR Logical_Operator_out9074_out1;

  Logical_Operator_out10867_out1 <= Logical_Operator_out8563_out1 XOR Logical_Operator_out9075_out1;

  Logical_Operator_out10868_out1 <= Logical_Operator_out8564_out1 XOR Logical_Operator_out9076_out1;

  Logical_Operator_out10869_out1 <= Logical_Operator_out8565_out1 XOR Logical_Operator_out9077_out1;

  Logical_Operator_out10870_out1 <= Logical_Operator_out8566_out1 XOR Logical_Operator_out9078_out1;

  Logical_Operator_out10871_out1 <= Logical_Operator_out8567_out1 XOR Logical_Operator_out9079_out1;

  Logical_Operator_out10872_out1 <= Logical_Operator_out8568_out1 XOR Logical_Operator_out9080_out1;

  Logical_Operator_out10873_out1 <= Logical_Operator_out8569_out1 XOR Logical_Operator_out9081_out1;

  Logical_Operator_out10874_out1 <= Logical_Operator_out8570_out1 XOR Logical_Operator_out9082_out1;

  Logical_Operator_out10875_out1 <= Logical_Operator_out8571_out1 XOR Logical_Operator_out9083_out1;

  Logical_Operator_out10876_out1 <= Logical_Operator_out8572_out1 XOR Logical_Operator_out9084_out1;

  Logical_Operator_out10877_out1 <= Logical_Operator_out8573_out1 XOR Logical_Operator_out9085_out1;

  Logical_Operator_out10878_out1 <= Logical_Operator_out8574_out1 XOR Logical_Operator_out9086_out1;

  Logical_Operator_out10879_out1 <= Logical_Operator_out8575_out1 XOR Logical_Operator_out9087_out1;

  Logical_Operator_out10880_out1 <= Logical_Operator_out8576_out1 XOR Logical_Operator_out9088_out1;

  Logical_Operator_out10881_out1 <= Logical_Operator_out8577_out1 XOR Logical_Operator_out9089_out1;

  Logical_Operator_out10882_out1 <= Logical_Operator_out8578_out1 XOR Logical_Operator_out9090_out1;

  Logical_Operator_out10883_out1 <= Logical_Operator_out8579_out1 XOR Logical_Operator_out9091_out1;

  Logical_Operator_out10884_out1 <= Logical_Operator_out8580_out1 XOR Logical_Operator_out9092_out1;

  Logical_Operator_out10885_out1 <= Logical_Operator_out8581_out1 XOR Logical_Operator_out9093_out1;

  Logical_Operator_out10886_out1 <= Logical_Operator_out8582_out1 XOR Logical_Operator_out9094_out1;

  Logical_Operator_out10887_out1 <= Logical_Operator_out8583_out1 XOR Logical_Operator_out9095_out1;

  Logical_Operator_out10888_out1 <= Logical_Operator_out8584_out1 XOR Logical_Operator_out9096_out1;

  Logical_Operator_out10889_out1 <= Logical_Operator_out8585_out1 XOR Logical_Operator_out9097_out1;

  Logical_Operator_out10890_out1 <= Logical_Operator_out8586_out1 XOR Logical_Operator_out9098_out1;

  Logical_Operator_out10891_out1 <= Logical_Operator_out8587_out1 XOR Logical_Operator_out9099_out1;

  Logical_Operator_out10892_out1 <= Logical_Operator_out8588_out1 XOR Logical_Operator_out9100_out1;

  Logical_Operator_out10893_out1 <= Logical_Operator_out8589_out1 XOR Logical_Operator_out9101_out1;

  Logical_Operator_out10894_out1 <= Logical_Operator_out8590_out1 XOR Logical_Operator_out9102_out1;

  Logical_Operator_out10895_out1 <= Logical_Operator_out8591_out1 XOR Logical_Operator_out9103_out1;

  Logical_Operator_out10896_out1 <= Logical_Operator_out8592_out1 XOR Logical_Operator_out9104_out1;

  Logical_Operator_out10897_out1 <= Logical_Operator_out8593_out1 XOR Logical_Operator_out9105_out1;

  Logical_Operator_out10898_out1 <= Logical_Operator_out8594_out1 XOR Logical_Operator_out9106_out1;

  Logical_Operator_out10899_out1 <= Logical_Operator_out8595_out1 XOR Logical_Operator_out9107_out1;

  Logical_Operator_out10900_out1 <= Logical_Operator_out8596_out1 XOR Logical_Operator_out9108_out1;

  Logical_Operator_out10901_out1 <= Logical_Operator_out8597_out1 XOR Logical_Operator_out9109_out1;

  Logical_Operator_out10902_out1 <= Logical_Operator_out8598_out1 XOR Logical_Operator_out9110_out1;

  Logical_Operator_out10903_out1 <= Logical_Operator_out8599_out1 XOR Logical_Operator_out9111_out1;

  Logical_Operator_out10904_out1 <= Logical_Operator_out8600_out1 XOR Logical_Operator_out9112_out1;

  Logical_Operator_out10905_out1 <= Logical_Operator_out8601_out1 XOR Logical_Operator_out9113_out1;

  Logical_Operator_out10906_out1 <= Logical_Operator_out8602_out1 XOR Logical_Operator_out9114_out1;

  Logical_Operator_out10907_out1 <= Logical_Operator_out8603_out1 XOR Logical_Operator_out9115_out1;

  Logical_Operator_out10908_out1 <= Logical_Operator_out8604_out1 XOR Logical_Operator_out9116_out1;

  Logical_Operator_out10909_out1 <= Logical_Operator_out8605_out1 XOR Logical_Operator_out9117_out1;

  Logical_Operator_out10910_out1 <= Logical_Operator_out8606_out1 XOR Logical_Operator_out9118_out1;

  Logical_Operator_out10911_out1 <= Logical_Operator_out8607_out1 XOR Logical_Operator_out9119_out1;

  Logical_Operator_out10912_out1 <= Logical_Operator_out8608_out1 XOR Logical_Operator_out9120_out1;

  Logical_Operator_out10913_out1 <= Logical_Operator_out8609_out1 XOR Logical_Operator_out9121_out1;

  Logical_Operator_out10914_out1 <= Logical_Operator_out8610_out1 XOR Logical_Operator_out9122_out1;

  Logical_Operator_out10915_out1 <= Logical_Operator_out8611_out1 XOR Logical_Operator_out9123_out1;

  Logical_Operator_out10916_out1 <= Logical_Operator_out8612_out1 XOR Logical_Operator_out9124_out1;

  Logical_Operator_out10917_out1 <= Logical_Operator_out8613_out1 XOR Logical_Operator_out9125_out1;

  Logical_Operator_out10918_out1 <= Logical_Operator_out8614_out1 XOR Logical_Operator_out9126_out1;

  Logical_Operator_out10919_out1 <= Logical_Operator_out8615_out1 XOR Logical_Operator_out9127_out1;

  Logical_Operator_out10920_out1 <= Logical_Operator_out8616_out1 XOR Logical_Operator_out9128_out1;

  Logical_Operator_out10921_out1 <= Logical_Operator_out8617_out1 XOR Logical_Operator_out9129_out1;

  Logical_Operator_out10922_out1 <= Logical_Operator_out8618_out1 XOR Logical_Operator_out9130_out1;

  Logical_Operator_out10923_out1 <= Logical_Operator_out8619_out1 XOR Logical_Operator_out9131_out1;

  Logical_Operator_out10924_out1 <= Logical_Operator_out8620_out1 XOR Logical_Operator_out9132_out1;

  Logical_Operator_out10925_out1 <= Logical_Operator_out8621_out1 XOR Logical_Operator_out9133_out1;

  Logical_Operator_out10926_out1 <= Logical_Operator_out8622_out1 XOR Logical_Operator_out9134_out1;

  Logical_Operator_out10927_out1 <= Logical_Operator_out8623_out1 XOR Logical_Operator_out9135_out1;

  Logical_Operator_out10928_out1 <= Logical_Operator_out8624_out1 XOR Logical_Operator_out9136_out1;

  Logical_Operator_out10929_out1 <= Logical_Operator_out8625_out1 XOR Logical_Operator_out9137_out1;

  Logical_Operator_out10930_out1 <= Logical_Operator_out8626_out1 XOR Logical_Operator_out9138_out1;

  Logical_Operator_out10931_out1 <= Logical_Operator_out8627_out1 XOR Logical_Operator_out9139_out1;

  Logical_Operator_out10932_out1 <= Logical_Operator_out8628_out1 XOR Logical_Operator_out9140_out1;

  Logical_Operator_out10933_out1 <= Logical_Operator_out8629_out1 XOR Logical_Operator_out9141_out1;

  Logical_Operator_out10934_out1 <= Logical_Operator_out8630_out1 XOR Logical_Operator_out9142_out1;

  Logical_Operator_out10935_out1 <= Logical_Operator_out8631_out1 XOR Logical_Operator_out9143_out1;

  Logical_Operator_out10936_out1 <= Logical_Operator_out8632_out1 XOR Logical_Operator_out9144_out1;

  Logical_Operator_out10937_out1 <= Logical_Operator_out8633_out1 XOR Logical_Operator_out9145_out1;

  Logical_Operator_out10938_out1 <= Logical_Operator_out8634_out1 XOR Logical_Operator_out9146_out1;

  Logical_Operator_out10939_out1 <= Logical_Operator_out8635_out1 XOR Logical_Operator_out9147_out1;

  Logical_Operator_out10940_out1 <= Logical_Operator_out8636_out1 XOR Logical_Operator_out9148_out1;

  Logical_Operator_out10941_out1 <= Logical_Operator_out8637_out1 XOR Logical_Operator_out9149_out1;

  Logical_Operator_out10942_out1 <= Logical_Operator_out8638_out1 XOR Logical_Operator_out9150_out1;

  Logical_Operator_out10943_out1 <= Logical_Operator_out8639_out1 XOR Logical_Operator_out9151_out1;

  Logical_Operator_out10944_out1 <= Logical_Operator_out8640_out1 XOR Logical_Operator_out9152_out1;

  Logical_Operator_out10945_out1 <= Logical_Operator_out8641_out1 XOR Logical_Operator_out9153_out1;

  Logical_Operator_out10946_out1 <= Logical_Operator_out8642_out1 XOR Logical_Operator_out9154_out1;

  Logical_Operator_out10947_out1 <= Logical_Operator_out8643_out1 XOR Logical_Operator_out9155_out1;

  Logical_Operator_out10948_out1 <= Logical_Operator_out8644_out1 XOR Logical_Operator_out9156_out1;

  Logical_Operator_out10949_out1 <= Logical_Operator_out8645_out1 XOR Logical_Operator_out9157_out1;

  Logical_Operator_out10950_out1 <= Logical_Operator_out8646_out1 XOR Logical_Operator_out9158_out1;

  Logical_Operator_out10951_out1 <= Logical_Operator_out8647_out1 XOR Logical_Operator_out9159_out1;

  Logical_Operator_out10952_out1 <= Logical_Operator_out8648_out1 XOR Logical_Operator_out9160_out1;

  Logical_Operator_out10953_out1 <= Logical_Operator_out8649_out1 XOR Logical_Operator_out9161_out1;

  Logical_Operator_out10954_out1 <= Logical_Operator_out8650_out1 XOR Logical_Operator_out9162_out1;

  Logical_Operator_out10955_out1 <= Logical_Operator_out8651_out1 XOR Logical_Operator_out9163_out1;

  Logical_Operator_out10956_out1 <= Logical_Operator_out8652_out1 XOR Logical_Operator_out9164_out1;

  Logical_Operator_out10957_out1 <= Logical_Operator_out8653_out1 XOR Logical_Operator_out9165_out1;

  Logical_Operator_out10958_out1 <= Logical_Operator_out8654_out1 XOR Logical_Operator_out9166_out1;

  Logical_Operator_out10959_out1 <= Logical_Operator_out8655_out1 XOR Logical_Operator_out9167_out1;

  Logical_Operator_out10960_out1 <= Logical_Operator_out8656_out1 XOR Logical_Operator_out9168_out1;

  Logical_Operator_out10961_out1 <= Logical_Operator_out8657_out1 XOR Logical_Operator_out9169_out1;

  Logical_Operator_out10962_out1 <= Logical_Operator_out8658_out1 XOR Logical_Operator_out9170_out1;

  Logical_Operator_out10963_out1 <= Logical_Operator_out8659_out1 XOR Logical_Operator_out9171_out1;

  Logical_Operator_out10964_out1 <= Logical_Operator_out8660_out1 XOR Logical_Operator_out9172_out1;

  Logical_Operator_out10965_out1 <= Logical_Operator_out8661_out1 XOR Logical_Operator_out9173_out1;

  Logical_Operator_out10966_out1 <= Logical_Operator_out8662_out1 XOR Logical_Operator_out9174_out1;

  Logical_Operator_out10967_out1 <= Logical_Operator_out8663_out1 XOR Logical_Operator_out9175_out1;

  Logical_Operator_out10968_out1 <= Logical_Operator_out8664_out1 XOR Logical_Operator_out9176_out1;

  Logical_Operator_out10969_out1 <= Logical_Operator_out8665_out1 XOR Logical_Operator_out9177_out1;

  Logical_Operator_out10970_out1 <= Logical_Operator_out8666_out1 XOR Logical_Operator_out9178_out1;

  Logical_Operator_out10971_out1 <= Logical_Operator_out8667_out1 XOR Logical_Operator_out9179_out1;

  Logical_Operator_out10972_out1 <= Logical_Operator_out8668_out1 XOR Logical_Operator_out9180_out1;

  Logical_Operator_out10973_out1 <= Logical_Operator_out8669_out1 XOR Logical_Operator_out9181_out1;

  Logical_Operator_out10974_out1 <= Logical_Operator_out8670_out1 XOR Logical_Operator_out9182_out1;

  Logical_Operator_out10975_out1 <= Logical_Operator_out8671_out1 XOR Logical_Operator_out9183_out1;

  Logical_Operator_out10976_out1 <= Logical_Operator_out8672_out1 XOR Logical_Operator_out9184_out1;

  Logical_Operator_out10977_out1 <= Logical_Operator_out8673_out1 XOR Logical_Operator_out9185_out1;

  Logical_Operator_out10978_out1 <= Logical_Operator_out8674_out1 XOR Logical_Operator_out9186_out1;

  Logical_Operator_out10979_out1 <= Logical_Operator_out8675_out1 XOR Logical_Operator_out9187_out1;

  Logical_Operator_out10980_out1 <= Logical_Operator_out8676_out1 XOR Logical_Operator_out9188_out1;

  Logical_Operator_out10981_out1 <= Logical_Operator_out8677_out1 XOR Logical_Operator_out9189_out1;

  Logical_Operator_out10982_out1 <= Logical_Operator_out8678_out1 XOR Logical_Operator_out9190_out1;

  Logical_Operator_out10983_out1 <= Logical_Operator_out8679_out1 XOR Logical_Operator_out9191_out1;

  Logical_Operator_out10984_out1 <= Logical_Operator_out8680_out1 XOR Logical_Operator_out9192_out1;

  Logical_Operator_out10985_out1 <= Logical_Operator_out8681_out1 XOR Logical_Operator_out9193_out1;

  Logical_Operator_out10986_out1 <= Logical_Operator_out8682_out1 XOR Logical_Operator_out9194_out1;

  Logical_Operator_out10987_out1 <= Logical_Operator_out8683_out1 XOR Logical_Operator_out9195_out1;

  Logical_Operator_out10988_out1 <= Logical_Operator_out8684_out1 XOR Logical_Operator_out9196_out1;

  Logical_Operator_out10989_out1 <= Logical_Operator_out8685_out1 XOR Logical_Operator_out9197_out1;

  Logical_Operator_out10990_out1 <= Logical_Operator_out8686_out1 XOR Logical_Operator_out9198_out1;

  Logical_Operator_out10991_out1 <= Logical_Operator_out8687_out1 XOR Logical_Operator_out9199_out1;

  Logical_Operator_out10992_out1 <= Logical_Operator_out8688_out1 XOR Logical_Operator_out9200_out1;

  Logical_Operator_out10993_out1 <= Logical_Operator_out8689_out1 XOR Logical_Operator_out9201_out1;

  Logical_Operator_out10994_out1 <= Logical_Operator_out8690_out1 XOR Logical_Operator_out9202_out1;

  Logical_Operator_out10995_out1 <= Logical_Operator_out8691_out1 XOR Logical_Operator_out9203_out1;

  Logical_Operator_out10996_out1 <= Logical_Operator_out8692_out1 XOR Logical_Operator_out9204_out1;

  Logical_Operator_out10997_out1 <= Logical_Operator_out8693_out1 XOR Logical_Operator_out9205_out1;

  Logical_Operator_out10998_out1 <= Logical_Operator_out8694_out1 XOR Logical_Operator_out9206_out1;

  Logical_Operator_out10999_out1 <= Logical_Operator_out8695_out1 XOR Logical_Operator_out9207_out1;

  Logical_Operator_out11000_out1 <= Logical_Operator_out8696_out1 XOR Logical_Operator_out9208_out1;

  Logical_Operator_out11001_out1 <= Logical_Operator_out8697_out1 XOR Logical_Operator_out9209_out1;

  Logical_Operator_out11002_out1 <= Logical_Operator_out8698_out1 XOR Logical_Operator_out9210_out1;

  Logical_Operator_out11003_out1 <= Logical_Operator_out8699_out1 XOR Logical_Operator_out9211_out1;

  Logical_Operator_out11004_out1 <= Logical_Operator_out8700_out1 XOR Logical_Operator_out9212_out1;

  Logical_Operator_out11005_out1 <= Logical_Operator_out8701_out1 XOR Logical_Operator_out9213_out1;

  Logical_Operator_out11006_out1 <= Logical_Operator_out8702_out1 XOR Logical_Operator_out9214_out1;

  Logical_Operator_out11007_out1 <= Logical_Operator_out8703_out1 XOR Logical_Operator_out9215_out1;

  Logical_Operator_out11008_out1 <= Logical_Operator_out8704_out1 XOR Logical_Operator_out9216_out1;

  Logical_Operator_out11009_out1 <= Logical_Operator_out7553_out1 XOR Logical_Operator_out8065_out1;

  Logical_Operator_out11010_out1 <= Logical_Operator_out7554_out1 XOR Logical_Operator_out8066_out1;

  Logical_Operator_out11011_out1 <= Logical_Operator_out7555_out1 XOR Logical_Operator_out8067_out1;

  Logical_Operator_out11012_out1 <= Logical_Operator_out7556_out1 XOR Logical_Operator_out8068_out1;

  Logical_Operator_out11013_out1 <= Logical_Operator_out7557_out1 XOR Logical_Operator_out8069_out1;

  Logical_Operator_out11014_out1 <= Logical_Operator_out7558_out1 XOR Logical_Operator_out8070_out1;

  Logical_Operator_out11015_out1 <= Logical_Operator_out7559_out1 XOR Logical_Operator_out8071_out1;

  Logical_Operator_out11016_out1 <= Logical_Operator_out7560_out1 XOR Logical_Operator_out8072_out1;

  Logical_Operator_out11017_out1 <= Logical_Operator_out7561_out1 XOR Logical_Operator_out8073_out1;

  Logical_Operator_out11018_out1 <= Logical_Operator_out7562_out1 XOR Logical_Operator_out8074_out1;

  Logical_Operator_out11019_out1 <= Logical_Operator_out7563_out1 XOR Logical_Operator_out8075_out1;

  Logical_Operator_out11020_out1 <= Logical_Operator_out7564_out1 XOR Logical_Operator_out8076_out1;

  Logical_Operator_out11021_out1 <= Logical_Operator_out7565_out1 XOR Logical_Operator_out8077_out1;

  Logical_Operator_out11022_out1 <= Logical_Operator_out7566_out1 XOR Logical_Operator_out8078_out1;

  Logical_Operator_out11023_out1 <= Logical_Operator_out7567_out1 XOR Logical_Operator_out8079_out1;

  Logical_Operator_out11024_out1 <= Logical_Operator_out7568_out1 XOR Logical_Operator_out8080_out1;

  Logical_Operator_out11025_out1 <= Logical_Operator_out7569_out1 XOR Logical_Operator_out8081_out1;

  Logical_Operator_out11026_out1 <= Logical_Operator_out7570_out1 XOR Logical_Operator_out8082_out1;

  Logical_Operator_out11027_out1 <= Logical_Operator_out7571_out1 XOR Logical_Operator_out8083_out1;

  Logical_Operator_out11028_out1 <= Logical_Operator_out7572_out1 XOR Logical_Operator_out8084_out1;

  Logical_Operator_out11029_out1 <= Logical_Operator_out7573_out1 XOR Logical_Operator_out8085_out1;

  Logical_Operator_out11030_out1 <= Logical_Operator_out7574_out1 XOR Logical_Operator_out8086_out1;

  Logical_Operator_out11031_out1 <= Logical_Operator_out7575_out1 XOR Logical_Operator_out8087_out1;

  Logical_Operator_out11032_out1 <= Logical_Operator_out7576_out1 XOR Logical_Operator_out8088_out1;

  Logical_Operator_out11033_out1 <= Logical_Operator_out7577_out1 XOR Logical_Operator_out8089_out1;

  Logical_Operator_out11034_out1 <= Logical_Operator_out7578_out1 XOR Logical_Operator_out8090_out1;

  Logical_Operator_out11035_out1 <= Logical_Operator_out7579_out1 XOR Logical_Operator_out8091_out1;

  Logical_Operator_out11036_out1 <= Logical_Operator_out7580_out1 XOR Logical_Operator_out8092_out1;

  Logical_Operator_out11037_out1 <= Logical_Operator_out7581_out1 XOR Logical_Operator_out8093_out1;

  Logical_Operator_out11038_out1 <= Logical_Operator_out7582_out1 XOR Logical_Operator_out8094_out1;

  Logical_Operator_out11039_out1 <= Logical_Operator_out7583_out1 XOR Logical_Operator_out8095_out1;

  Logical_Operator_out11040_out1 <= Logical_Operator_out7584_out1 XOR Logical_Operator_out8096_out1;

  Logical_Operator_out11041_out1 <= Logical_Operator_out7585_out1 XOR Logical_Operator_out8097_out1;

  Logical_Operator_out11042_out1 <= Logical_Operator_out7586_out1 XOR Logical_Operator_out8098_out1;

  Logical_Operator_out11043_out1 <= Logical_Operator_out7587_out1 XOR Logical_Operator_out8099_out1;

  Logical_Operator_out11044_out1 <= Logical_Operator_out7588_out1 XOR Logical_Operator_out8100_out1;

  Logical_Operator_out11045_out1 <= Logical_Operator_out7589_out1 XOR Logical_Operator_out8101_out1;

  Logical_Operator_out11046_out1 <= Logical_Operator_out7590_out1 XOR Logical_Operator_out8102_out1;

  Logical_Operator_out11047_out1 <= Logical_Operator_out7591_out1 XOR Logical_Operator_out8103_out1;

  Logical_Operator_out11048_out1 <= Logical_Operator_out7592_out1 XOR Logical_Operator_out8104_out1;

  Logical_Operator_out11049_out1 <= Logical_Operator_out7593_out1 XOR Logical_Operator_out8105_out1;

  Logical_Operator_out11050_out1 <= Logical_Operator_out7594_out1 XOR Logical_Operator_out8106_out1;

  Logical_Operator_out11051_out1 <= Logical_Operator_out7595_out1 XOR Logical_Operator_out8107_out1;

  Logical_Operator_out11052_out1 <= Logical_Operator_out7596_out1 XOR Logical_Operator_out8108_out1;

  Logical_Operator_out11053_out1 <= Logical_Operator_out7597_out1 XOR Logical_Operator_out8109_out1;

  Logical_Operator_out11054_out1 <= Logical_Operator_out7598_out1 XOR Logical_Operator_out8110_out1;

  Logical_Operator_out11055_out1 <= Logical_Operator_out7599_out1 XOR Logical_Operator_out8111_out1;

  Logical_Operator_out11056_out1 <= Logical_Operator_out7600_out1 XOR Logical_Operator_out8112_out1;

  Logical_Operator_out11057_out1 <= Logical_Operator_out7601_out1 XOR Logical_Operator_out8113_out1;

  Logical_Operator_out11058_out1 <= Logical_Operator_out7602_out1 XOR Logical_Operator_out8114_out1;

  Logical_Operator_out11059_out1 <= Logical_Operator_out7603_out1 XOR Logical_Operator_out8115_out1;

  Logical_Operator_out11060_out1 <= Logical_Operator_out7604_out1 XOR Logical_Operator_out8116_out1;

  Logical_Operator_out11061_out1 <= Logical_Operator_out7605_out1 XOR Logical_Operator_out8117_out1;

  Logical_Operator_out11062_out1 <= Logical_Operator_out7606_out1 XOR Logical_Operator_out8118_out1;

  Logical_Operator_out11063_out1 <= Logical_Operator_out7607_out1 XOR Logical_Operator_out8119_out1;

  Logical_Operator_out11064_out1 <= Logical_Operator_out7608_out1 XOR Logical_Operator_out8120_out1;

  Logical_Operator_out11065_out1 <= Logical_Operator_out7609_out1 XOR Logical_Operator_out8121_out1;

  Logical_Operator_out11066_out1 <= Logical_Operator_out7610_out1 XOR Logical_Operator_out8122_out1;

  Logical_Operator_out11067_out1 <= Logical_Operator_out7611_out1 XOR Logical_Operator_out8123_out1;

  Logical_Operator_out11068_out1 <= Logical_Operator_out7612_out1 XOR Logical_Operator_out8124_out1;

  Logical_Operator_out11069_out1 <= Logical_Operator_out7613_out1 XOR Logical_Operator_out8125_out1;

  Logical_Operator_out11070_out1 <= Logical_Operator_out7614_out1 XOR Logical_Operator_out8126_out1;

  Logical_Operator_out11071_out1 <= Logical_Operator_out7615_out1 XOR Logical_Operator_out8127_out1;

  Logical_Operator_out11072_out1 <= Logical_Operator_out7616_out1 XOR Logical_Operator_out8128_out1;

  Logical_Operator_out11073_out1 <= Logical_Operator_out7617_out1 XOR Logical_Operator_out8129_out1;

  Logical_Operator_out11074_out1 <= Logical_Operator_out7618_out1 XOR Logical_Operator_out8130_out1;

  Logical_Operator_out11075_out1 <= Logical_Operator_out7619_out1 XOR Logical_Operator_out8131_out1;

  Logical_Operator_out11076_out1 <= Logical_Operator_out7620_out1 XOR Logical_Operator_out8132_out1;

  Logical_Operator_out11077_out1 <= Logical_Operator_out7621_out1 XOR Logical_Operator_out8133_out1;

  Logical_Operator_out11078_out1 <= Logical_Operator_out7622_out1 XOR Logical_Operator_out8134_out1;

  Logical_Operator_out11079_out1 <= Logical_Operator_out7623_out1 XOR Logical_Operator_out8135_out1;

  Logical_Operator_out11080_out1 <= Logical_Operator_out7624_out1 XOR Logical_Operator_out8136_out1;

  Logical_Operator_out11081_out1 <= Logical_Operator_out7625_out1 XOR Logical_Operator_out8137_out1;

  Logical_Operator_out11082_out1 <= Logical_Operator_out7626_out1 XOR Logical_Operator_out8138_out1;

  Logical_Operator_out11083_out1 <= Logical_Operator_out7627_out1 XOR Logical_Operator_out8139_out1;

  Logical_Operator_out11084_out1 <= Logical_Operator_out7628_out1 XOR Logical_Operator_out8140_out1;

  Logical_Operator_out11085_out1 <= Logical_Operator_out7629_out1 XOR Logical_Operator_out8141_out1;

  Logical_Operator_out11086_out1 <= Logical_Operator_out7630_out1 XOR Logical_Operator_out8142_out1;

  Logical_Operator_out11087_out1 <= Logical_Operator_out7631_out1 XOR Logical_Operator_out8143_out1;

  Logical_Operator_out11088_out1 <= Logical_Operator_out7632_out1 XOR Logical_Operator_out8144_out1;

  Logical_Operator_out11089_out1 <= Logical_Operator_out7633_out1 XOR Logical_Operator_out8145_out1;

  Logical_Operator_out11090_out1 <= Logical_Operator_out7634_out1 XOR Logical_Operator_out8146_out1;

  Logical_Operator_out11091_out1 <= Logical_Operator_out7635_out1 XOR Logical_Operator_out8147_out1;

  Logical_Operator_out11092_out1 <= Logical_Operator_out7636_out1 XOR Logical_Operator_out8148_out1;

  Logical_Operator_out11093_out1 <= Logical_Operator_out7637_out1 XOR Logical_Operator_out8149_out1;

  Logical_Operator_out11094_out1 <= Logical_Operator_out7638_out1 XOR Logical_Operator_out8150_out1;

  Logical_Operator_out11095_out1 <= Logical_Operator_out7639_out1 XOR Logical_Operator_out8151_out1;

  Logical_Operator_out11096_out1 <= Logical_Operator_out7640_out1 XOR Logical_Operator_out8152_out1;

  Logical_Operator_out11097_out1 <= Logical_Operator_out7641_out1 XOR Logical_Operator_out8153_out1;

  Logical_Operator_out11098_out1 <= Logical_Operator_out7642_out1 XOR Logical_Operator_out8154_out1;

  Logical_Operator_out11099_out1 <= Logical_Operator_out7643_out1 XOR Logical_Operator_out8155_out1;

  Logical_Operator_out11100_out1 <= Logical_Operator_out7644_out1 XOR Logical_Operator_out8156_out1;

  Logical_Operator_out11101_out1 <= Logical_Operator_out7645_out1 XOR Logical_Operator_out8157_out1;

  Logical_Operator_out11102_out1 <= Logical_Operator_out7646_out1 XOR Logical_Operator_out8158_out1;

  Logical_Operator_out11103_out1 <= Logical_Operator_out7647_out1 XOR Logical_Operator_out8159_out1;

  Logical_Operator_out11104_out1 <= Logical_Operator_out7648_out1 XOR Logical_Operator_out8160_out1;

  Logical_Operator_out11105_out1 <= Logical_Operator_out7649_out1 XOR Logical_Operator_out8161_out1;

  Logical_Operator_out11106_out1 <= Logical_Operator_out7650_out1 XOR Logical_Operator_out8162_out1;

  Logical_Operator_out11107_out1 <= Logical_Operator_out7651_out1 XOR Logical_Operator_out8163_out1;

  Logical_Operator_out11108_out1 <= Logical_Operator_out7652_out1 XOR Logical_Operator_out8164_out1;

  Logical_Operator_out11109_out1 <= Logical_Operator_out7653_out1 XOR Logical_Operator_out8165_out1;

  Logical_Operator_out11110_out1 <= Logical_Operator_out7654_out1 XOR Logical_Operator_out8166_out1;

  Logical_Operator_out11111_out1 <= Logical_Operator_out7655_out1 XOR Logical_Operator_out8167_out1;

  Logical_Operator_out11112_out1 <= Logical_Operator_out7656_out1 XOR Logical_Operator_out8168_out1;

  Logical_Operator_out11113_out1 <= Logical_Operator_out7657_out1 XOR Logical_Operator_out8169_out1;

  Logical_Operator_out11114_out1 <= Logical_Operator_out7658_out1 XOR Logical_Operator_out8170_out1;

  Logical_Operator_out11115_out1 <= Logical_Operator_out7659_out1 XOR Logical_Operator_out8171_out1;

  Logical_Operator_out11116_out1 <= Logical_Operator_out7660_out1 XOR Logical_Operator_out8172_out1;

  Logical_Operator_out11117_out1 <= Logical_Operator_out7661_out1 XOR Logical_Operator_out8173_out1;

  Logical_Operator_out11118_out1 <= Logical_Operator_out7662_out1 XOR Logical_Operator_out8174_out1;

  Logical_Operator_out11119_out1 <= Logical_Operator_out7663_out1 XOR Logical_Operator_out8175_out1;

  Logical_Operator_out11120_out1 <= Logical_Operator_out7664_out1 XOR Logical_Operator_out8176_out1;

  Logical_Operator_out11121_out1 <= Logical_Operator_out7665_out1 XOR Logical_Operator_out8177_out1;

  Logical_Operator_out11122_out1 <= Logical_Operator_out7666_out1 XOR Logical_Operator_out8178_out1;

  Logical_Operator_out11123_out1 <= Logical_Operator_out7667_out1 XOR Logical_Operator_out8179_out1;

  Logical_Operator_out11124_out1 <= Logical_Operator_out7668_out1 XOR Logical_Operator_out8180_out1;

  Logical_Operator_out11125_out1 <= Logical_Operator_out7669_out1 XOR Logical_Operator_out8181_out1;

  Logical_Operator_out11126_out1 <= Logical_Operator_out7670_out1 XOR Logical_Operator_out8182_out1;

  Logical_Operator_out11127_out1 <= Logical_Operator_out7671_out1 XOR Logical_Operator_out8183_out1;

  Logical_Operator_out11128_out1 <= Logical_Operator_out7672_out1 XOR Logical_Operator_out8184_out1;

  Logical_Operator_out11129_out1 <= Logical_Operator_out7673_out1 XOR Logical_Operator_out8185_out1;

  Logical_Operator_out11130_out1 <= Logical_Operator_out7674_out1 XOR Logical_Operator_out8186_out1;

  Logical_Operator_out11131_out1 <= Logical_Operator_out7675_out1 XOR Logical_Operator_out8187_out1;

  Logical_Operator_out11132_out1 <= Logical_Operator_out7676_out1 XOR Logical_Operator_out8188_out1;

  Logical_Operator_out11133_out1 <= Logical_Operator_out7677_out1 XOR Logical_Operator_out8189_out1;

  Logical_Operator_out11134_out1 <= Logical_Operator_out7678_out1 XOR Logical_Operator_out8190_out1;

  Logical_Operator_out11135_out1 <= Logical_Operator_out7679_out1 XOR Logical_Operator_out8191_out1;

  Logical_Operator_out11136_out1 <= Logical_Operator_out7680_out1 XOR Logical_Operator_out8192_out1;

  Logical_Operator_out11137_out1 <= Logical_Operator_out6593_out1 XOR Logical_Operator_out7105_out1;

  Logical_Operator_out11138_out1 <= Logical_Operator_out6594_out1 XOR Logical_Operator_out7106_out1;

  Logical_Operator_out11139_out1 <= Logical_Operator_out6595_out1 XOR Logical_Operator_out7107_out1;

  Logical_Operator_out11140_out1 <= Logical_Operator_out6596_out1 XOR Logical_Operator_out7108_out1;

  Logical_Operator_out11141_out1 <= Logical_Operator_out6597_out1 XOR Logical_Operator_out7109_out1;

  Logical_Operator_out11142_out1 <= Logical_Operator_out6598_out1 XOR Logical_Operator_out7110_out1;

  Logical_Operator_out11143_out1 <= Logical_Operator_out6599_out1 XOR Logical_Operator_out7111_out1;

  Logical_Operator_out11144_out1 <= Logical_Operator_out6600_out1 XOR Logical_Operator_out7112_out1;

  Logical_Operator_out11145_out1 <= Logical_Operator_out6601_out1 XOR Logical_Operator_out7113_out1;

  Logical_Operator_out11146_out1 <= Logical_Operator_out6602_out1 XOR Logical_Operator_out7114_out1;

  Logical_Operator_out11147_out1 <= Logical_Operator_out6603_out1 XOR Logical_Operator_out7115_out1;

  Logical_Operator_out11148_out1 <= Logical_Operator_out6604_out1 XOR Logical_Operator_out7116_out1;

  Logical_Operator_out11149_out1 <= Logical_Operator_out6605_out1 XOR Logical_Operator_out7117_out1;

  Logical_Operator_out11150_out1 <= Logical_Operator_out6606_out1 XOR Logical_Operator_out7118_out1;

  Logical_Operator_out11151_out1 <= Logical_Operator_out6607_out1 XOR Logical_Operator_out7119_out1;

  Logical_Operator_out11152_out1 <= Logical_Operator_out6608_out1 XOR Logical_Operator_out7120_out1;

  Logical_Operator_out11153_out1 <= Logical_Operator_out6609_out1 XOR Logical_Operator_out7121_out1;

  Logical_Operator_out11154_out1 <= Logical_Operator_out6610_out1 XOR Logical_Operator_out7122_out1;

  Logical_Operator_out11155_out1 <= Logical_Operator_out6611_out1 XOR Logical_Operator_out7123_out1;

  Logical_Operator_out11156_out1 <= Logical_Operator_out6612_out1 XOR Logical_Operator_out7124_out1;

  Logical_Operator_out11157_out1 <= Logical_Operator_out6613_out1 XOR Logical_Operator_out7125_out1;

  Logical_Operator_out11158_out1 <= Logical_Operator_out6614_out1 XOR Logical_Operator_out7126_out1;

  Logical_Operator_out11159_out1 <= Logical_Operator_out6615_out1 XOR Logical_Operator_out7127_out1;

  Logical_Operator_out11160_out1 <= Logical_Operator_out6616_out1 XOR Logical_Operator_out7128_out1;

  Logical_Operator_out11161_out1 <= Logical_Operator_out6617_out1 XOR Logical_Operator_out7129_out1;

  Logical_Operator_out11162_out1 <= Logical_Operator_out6618_out1 XOR Logical_Operator_out7130_out1;

  Logical_Operator_out11163_out1 <= Logical_Operator_out6619_out1 XOR Logical_Operator_out7131_out1;

  Logical_Operator_out11164_out1 <= Logical_Operator_out6620_out1 XOR Logical_Operator_out7132_out1;

  Logical_Operator_out11165_out1 <= Logical_Operator_out6621_out1 XOR Logical_Operator_out7133_out1;

  Logical_Operator_out11166_out1 <= Logical_Operator_out6622_out1 XOR Logical_Operator_out7134_out1;

  Logical_Operator_out11167_out1 <= Logical_Operator_out6623_out1 XOR Logical_Operator_out7135_out1;

  Logical_Operator_out11168_out1 <= Logical_Operator_out6624_out1 XOR Logical_Operator_out7136_out1;

  Logical_Operator_out11169_out1 <= Logical_Operator_out6625_out1 XOR Logical_Operator_out7137_out1;

  Logical_Operator_out11170_out1 <= Logical_Operator_out6626_out1 XOR Logical_Operator_out7138_out1;

  Logical_Operator_out11171_out1 <= Logical_Operator_out6627_out1 XOR Logical_Operator_out7139_out1;

  Logical_Operator_out11172_out1 <= Logical_Operator_out6628_out1 XOR Logical_Operator_out7140_out1;

  Logical_Operator_out11173_out1 <= Logical_Operator_out6629_out1 XOR Logical_Operator_out7141_out1;

  Logical_Operator_out11174_out1 <= Logical_Operator_out6630_out1 XOR Logical_Operator_out7142_out1;

  Logical_Operator_out11175_out1 <= Logical_Operator_out6631_out1 XOR Logical_Operator_out7143_out1;

  Logical_Operator_out11176_out1 <= Logical_Operator_out6632_out1 XOR Logical_Operator_out7144_out1;

  Logical_Operator_out11177_out1 <= Logical_Operator_out6633_out1 XOR Logical_Operator_out7145_out1;

  Logical_Operator_out11178_out1 <= Logical_Operator_out6634_out1 XOR Logical_Operator_out7146_out1;

  Logical_Operator_out11179_out1 <= Logical_Operator_out6635_out1 XOR Logical_Operator_out7147_out1;

  Logical_Operator_out11180_out1 <= Logical_Operator_out6636_out1 XOR Logical_Operator_out7148_out1;

  Logical_Operator_out11181_out1 <= Logical_Operator_out6637_out1 XOR Logical_Operator_out7149_out1;

  Logical_Operator_out11182_out1 <= Logical_Operator_out6638_out1 XOR Logical_Operator_out7150_out1;

  Logical_Operator_out11183_out1 <= Logical_Operator_out6639_out1 XOR Logical_Operator_out7151_out1;

  Logical_Operator_out11184_out1 <= Logical_Operator_out6640_out1 XOR Logical_Operator_out7152_out1;

  Logical_Operator_out11185_out1 <= Logical_Operator_out6641_out1 XOR Logical_Operator_out7153_out1;

  Logical_Operator_out11186_out1 <= Logical_Operator_out6642_out1 XOR Logical_Operator_out7154_out1;

  Logical_Operator_out11187_out1 <= Logical_Operator_out6643_out1 XOR Logical_Operator_out7155_out1;

  Logical_Operator_out11188_out1 <= Logical_Operator_out6644_out1 XOR Logical_Operator_out7156_out1;

  Logical_Operator_out11189_out1 <= Logical_Operator_out6645_out1 XOR Logical_Operator_out7157_out1;

  Logical_Operator_out11190_out1 <= Logical_Operator_out6646_out1 XOR Logical_Operator_out7158_out1;

  Logical_Operator_out11191_out1 <= Logical_Operator_out6647_out1 XOR Logical_Operator_out7159_out1;

  Logical_Operator_out11192_out1 <= Logical_Operator_out6648_out1 XOR Logical_Operator_out7160_out1;

  Logical_Operator_out11193_out1 <= Logical_Operator_out6649_out1 XOR Logical_Operator_out7161_out1;

  Logical_Operator_out11194_out1 <= Logical_Operator_out6650_out1 XOR Logical_Operator_out7162_out1;

  Logical_Operator_out11195_out1 <= Logical_Operator_out6651_out1 XOR Logical_Operator_out7163_out1;

  Logical_Operator_out11196_out1 <= Logical_Operator_out6652_out1 XOR Logical_Operator_out7164_out1;

  Logical_Operator_out11197_out1 <= Logical_Operator_out6653_out1 XOR Logical_Operator_out7165_out1;

  Logical_Operator_out11198_out1 <= Logical_Operator_out6654_out1 XOR Logical_Operator_out7166_out1;

  Logical_Operator_out11199_out1 <= Logical_Operator_out6655_out1 XOR Logical_Operator_out7167_out1;

  Logical_Operator_out11200_out1 <= Logical_Operator_out6656_out1 XOR Logical_Operator_out7168_out1;

  Logical_Operator_out11201_out1 <= Logical_Operator_out5601_out1 XOR Logical_Operator_out6113_out1;

  Logical_Operator_out11202_out1 <= Logical_Operator_out5602_out1 XOR Logical_Operator_out6114_out1;

  Logical_Operator_out11203_out1 <= Logical_Operator_out5603_out1 XOR Logical_Operator_out6115_out1;

  Logical_Operator_out11204_out1 <= Logical_Operator_out5604_out1 XOR Logical_Operator_out6116_out1;

  Logical_Operator_out11205_out1 <= Logical_Operator_out5605_out1 XOR Logical_Operator_out6117_out1;

  Logical_Operator_out11206_out1 <= Logical_Operator_out5606_out1 XOR Logical_Operator_out6118_out1;

  Logical_Operator_out11207_out1 <= Logical_Operator_out5607_out1 XOR Logical_Operator_out6119_out1;

  Logical_Operator_out11208_out1 <= Logical_Operator_out5608_out1 XOR Logical_Operator_out6120_out1;

  Logical_Operator_out11209_out1 <= Logical_Operator_out5609_out1 XOR Logical_Operator_out6121_out1;

  Logical_Operator_out11210_out1 <= Logical_Operator_out5610_out1 XOR Logical_Operator_out6122_out1;

  Logical_Operator_out11211_out1 <= Logical_Operator_out5611_out1 XOR Logical_Operator_out6123_out1;

  Logical_Operator_out11212_out1 <= Logical_Operator_out5612_out1 XOR Logical_Operator_out6124_out1;

  Logical_Operator_out11213_out1 <= Logical_Operator_out5613_out1 XOR Logical_Operator_out6125_out1;

  Logical_Operator_out11214_out1 <= Logical_Operator_out5614_out1 XOR Logical_Operator_out6126_out1;

  Logical_Operator_out11215_out1 <= Logical_Operator_out5615_out1 XOR Logical_Operator_out6127_out1;

  Logical_Operator_out11216_out1 <= Logical_Operator_out5616_out1 XOR Logical_Operator_out6128_out1;

  Logical_Operator_out11217_out1 <= Logical_Operator_out5617_out1 XOR Logical_Operator_out6129_out1;

  Logical_Operator_out11218_out1 <= Logical_Operator_out5618_out1 XOR Logical_Operator_out6130_out1;

  Logical_Operator_out11219_out1 <= Logical_Operator_out5619_out1 XOR Logical_Operator_out6131_out1;

  Logical_Operator_out11220_out1 <= Logical_Operator_out5620_out1 XOR Logical_Operator_out6132_out1;

  Logical_Operator_out11221_out1 <= Logical_Operator_out5621_out1 XOR Logical_Operator_out6133_out1;

  Logical_Operator_out11222_out1 <= Logical_Operator_out5622_out1 XOR Logical_Operator_out6134_out1;

  Logical_Operator_out11223_out1 <= Logical_Operator_out5623_out1 XOR Logical_Operator_out6135_out1;

  Logical_Operator_out11224_out1 <= Logical_Operator_out5624_out1 XOR Logical_Operator_out6136_out1;

  Logical_Operator_out11225_out1 <= Logical_Operator_out5625_out1 XOR Logical_Operator_out6137_out1;

  Logical_Operator_out11226_out1 <= Logical_Operator_out5626_out1 XOR Logical_Operator_out6138_out1;

  Logical_Operator_out11227_out1 <= Logical_Operator_out5627_out1 XOR Logical_Operator_out6139_out1;

  Logical_Operator_out11228_out1 <= Logical_Operator_out5628_out1 XOR Logical_Operator_out6140_out1;

  Logical_Operator_out11229_out1 <= Logical_Operator_out5629_out1 XOR Logical_Operator_out6141_out1;

  Logical_Operator_out11230_out1 <= Logical_Operator_out5630_out1 XOR Logical_Operator_out6142_out1;

  Logical_Operator_out11231_out1 <= Logical_Operator_out5631_out1 XOR Logical_Operator_out6143_out1;

  Logical_Operator_out11232_out1 <= Logical_Operator_out5632_out1 XOR Logical_Operator_out6144_out1;

  Logical_Operator_out11233_out1 <= Logical_Operator_out4593_out1 XOR Logical_Operator_out5105_out1;

  Logical_Operator_out11234_out1 <= Logical_Operator_out4594_out1 XOR Logical_Operator_out5106_out1;

  Logical_Operator_out11235_out1 <= Logical_Operator_out4595_out1 XOR Logical_Operator_out5107_out1;

  Logical_Operator_out11236_out1 <= Logical_Operator_out4596_out1 XOR Logical_Operator_out5108_out1;

  Logical_Operator_out11237_out1 <= Logical_Operator_out4597_out1 XOR Logical_Operator_out5109_out1;

  Logical_Operator_out11238_out1 <= Logical_Operator_out4598_out1 XOR Logical_Operator_out5110_out1;

  Logical_Operator_out11239_out1 <= Logical_Operator_out4599_out1 XOR Logical_Operator_out5111_out1;

  Logical_Operator_out11240_out1 <= Logical_Operator_out4600_out1 XOR Logical_Operator_out5112_out1;

  Logical_Operator_out11241_out1 <= Logical_Operator_out4601_out1 XOR Logical_Operator_out5113_out1;

  Logical_Operator_out11242_out1 <= Logical_Operator_out4602_out1 XOR Logical_Operator_out5114_out1;

  Logical_Operator_out11243_out1 <= Logical_Operator_out4603_out1 XOR Logical_Operator_out5115_out1;

  Logical_Operator_out11244_out1 <= Logical_Operator_out4604_out1 XOR Logical_Operator_out5116_out1;

  Logical_Operator_out11245_out1 <= Logical_Operator_out4605_out1 XOR Logical_Operator_out5117_out1;

  Logical_Operator_out11246_out1 <= Logical_Operator_out4606_out1 XOR Logical_Operator_out5118_out1;

  Logical_Operator_out11247_out1 <= Logical_Operator_out4607_out1 XOR Logical_Operator_out5119_out1;

  Logical_Operator_out11248_out1 <= Logical_Operator_out4608_out1 XOR Logical_Operator_out5120_out1;

  Logical_Operator_out11249_out1 <= Logical_Operator_out3577_out1 XOR Logical_Operator_out4089_out1;

  Logical_Operator_out11250_out1 <= Logical_Operator_out3578_out1 XOR Logical_Operator_out4090_out1;

  Logical_Operator_out11251_out1 <= Logical_Operator_out3579_out1 XOR Logical_Operator_out4091_out1;

  Logical_Operator_out11252_out1 <= Logical_Operator_out3580_out1 XOR Logical_Operator_out4092_out1;

  Logical_Operator_out11253_out1 <= Logical_Operator_out3581_out1 XOR Logical_Operator_out4093_out1;

  Logical_Operator_out11254_out1 <= Logical_Operator_out3582_out1 XOR Logical_Operator_out4094_out1;

  Logical_Operator_out11255_out1 <= Logical_Operator_out3583_out1 XOR Logical_Operator_out4095_out1;

  Logical_Operator_out11256_out1 <= Logical_Operator_out3584_out1 XOR Logical_Operator_out4096_out1;

  Logical_Operator_out11257_out1 <= Logical_Operator_out2557_out1 XOR Logical_Operator_out3069_out1;

  Logical_Operator_out11258_out1 <= Logical_Operator_out2558_out1 XOR Logical_Operator_out3070_out1;

  Logical_Operator_out11259_out1 <= Logical_Operator_out2559_out1 XOR Logical_Operator_out3071_out1;

  Logical_Operator_out11260_out1 <= Logical_Operator_out2560_out1 XOR Logical_Operator_out3072_out1;

  Logical_Operator_out11261_out1 <= Logical_Operator_out1535_out1 XOR Logical_Operator_out2047_out1;

  Logical_Operator_out11262_out1 <= Logical_Operator_out1536_out1 XOR Logical_Operator_out2048_out1;

  Logical_Operator_out11263_out1 <= Logical_Operator_out512_out1 XOR Logical_Operator_out1024_out1;

  Logical_Operator_out11264_out1 <= in1024 XOR in2048;

  out1 <= Logical_Operator_out10241_out1;

  out2 <= Logical_Operator_out10242_out1;

  out3 <= Logical_Operator_out10243_out1;

  out4 <= Logical_Operator_out10244_out1;

  out5 <= Logical_Operator_out10245_out1;

  out6 <= Logical_Operator_out10246_out1;

  out7 <= Logical_Operator_out10247_out1;

  out8 <= Logical_Operator_out10248_out1;

  out9 <= Logical_Operator_out10249_out1;

  out10 <= Logical_Operator_out10250_out1;

  out11 <= Logical_Operator_out10251_out1;

  out12 <= Logical_Operator_out10252_out1;

  out13 <= Logical_Operator_out10253_out1;

  out14 <= Logical_Operator_out10254_out1;

  out15 <= Logical_Operator_out10255_out1;

  out16 <= Logical_Operator_out10256_out1;

  out17 <= Logical_Operator_out10257_out1;

  out18 <= Logical_Operator_out10258_out1;

  out19 <= Logical_Operator_out10259_out1;

  out20 <= Logical_Operator_out10260_out1;

  out21 <= Logical_Operator_out10261_out1;

  out22 <= Logical_Operator_out10262_out1;

  out23 <= Logical_Operator_out10263_out1;

  out24 <= Logical_Operator_out10264_out1;

  out25 <= Logical_Operator_out10265_out1;

  out26 <= Logical_Operator_out10266_out1;

  out27 <= Logical_Operator_out10267_out1;

  out28 <= Logical_Operator_out10268_out1;

  out29 <= Logical_Operator_out10269_out1;

  out30 <= Logical_Operator_out10270_out1;

  out31 <= Logical_Operator_out10271_out1;

  out32 <= Logical_Operator_out10272_out1;

  out33 <= Logical_Operator_out10273_out1;

  out34 <= Logical_Operator_out10274_out1;

  out35 <= Logical_Operator_out10275_out1;

  out36 <= Logical_Operator_out10276_out1;

  out37 <= Logical_Operator_out10277_out1;

  out38 <= Logical_Operator_out10278_out1;

  out39 <= Logical_Operator_out10279_out1;

  out40 <= Logical_Operator_out10280_out1;

  out41 <= Logical_Operator_out10281_out1;

  out42 <= Logical_Operator_out10282_out1;

  out43 <= Logical_Operator_out10283_out1;

  out44 <= Logical_Operator_out10284_out1;

  out45 <= Logical_Operator_out10285_out1;

  out46 <= Logical_Operator_out10286_out1;

  out47 <= Logical_Operator_out10287_out1;

  out48 <= Logical_Operator_out10288_out1;

  out49 <= Logical_Operator_out10289_out1;

  out50 <= Logical_Operator_out10290_out1;

  out51 <= Logical_Operator_out10291_out1;

  out52 <= Logical_Operator_out10292_out1;

  out53 <= Logical_Operator_out10293_out1;

  out54 <= Logical_Operator_out10294_out1;

  out55 <= Logical_Operator_out10295_out1;

  out56 <= Logical_Operator_out10296_out1;

  out57 <= Logical_Operator_out10297_out1;

  out58 <= Logical_Operator_out10298_out1;

  out59 <= Logical_Operator_out10299_out1;

  out60 <= Logical_Operator_out10300_out1;

  out61 <= Logical_Operator_out10301_out1;

  out62 <= Logical_Operator_out10302_out1;

  out63 <= Logical_Operator_out10303_out1;

  out64 <= Logical_Operator_out10304_out1;

  out65 <= Logical_Operator_out10305_out1;

  out66 <= Logical_Operator_out10306_out1;

  out67 <= Logical_Operator_out10307_out1;

  out68 <= Logical_Operator_out10308_out1;

  out69 <= Logical_Operator_out10309_out1;

  out70 <= Logical_Operator_out10310_out1;

  out71 <= Logical_Operator_out10311_out1;

  out72 <= Logical_Operator_out10312_out1;

  out73 <= Logical_Operator_out10313_out1;

  out74 <= Logical_Operator_out10314_out1;

  out75 <= Logical_Operator_out10315_out1;

  out76 <= Logical_Operator_out10316_out1;

  out77 <= Logical_Operator_out10317_out1;

  out78 <= Logical_Operator_out10318_out1;

  out79 <= Logical_Operator_out10319_out1;

  out80 <= Logical_Operator_out10320_out1;

  out81 <= Logical_Operator_out10321_out1;

  out82 <= Logical_Operator_out10322_out1;

  out83 <= Logical_Operator_out10323_out1;

  out84 <= Logical_Operator_out10324_out1;

  out85 <= Logical_Operator_out10325_out1;

  out86 <= Logical_Operator_out10326_out1;

  out87 <= Logical_Operator_out10327_out1;

  out88 <= Logical_Operator_out10328_out1;

  out89 <= Logical_Operator_out10329_out1;

  out90 <= Logical_Operator_out10330_out1;

  out91 <= Logical_Operator_out10331_out1;

  out92 <= Logical_Operator_out10332_out1;

  out93 <= Logical_Operator_out10333_out1;

  out94 <= Logical_Operator_out10334_out1;

  out95 <= Logical_Operator_out10335_out1;

  out96 <= Logical_Operator_out10336_out1;

  out97 <= Logical_Operator_out10337_out1;

  out98 <= Logical_Operator_out10338_out1;

  out99 <= Logical_Operator_out10339_out1;

  out100 <= Logical_Operator_out10340_out1;

  out101 <= Logical_Operator_out10341_out1;

  out102 <= Logical_Operator_out10342_out1;

  out103 <= Logical_Operator_out10343_out1;

  out104 <= Logical_Operator_out10344_out1;

  out105 <= Logical_Operator_out10345_out1;

  out106 <= Logical_Operator_out10346_out1;

  out107 <= Logical_Operator_out10347_out1;

  out108 <= Logical_Operator_out10348_out1;

  out109 <= Logical_Operator_out10349_out1;

  out110 <= Logical_Operator_out10350_out1;

  out111 <= Logical_Operator_out10351_out1;

  out112 <= Logical_Operator_out10352_out1;

  out113 <= Logical_Operator_out10353_out1;

  out114 <= Logical_Operator_out10354_out1;

  out115 <= Logical_Operator_out10355_out1;

  out116 <= Logical_Operator_out10356_out1;

  out117 <= Logical_Operator_out10357_out1;

  out118 <= Logical_Operator_out10358_out1;

  out119 <= Logical_Operator_out10359_out1;

  out120 <= Logical_Operator_out10360_out1;

  out121 <= Logical_Operator_out10361_out1;

  out122 <= Logical_Operator_out10362_out1;

  out123 <= Logical_Operator_out10363_out1;

  out124 <= Logical_Operator_out10364_out1;

  out125 <= Logical_Operator_out10365_out1;

  out126 <= Logical_Operator_out10366_out1;

  out127 <= Logical_Operator_out10367_out1;

  out128 <= Logical_Operator_out10368_out1;

  out129 <= Logical_Operator_out10369_out1;

  out130 <= Logical_Operator_out10370_out1;

  out131 <= Logical_Operator_out10371_out1;

  out132 <= Logical_Operator_out10372_out1;

  out133 <= Logical_Operator_out10373_out1;

  out134 <= Logical_Operator_out10374_out1;

  out135 <= Logical_Operator_out10375_out1;

  out136 <= Logical_Operator_out10376_out1;

  out137 <= Logical_Operator_out10377_out1;

  out138 <= Logical_Operator_out10378_out1;

  out139 <= Logical_Operator_out10379_out1;

  out140 <= Logical_Operator_out10380_out1;

  out141 <= Logical_Operator_out10381_out1;

  out142 <= Logical_Operator_out10382_out1;

  out143 <= Logical_Operator_out10383_out1;

  out144 <= Logical_Operator_out10384_out1;

  out145 <= Logical_Operator_out10385_out1;

  out146 <= Logical_Operator_out10386_out1;

  out147 <= Logical_Operator_out10387_out1;

  out148 <= Logical_Operator_out10388_out1;

  out149 <= Logical_Operator_out10389_out1;

  out150 <= Logical_Operator_out10390_out1;

  out151 <= Logical_Operator_out10391_out1;

  out152 <= Logical_Operator_out10392_out1;

  out153 <= Logical_Operator_out10393_out1;

  out154 <= Logical_Operator_out10394_out1;

  out155 <= Logical_Operator_out10395_out1;

  out156 <= Logical_Operator_out10396_out1;

  out157 <= Logical_Operator_out10397_out1;

  out158 <= Logical_Operator_out10398_out1;

  out159 <= Logical_Operator_out10399_out1;

  out160 <= Logical_Operator_out10400_out1;

  out161 <= Logical_Operator_out10401_out1;

  out162 <= Logical_Operator_out10402_out1;

  out163 <= Logical_Operator_out10403_out1;

  out164 <= Logical_Operator_out10404_out1;

  out165 <= Logical_Operator_out10405_out1;

  out166 <= Logical_Operator_out10406_out1;

  out167 <= Logical_Operator_out10407_out1;

  out168 <= Logical_Operator_out10408_out1;

  out169 <= Logical_Operator_out10409_out1;

  out170 <= Logical_Operator_out10410_out1;

  out171 <= Logical_Operator_out10411_out1;

  out172 <= Logical_Operator_out10412_out1;

  out173 <= Logical_Operator_out10413_out1;

  out174 <= Logical_Operator_out10414_out1;

  out175 <= Logical_Operator_out10415_out1;

  out176 <= Logical_Operator_out10416_out1;

  out177 <= Logical_Operator_out10417_out1;

  out178 <= Logical_Operator_out10418_out1;

  out179 <= Logical_Operator_out10419_out1;

  out180 <= Logical_Operator_out10420_out1;

  out181 <= Logical_Operator_out10421_out1;

  out182 <= Logical_Operator_out10422_out1;

  out183 <= Logical_Operator_out10423_out1;

  out184 <= Logical_Operator_out10424_out1;

  out185 <= Logical_Operator_out10425_out1;

  out186 <= Logical_Operator_out10426_out1;

  out187 <= Logical_Operator_out10427_out1;

  out188 <= Logical_Operator_out10428_out1;

  out189 <= Logical_Operator_out10429_out1;

  out190 <= Logical_Operator_out10430_out1;

  out191 <= Logical_Operator_out10431_out1;

  out192 <= Logical_Operator_out10432_out1;

  out193 <= Logical_Operator_out10433_out1;

  out194 <= Logical_Operator_out10434_out1;

  out195 <= Logical_Operator_out10435_out1;

  out196 <= Logical_Operator_out10436_out1;

  out197 <= Logical_Operator_out10437_out1;

  out198 <= Logical_Operator_out10438_out1;

  out199 <= Logical_Operator_out10439_out1;

  out200 <= Logical_Operator_out10440_out1;

  out201 <= Logical_Operator_out10441_out1;

  out202 <= Logical_Operator_out10442_out1;

  out203 <= Logical_Operator_out10443_out1;

  out204 <= Logical_Operator_out10444_out1;

  out205 <= Logical_Operator_out10445_out1;

  out206 <= Logical_Operator_out10446_out1;

  out207 <= Logical_Operator_out10447_out1;

  out208 <= Logical_Operator_out10448_out1;

  out209 <= Logical_Operator_out10449_out1;

  out210 <= Logical_Operator_out10450_out1;

  out211 <= Logical_Operator_out10451_out1;

  out212 <= Logical_Operator_out10452_out1;

  out213 <= Logical_Operator_out10453_out1;

  out214 <= Logical_Operator_out10454_out1;

  out215 <= Logical_Operator_out10455_out1;

  out216 <= Logical_Operator_out10456_out1;

  out217 <= Logical_Operator_out10457_out1;

  out218 <= Logical_Operator_out10458_out1;

  out219 <= Logical_Operator_out10459_out1;

  out220 <= Logical_Operator_out10460_out1;

  out221 <= Logical_Operator_out10461_out1;

  out222 <= Logical_Operator_out10462_out1;

  out223 <= Logical_Operator_out10463_out1;

  out224 <= Logical_Operator_out10464_out1;

  out225 <= Logical_Operator_out10465_out1;

  out226 <= Logical_Operator_out10466_out1;

  out227 <= Logical_Operator_out10467_out1;

  out228 <= Logical_Operator_out10468_out1;

  out229 <= Logical_Operator_out10469_out1;

  out230 <= Logical_Operator_out10470_out1;

  out231 <= Logical_Operator_out10471_out1;

  out232 <= Logical_Operator_out10472_out1;

  out233 <= Logical_Operator_out10473_out1;

  out234 <= Logical_Operator_out10474_out1;

  out235 <= Logical_Operator_out10475_out1;

  out236 <= Logical_Operator_out10476_out1;

  out237 <= Logical_Operator_out10477_out1;

  out238 <= Logical_Operator_out10478_out1;

  out239 <= Logical_Operator_out10479_out1;

  out240 <= Logical_Operator_out10480_out1;

  out241 <= Logical_Operator_out10481_out1;

  out242 <= Logical_Operator_out10482_out1;

  out243 <= Logical_Operator_out10483_out1;

  out244 <= Logical_Operator_out10484_out1;

  out245 <= Logical_Operator_out10485_out1;

  out246 <= Logical_Operator_out10486_out1;

  out247 <= Logical_Operator_out10487_out1;

  out248 <= Logical_Operator_out10488_out1;

  out249 <= Logical_Operator_out10489_out1;

  out250 <= Logical_Operator_out10490_out1;

  out251 <= Logical_Operator_out10491_out1;

  out252 <= Logical_Operator_out10492_out1;

  out253 <= Logical_Operator_out10493_out1;

  out254 <= Logical_Operator_out10494_out1;

  out255 <= Logical_Operator_out10495_out1;

  out256 <= Logical_Operator_out10496_out1;

  out257 <= Logical_Operator_out10497_out1;

  out258 <= Logical_Operator_out10498_out1;

  out259 <= Logical_Operator_out10499_out1;

  out260 <= Logical_Operator_out10500_out1;

  out261 <= Logical_Operator_out10501_out1;

  out262 <= Logical_Operator_out10502_out1;

  out263 <= Logical_Operator_out10503_out1;

  out264 <= Logical_Operator_out10504_out1;

  out265 <= Logical_Operator_out10505_out1;

  out266 <= Logical_Operator_out10506_out1;

  out267 <= Logical_Operator_out10507_out1;

  out268 <= Logical_Operator_out10508_out1;

  out269 <= Logical_Operator_out10509_out1;

  out270 <= Logical_Operator_out10510_out1;

  out271 <= Logical_Operator_out10511_out1;

  out272 <= Logical_Operator_out10512_out1;

  out273 <= Logical_Operator_out10513_out1;

  out274 <= Logical_Operator_out10514_out1;

  out275 <= Logical_Operator_out10515_out1;

  out276 <= Logical_Operator_out10516_out1;

  out277 <= Logical_Operator_out10517_out1;

  out278 <= Logical_Operator_out10518_out1;

  out279 <= Logical_Operator_out10519_out1;

  out280 <= Logical_Operator_out10520_out1;

  out281 <= Logical_Operator_out10521_out1;

  out282 <= Logical_Operator_out10522_out1;

  out283 <= Logical_Operator_out10523_out1;

  out284 <= Logical_Operator_out10524_out1;

  out285 <= Logical_Operator_out10525_out1;

  out286 <= Logical_Operator_out10526_out1;

  out287 <= Logical_Operator_out10527_out1;

  out288 <= Logical_Operator_out10528_out1;

  out289 <= Logical_Operator_out10529_out1;

  out290 <= Logical_Operator_out10530_out1;

  out291 <= Logical_Operator_out10531_out1;

  out292 <= Logical_Operator_out10532_out1;

  out293 <= Logical_Operator_out10533_out1;

  out294 <= Logical_Operator_out10534_out1;

  out295 <= Logical_Operator_out10535_out1;

  out296 <= Logical_Operator_out10536_out1;

  out297 <= Logical_Operator_out10537_out1;

  out298 <= Logical_Operator_out10538_out1;

  out299 <= Logical_Operator_out10539_out1;

  out300 <= Logical_Operator_out10540_out1;

  out301 <= Logical_Operator_out10541_out1;

  out302 <= Logical_Operator_out10542_out1;

  out303 <= Logical_Operator_out10543_out1;

  out304 <= Logical_Operator_out10544_out1;

  out305 <= Logical_Operator_out10545_out1;

  out306 <= Logical_Operator_out10546_out1;

  out307 <= Logical_Operator_out10547_out1;

  out308 <= Logical_Operator_out10548_out1;

  out309 <= Logical_Operator_out10549_out1;

  out310 <= Logical_Operator_out10550_out1;

  out311 <= Logical_Operator_out10551_out1;

  out312 <= Logical_Operator_out10552_out1;

  out313 <= Logical_Operator_out10553_out1;

  out314 <= Logical_Operator_out10554_out1;

  out315 <= Logical_Operator_out10555_out1;

  out316 <= Logical_Operator_out10556_out1;

  out317 <= Logical_Operator_out10557_out1;

  out318 <= Logical_Operator_out10558_out1;

  out319 <= Logical_Operator_out10559_out1;

  out320 <= Logical_Operator_out10560_out1;

  out321 <= Logical_Operator_out10561_out1;

  out322 <= Logical_Operator_out10562_out1;

  out323 <= Logical_Operator_out10563_out1;

  out324 <= Logical_Operator_out10564_out1;

  out325 <= Logical_Operator_out10565_out1;

  out326 <= Logical_Operator_out10566_out1;

  out327 <= Logical_Operator_out10567_out1;

  out328 <= Logical_Operator_out10568_out1;

  out329 <= Logical_Operator_out10569_out1;

  out330 <= Logical_Operator_out10570_out1;

  out331 <= Logical_Operator_out10571_out1;

  out332 <= Logical_Operator_out10572_out1;

  out333 <= Logical_Operator_out10573_out1;

  out334 <= Logical_Operator_out10574_out1;

  out335 <= Logical_Operator_out10575_out1;

  out336 <= Logical_Operator_out10576_out1;

  out337 <= Logical_Operator_out10577_out1;

  out338 <= Logical_Operator_out10578_out1;

  out339 <= Logical_Operator_out10579_out1;

  out340 <= Logical_Operator_out10580_out1;

  out341 <= Logical_Operator_out10581_out1;

  out342 <= Logical_Operator_out10582_out1;

  out343 <= Logical_Operator_out10583_out1;

  out344 <= Logical_Operator_out10584_out1;

  out345 <= Logical_Operator_out10585_out1;

  out346 <= Logical_Operator_out10586_out1;

  out347 <= Logical_Operator_out10587_out1;

  out348 <= Logical_Operator_out10588_out1;

  out349 <= Logical_Operator_out10589_out1;

  out350 <= Logical_Operator_out10590_out1;

  out351 <= Logical_Operator_out10591_out1;

  out352 <= Logical_Operator_out10592_out1;

  out353 <= Logical_Operator_out10593_out1;

  out354 <= Logical_Operator_out10594_out1;

  out355 <= Logical_Operator_out10595_out1;

  out356 <= Logical_Operator_out10596_out1;

  out357 <= Logical_Operator_out10597_out1;

  out358 <= Logical_Operator_out10598_out1;

  out359 <= Logical_Operator_out10599_out1;

  out360 <= Logical_Operator_out10600_out1;

  out361 <= Logical_Operator_out10601_out1;

  out362 <= Logical_Operator_out10602_out1;

  out363 <= Logical_Operator_out10603_out1;

  out364 <= Logical_Operator_out10604_out1;

  out365 <= Logical_Operator_out10605_out1;

  out366 <= Logical_Operator_out10606_out1;

  out367 <= Logical_Operator_out10607_out1;

  out368 <= Logical_Operator_out10608_out1;

  out369 <= Logical_Operator_out10609_out1;

  out370 <= Logical_Operator_out10610_out1;

  out371 <= Logical_Operator_out10611_out1;

  out372 <= Logical_Operator_out10612_out1;

  out373 <= Logical_Operator_out10613_out1;

  out374 <= Logical_Operator_out10614_out1;

  out375 <= Logical_Operator_out10615_out1;

  out376 <= Logical_Operator_out10616_out1;

  out377 <= Logical_Operator_out10617_out1;

  out378 <= Logical_Operator_out10618_out1;

  out379 <= Logical_Operator_out10619_out1;

  out380 <= Logical_Operator_out10620_out1;

  out381 <= Logical_Operator_out10621_out1;

  out382 <= Logical_Operator_out10622_out1;

  out383 <= Logical_Operator_out10623_out1;

  out384 <= Logical_Operator_out10624_out1;

  out385 <= Logical_Operator_out10625_out1;

  out386 <= Logical_Operator_out10626_out1;

  out387 <= Logical_Operator_out10627_out1;

  out388 <= Logical_Operator_out10628_out1;

  out389 <= Logical_Operator_out10629_out1;

  out390 <= Logical_Operator_out10630_out1;

  out391 <= Logical_Operator_out10631_out1;

  out392 <= Logical_Operator_out10632_out1;

  out393 <= Logical_Operator_out10633_out1;

  out394 <= Logical_Operator_out10634_out1;

  out395 <= Logical_Operator_out10635_out1;

  out396 <= Logical_Operator_out10636_out1;

  out397 <= Logical_Operator_out10637_out1;

  out398 <= Logical_Operator_out10638_out1;

  out399 <= Logical_Operator_out10639_out1;

  out400 <= Logical_Operator_out10640_out1;

  out401 <= Logical_Operator_out10641_out1;

  out402 <= Logical_Operator_out10642_out1;

  out403 <= Logical_Operator_out10643_out1;

  out404 <= Logical_Operator_out10644_out1;

  out405 <= Logical_Operator_out10645_out1;

  out406 <= Logical_Operator_out10646_out1;

  out407 <= Logical_Operator_out10647_out1;

  out408 <= Logical_Operator_out10648_out1;

  out409 <= Logical_Operator_out10649_out1;

  out410 <= Logical_Operator_out10650_out1;

  out411 <= Logical_Operator_out10651_out1;

  out412 <= Logical_Operator_out10652_out1;

  out413 <= Logical_Operator_out10653_out1;

  out414 <= Logical_Operator_out10654_out1;

  out415 <= Logical_Operator_out10655_out1;

  out416 <= Logical_Operator_out10656_out1;

  out417 <= Logical_Operator_out10657_out1;

  out418 <= Logical_Operator_out10658_out1;

  out419 <= Logical_Operator_out10659_out1;

  out420 <= Logical_Operator_out10660_out1;

  out421 <= Logical_Operator_out10661_out1;

  out422 <= Logical_Operator_out10662_out1;

  out423 <= Logical_Operator_out10663_out1;

  out424 <= Logical_Operator_out10664_out1;

  out425 <= Logical_Operator_out10665_out1;

  out426 <= Logical_Operator_out10666_out1;

  out427 <= Logical_Operator_out10667_out1;

  out428 <= Logical_Operator_out10668_out1;

  out429 <= Logical_Operator_out10669_out1;

  out430 <= Logical_Operator_out10670_out1;

  out431 <= Logical_Operator_out10671_out1;

  out432 <= Logical_Operator_out10672_out1;

  out433 <= Logical_Operator_out10673_out1;

  out434 <= Logical_Operator_out10674_out1;

  out435 <= Logical_Operator_out10675_out1;

  out436 <= Logical_Operator_out10676_out1;

  out437 <= Logical_Operator_out10677_out1;

  out438 <= Logical_Operator_out10678_out1;

  out439 <= Logical_Operator_out10679_out1;

  out440 <= Logical_Operator_out10680_out1;

  out441 <= Logical_Operator_out10681_out1;

  out442 <= Logical_Operator_out10682_out1;

  out443 <= Logical_Operator_out10683_out1;

  out444 <= Logical_Operator_out10684_out1;

  out445 <= Logical_Operator_out10685_out1;

  out446 <= Logical_Operator_out10686_out1;

  out447 <= Logical_Operator_out10687_out1;

  out448 <= Logical_Operator_out10688_out1;

  out449 <= Logical_Operator_out10689_out1;

  out450 <= Logical_Operator_out10690_out1;

  out451 <= Logical_Operator_out10691_out1;

  out452 <= Logical_Operator_out10692_out1;

  out453 <= Logical_Operator_out10693_out1;

  out454 <= Logical_Operator_out10694_out1;

  out455 <= Logical_Operator_out10695_out1;

  out456 <= Logical_Operator_out10696_out1;

  out457 <= Logical_Operator_out10697_out1;

  out458 <= Logical_Operator_out10698_out1;

  out459 <= Logical_Operator_out10699_out1;

  out460 <= Logical_Operator_out10700_out1;

  out461 <= Logical_Operator_out10701_out1;

  out462 <= Logical_Operator_out10702_out1;

  out463 <= Logical_Operator_out10703_out1;

  out464 <= Logical_Operator_out10704_out1;

  out465 <= Logical_Operator_out10705_out1;

  out466 <= Logical_Operator_out10706_out1;

  out467 <= Logical_Operator_out10707_out1;

  out468 <= Logical_Operator_out10708_out1;

  out469 <= Logical_Operator_out10709_out1;

  out470 <= Logical_Operator_out10710_out1;

  out471 <= Logical_Operator_out10711_out1;

  out472 <= Logical_Operator_out10712_out1;

  out473 <= Logical_Operator_out10713_out1;

  out474 <= Logical_Operator_out10714_out1;

  out475 <= Logical_Operator_out10715_out1;

  out476 <= Logical_Operator_out10716_out1;

  out477 <= Logical_Operator_out10717_out1;

  out478 <= Logical_Operator_out10718_out1;

  out479 <= Logical_Operator_out10719_out1;

  out480 <= Logical_Operator_out10720_out1;

  out481 <= Logical_Operator_out10721_out1;

  out482 <= Logical_Operator_out10722_out1;

  out483 <= Logical_Operator_out10723_out1;

  out484 <= Logical_Operator_out10724_out1;

  out485 <= Logical_Operator_out10725_out1;

  out486 <= Logical_Operator_out10726_out1;

  out487 <= Logical_Operator_out10727_out1;

  out488 <= Logical_Operator_out10728_out1;

  out489 <= Logical_Operator_out10729_out1;

  out490 <= Logical_Operator_out10730_out1;

  out491 <= Logical_Operator_out10731_out1;

  out492 <= Logical_Operator_out10732_out1;

  out493 <= Logical_Operator_out10733_out1;

  out494 <= Logical_Operator_out10734_out1;

  out495 <= Logical_Operator_out10735_out1;

  out496 <= Logical_Operator_out10736_out1;

  out497 <= Logical_Operator_out10737_out1;

  out498 <= Logical_Operator_out10738_out1;

  out499 <= Logical_Operator_out10739_out1;

  out500 <= Logical_Operator_out10740_out1;

  out501 <= Logical_Operator_out10741_out1;

  out502 <= Logical_Operator_out10742_out1;

  out503 <= Logical_Operator_out10743_out1;

  out504 <= Logical_Operator_out10744_out1;

  out505 <= Logical_Operator_out10745_out1;

  out506 <= Logical_Operator_out10746_out1;

  out507 <= Logical_Operator_out10747_out1;

  out508 <= Logical_Operator_out10748_out1;

  out509 <= Logical_Operator_out10749_out1;

  out510 <= Logical_Operator_out10750_out1;

  out511 <= Logical_Operator_out10751_out1;

  out512 <= Logical_Operator_out10752_out1;

  out513 <= Logical_Operator_out10753_out1;

  out514 <= Logical_Operator_out10754_out1;

  out515 <= Logical_Operator_out10755_out1;

  out516 <= Logical_Operator_out10756_out1;

  out517 <= Logical_Operator_out10757_out1;

  out518 <= Logical_Operator_out10758_out1;

  out519 <= Logical_Operator_out10759_out1;

  out520 <= Logical_Operator_out10760_out1;

  out521 <= Logical_Operator_out10761_out1;

  out522 <= Logical_Operator_out10762_out1;

  out523 <= Logical_Operator_out10763_out1;

  out524 <= Logical_Operator_out10764_out1;

  out525 <= Logical_Operator_out10765_out1;

  out526 <= Logical_Operator_out10766_out1;

  out527 <= Logical_Operator_out10767_out1;

  out528 <= Logical_Operator_out10768_out1;

  out529 <= Logical_Operator_out10769_out1;

  out530 <= Logical_Operator_out10770_out1;

  out531 <= Logical_Operator_out10771_out1;

  out532 <= Logical_Operator_out10772_out1;

  out533 <= Logical_Operator_out10773_out1;

  out534 <= Logical_Operator_out10774_out1;

  out535 <= Logical_Operator_out10775_out1;

  out536 <= Logical_Operator_out10776_out1;

  out537 <= Logical_Operator_out10777_out1;

  out538 <= Logical_Operator_out10778_out1;

  out539 <= Logical_Operator_out10779_out1;

  out540 <= Logical_Operator_out10780_out1;

  out541 <= Logical_Operator_out10781_out1;

  out542 <= Logical_Operator_out10782_out1;

  out543 <= Logical_Operator_out10783_out1;

  out544 <= Logical_Operator_out10784_out1;

  out545 <= Logical_Operator_out10785_out1;

  out546 <= Logical_Operator_out10786_out1;

  out547 <= Logical_Operator_out10787_out1;

  out548 <= Logical_Operator_out10788_out1;

  out549 <= Logical_Operator_out10789_out1;

  out550 <= Logical_Operator_out10790_out1;

  out551 <= Logical_Operator_out10791_out1;

  out552 <= Logical_Operator_out10792_out1;

  out553 <= Logical_Operator_out10793_out1;

  out554 <= Logical_Operator_out10794_out1;

  out555 <= Logical_Operator_out10795_out1;

  out556 <= Logical_Operator_out10796_out1;

  out557 <= Logical_Operator_out10797_out1;

  out558 <= Logical_Operator_out10798_out1;

  out559 <= Logical_Operator_out10799_out1;

  out560 <= Logical_Operator_out10800_out1;

  out561 <= Logical_Operator_out10801_out1;

  out562 <= Logical_Operator_out10802_out1;

  out563 <= Logical_Operator_out10803_out1;

  out564 <= Logical_Operator_out10804_out1;

  out565 <= Logical_Operator_out10805_out1;

  out566 <= Logical_Operator_out10806_out1;

  out567 <= Logical_Operator_out10807_out1;

  out568 <= Logical_Operator_out10808_out1;

  out569 <= Logical_Operator_out10809_out1;

  out570 <= Logical_Operator_out10810_out1;

  out571 <= Logical_Operator_out10811_out1;

  out572 <= Logical_Operator_out10812_out1;

  out573 <= Logical_Operator_out10813_out1;

  out574 <= Logical_Operator_out10814_out1;

  out575 <= Logical_Operator_out10815_out1;

  out576 <= Logical_Operator_out10816_out1;

  out577 <= Logical_Operator_out10817_out1;

  out578 <= Logical_Operator_out10818_out1;

  out579 <= Logical_Operator_out10819_out1;

  out580 <= Logical_Operator_out10820_out1;

  out581 <= Logical_Operator_out10821_out1;

  out582 <= Logical_Operator_out10822_out1;

  out583 <= Logical_Operator_out10823_out1;

  out584 <= Logical_Operator_out10824_out1;

  out585 <= Logical_Operator_out10825_out1;

  out586 <= Logical_Operator_out10826_out1;

  out587 <= Logical_Operator_out10827_out1;

  out588 <= Logical_Operator_out10828_out1;

  out589 <= Logical_Operator_out10829_out1;

  out590 <= Logical_Operator_out10830_out1;

  out591 <= Logical_Operator_out10831_out1;

  out592 <= Logical_Operator_out10832_out1;

  out593 <= Logical_Operator_out10833_out1;

  out594 <= Logical_Operator_out10834_out1;

  out595 <= Logical_Operator_out10835_out1;

  out596 <= Logical_Operator_out10836_out1;

  out597 <= Logical_Operator_out10837_out1;

  out598 <= Logical_Operator_out10838_out1;

  out599 <= Logical_Operator_out10839_out1;

  out600 <= Logical_Operator_out10840_out1;

  out601 <= Logical_Operator_out10841_out1;

  out602 <= Logical_Operator_out10842_out1;

  out603 <= Logical_Operator_out10843_out1;

  out604 <= Logical_Operator_out10844_out1;

  out605 <= Logical_Operator_out10845_out1;

  out606 <= Logical_Operator_out10846_out1;

  out607 <= Logical_Operator_out10847_out1;

  out608 <= Logical_Operator_out10848_out1;

  out609 <= Logical_Operator_out10849_out1;

  out610 <= Logical_Operator_out10850_out1;

  out611 <= Logical_Operator_out10851_out1;

  out612 <= Logical_Operator_out10852_out1;

  out613 <= Logical_Operator_out10853_out1;

  out614 <= Logical_Operator_out10854_out1;

  out615 <= Logical_Operator_out10855_out1;

  out616 <= Logical_Operator_out10856_out1;

  out617 <= Logical_Operator_out10857_out1;

  out618 <= Logical_Operator_out10858_out1;

  out619 <= Logical_Operator_out10859_out1;

  out620 <= Logical_Operator_out10860_out1;

  out621 <= Logical_Operator_out10861_out1;

  out622 <= Logical_Operator_out10862_out1;

  out623 <= Logical_Operator_out10863_out1;

  out624 <= Logical_Operator_out10864_out1;

  out625 <= Logical_Operator_out10865_out1;

  out626 <= Logical_Operator_out10866_out1;

  out627 <= Logical_Operator_out10867_out1;

  out628 <= Logical_Operator_out10868_out1;

  out629 <= Logical_Operator_out10869_out1;

  out630 <= Logical_Operator_out10870_out1;

  out631 <= Logical_Operator_out10871_out1;

  out632 <= Logical_Operator_out10872_out1;

  out633 <= Logical_Operator_out10873_out1;

  out634 <= Logical_Operator_out10874_out1;

  out635 <= Logical_Operator_out10875_out1;

  out636 <= Logical_Operator_out10876_out1;

  out637 <= Logical_Operator_out10877_out1;

  out638 <= Logical_Operator_out10878_out1;

  out639 <= Logical_Operator_out10879_out1;

  out640 <= Logical_Operator_out10880_out1;

  out641 <= Logical_Operator_out10881_out1;

  out642 <= Logical_Operator_out10882_out1;

  out643 <= Logical_Operator_out10883_out1;

  out644 <= Logical_Operator_out10884_out1;

  out645 <= Logical_Operator_out10885_out1;

  out646 <= Logical_Operator_out10886_out1;

  out647 <= Logical_Operator_out10887_out1;

  out648 <= Logical_Operator_out10888_out1;

  out649 <= Logical_Operator_out10889_out1;

  out650 <= Logical_Operator_out10890_out1;

  out651 <= Logical_Operator_out10891_out1;

  out652 <= Logical_Operator_out10892_out1;

  out653 <= Logical_Operator_out10893_out1;

  out654 <= Logical_Operator_out10894_out1;

  out655 <= Logical_Operator_out10895_out1;

  out656 <= Logical_Operator_out10896_out1;

  out657 <= Logical_Operator_out10897_out1;

  out658 <= Logical_Operator_out10898_out1;

  out659 <= Logical_Operator_out10899_out1;

  out660 <= Logical_Operator_out10900_out1;

  out661 <= Logical_Operator_out10901_out1;

  out662 <= Logical_Operator_out10902_out1;

  out663 <= Logical_Operator_out10903_out1;

  out664 <= Logical_Operator_out10904_out1;

  out665 <= Logical_Operator_out10905_out1;

  out666 <= Logical_Operator_out10906_out1;

  out667 <= Logical_Operator_out10907_out1;

  out668 <= Logical_Operator_out10908_out1;

  out669 <= Logical_Operator_out10909_out1;

  out670 <= Logical_Operator_out10910_out1;

  out671 <= Logical_Operator_out10911_out1;

  out672 <= Logical_Operator_out10912_out1;

  out673 <= Logical_Operator_out10913_out1;

  out674 <= Logical_Operator_out10914_out1;

  out675 <= Logical_Operator_out10915_out1;

  out676 <= Logical_Operator_out10916_out1;

  out677 <= Logical_Operator_out10917_out1;

  out678 <= Logical_Operator_out10918_out1;

  out679 <= Logical_Operator_out10919_out1;

  out680 <= Logical_Operator_out10920_out1;

  out681 <= Logical_Operator_out10921_out1;

  out682 <= Logical_Operator_out10922_out1;

  out683 <= Logical_Operator_out10923_out1;

  out684 <= Logical_Operator_out10924_out1;

  out685 <= Logical_Operator_out10925_out1;

  out686 <= Logical_Operator_out10926_out1;

  out687 <= Logical_Operator_out10927_out1;

  out688 <= Logical_Operator_out10928_out1;

  out689 <= Logical_Operator_out10929_out1;

  out690 <= Logical_Operator_out10930_out1;

  out691 <= Logical_Operator_out10931_out1;

  out692 <= Logical_Operator_out10932_out1;

  out693 <= Logical_Operator_out10933_out1;

  out694 <= Logical_Operator_out10934_out1;

  out695 <= Logical_Operator_out10935_out1;

  out696 <= Logical_Operator_out10936_out1;

  out697 <= Logical_Operator_out10937_out1;

  out698 <= Logical_Operator_out10938_out1;

  out699 <= Logical_Operator_out10939_out1;

  out700 <= Logical_Operator_out10940_out1;

  out701 <= Logical_Operator_out10941_out1;

  out702 <= Logical_Operator_out10942_out1;

  out703 <= Logical_Operator_out10943_out1;

  out704 <= Logical_Operator_out10944_out1;

  out705 <= Logical_Operator_out10945_out1;

  out706 <= Logical_Operator_out10946_out1;

  out707 <= Logical_Operator_out10947_out1;

  out708 <= Logical_Operator_out10948_out1;

  out709 <= Logical_Operator_out10949_out1;

  out710 <= Logical_Operator_out10950_out1;

  out711 <= Logical_Operator_out10951_out1;

  out712 <= Logical_Operator_out10952_out1;

  out713 <= Logical_Operator_out10953_out1;

  out714 <= Logical_Operator_out10954_out1;

  out715 <= Logical_Operator_out10955_out1;

  out716 <= Logical_Operator_out10956_out1;

  out717 <= Logical_Operator_out10957_out1;

  out718 <= Logical_Operator_out10958_out1;

  out719 <= Logical_Operator_out10959_out1;

  out720 <= Logical_Operator_out10960_out1;

  out721 <= Logical_Operator_out10961_out1;

  out722 <= Logical_Operator_out10962_out1;

  out723 <= Logical_Operator_out10963_out1;

  out724 <= Logical_Operator_out10964_out1;

  out725 <= Logical_Operator_out10965_out1;

  out726 <= Logical_Operator_out10966_out1;

  out727 <= Logical_Operator_out10967_out1;

  out728 <= Logical_Operator_out10968_out1;

  out729 <= Logical_Operator_out10969_out1;

  out730 <= Logical_Operator_out10970_out1;

  out731 <= Logical_Operator_out10971_out1;

  out732 <= Logical_Operator_out10972_out1;

  out733 <= Logical_Operator_out10973_out1;

  out734 <= Logical_Operator_out10974_out1;

  out735 <= Logical_Operator_out10975_out1;

  out736 <= Logical_Operator_out10976_out1;

  out737 <= Logical_Operator_out10977_out1;

  out738 <= Logical_Operator_out10978_out1;

  out739 <= Logical_Operator_out10979_out1;

  out740 <= Logical_Operator_out10980_out1;

  out741 <= Logical_Operator_out10981_out1;

  out742 <= Logical_Operator_out10982_out1;

  out743 <= Logical_Operator_out10983_out1;

  out744 <= Logical_Operator_out10984_out1;

  out745 <= Logical_Operator_out10985_out1;

  out746 <= Logical_Operator_out10986_out1;

  out747 <= Logical_Operator_out10987_out1;

  out748 <= Logical_Operator_out10988_out1;

  out749 <= Logical_Operator_out10989_out1;

  out750 <= Logical_Operator_out10990_out1;

  out751 <= Logical_Operator_out10991_out1;

  out752 <= Logical_Operator_out10992_out1;

  out753 <= Logical_Operator_out10993_out1;

  out754 <= Logical_Operator_out10994_out1;

  out755 <= Logical_Operator_out10995_out1;

  out756 <= Logical_Operator_out10996_out1;

  out757 <= Logical_Operator_out10997_out1;

  out758 <= Logical_Operator_out10998_out1;

  out759 <= Logical_Operator_out10999_out1;

  out760 <= Logical_Operator_out11000_out1;

  out761 <= Logical_Operator_out11001_out1;

  out762 <= Logical_Operator_out11002_out1;

  out763 <= Logical_Operator_out11003_out1;

  out764 <= Logical_Operator_out11004_out1;

  out765 <= Logical_Operator_out11005_out1;

  out766 <= Logical_Operator_out11006_out1;

  out767 <= Logical_Operator_out11007_out1;

  out768 <= Logical_Operator_out11008_out1;

  out769 <= Logical_Operator_out11009_out1;

  out770 <= Logical_Operator_out11010_out1;

  out771 <= Logical_Operator_out11011_out1;

  out772 <= Logical_Operator_out11012_out1;

  out773 <= Logical_Operator_out11013_out1;

  out774 <= Logical_Operator_out11014_out1;

  out775 <= Logical_Operator_out11015_out1;

  out776 <= Logical_Operator_out11016_out1;

  out777 <= Logical_Operator_out11017_out1;

  out778 <= Logical_Operator_out11018_out1;

  out779 <= Logical_Operator_out11019_out1;

  out780 <= Logical_Operator_out11020_out1;

  out781 <= Logical_Operator_out11021_out1;

  out782 <= Logical_Operator_out11022_out1;

  out783 <= Logical_Operator_out11023_out1;

  out784 <= Logical_Operator_out11024_out1;

  out785 <= Logical_Operator_out11025_out1;

  out786 <= Logical_Operator_out11026_out1;

  out787 <= Logical_Operator_out11027_out1;

  out788 <= Logical_Operator_out11028_out1;

  out789 <= Logical_Operator_out11029_out1;

  out790 <= Logical_Operator_out11030_out1;

  out791 <= Logical_Operator_out11031_out1;

  out792 <= Logical_Operator_out11032_out1;

  out793 <= Logical_Operator_out11033_out1;

  out794 <= Logical_Operator_out11034_out1;

  out795 <= Logical_Operator_out11035_out1;

  out796 <= Logical_Operator_out11036_out1;

  out797 <= Logical_Operator_out11037_out1;

  out798 <= Logical_Operator_out11038_out1;

  out799 <= Logical_Operator_out11039_out1;

  out800 <= Logical_Operator_out11040_out1;

  out801 <= Logical_Operator_out11041_out1;

  out802 <= Logical_Operator_out11042_out1;

  out803 <= Logical_Operator_out11043_out1;

  out804 <= Logical_Operator_out11044_out1;

  out805 <= Logical_Operator_out11045_out1;

  out806 <= Logical_Operator_out11046_out1;

  out807 <= Logical_Operator_out11047_out1;

  out808 <= Logical_Operator_out11048_out1;

  out809 <= Logical_Operator_out11049_out1;

  out810 <= Logical_Operator_out11050_out1;

  out811 <= Logical_Operator_out11051_out1;

  out812 <= Logical_Operator_out11052_out1;

  out813 <= Logical_Operator_out11053_out1;

  out814 <= Logical_Operator_out11054_out1;

  out815 <= Logical_Operator_out11055_out1;

  out816 <= Logical_Operator_out11056_out1;

  out817 <= Logical_Operator_out11057_out1;

  out818 <= Logical_Operator_out11058_out1;

  out819 <= Logical_Operator_out11059_out1;

  out820 <= Logical_Operator_out11060_out1;

  out821 <= Logical_Operator_out11061_out1;

  out822 <= Logical_Operator_out11062_out1;

  out823 <= Logical_Operator_out11063_out1;

  out824 <= Logical_Operator_out11064_out1;

  out825 <= Logical_Operator_out11065_out1;

  out826 <= Logical_Operator_out11066_out1;

  out827 <= Logical_Operator_out11067_out1;

  out828 <= Logical_Operator_out11068_out1;

  out829 <= Logical_Operator_out11069_out1;

  out830 <= Logical_Operator_out11070_out1;

  out831 <= Logical_Operator_out11071_out1;

  out832 <= Logical_Operator_out11072_out1;

  out833 <= Logical_Operator_out11073_out1;

  out834 <= Logical_Operator_out11074_out1;

  out835 <= Logical_Operator_out11075_out1;

  out836 <= Logical_Operator_out11076_out1;

  out837 <= Logical_Operator_out11077_out1;

  out838 <= Logical_Operator_out11078_out1;

  out839 <= Logical_Operator_out11079_out1;

  out840 <= Logical_Operator_out11080_out1;

  out841 <= Logical_Operator_out11081_out1;

  out842 <= Logical_Operator_out11082_out1;

  out843 <= Logical_Operator_out11083_out1;

  out844 <= Logical_Operator_out11084_out1;

  out845 <= Logical_Operator_out11085_out1;

  out846 <= Logical_Operator_out11086_out1;

  out847 <= Logical_Operator_out11087_out1;

  out848 <= Logical_Operator_out11088_out1;

  out849 <= Logical_Operator_out11089_out1;

  out850 <= Logical_Operator_out11090_out1;

  out851 <= Logical_Operator_out11091_out1;

  out852 <= Logical_Operator_out11092_out1;

  out853 <= Logical_Operator_out11093_out1;

  out854 <= Logical_Operator_out11094_out1;

  out855 <= Logical_Operator_out11095_out1;

  out856 <= Logical_Operator_out11096_out1;

  out857 <= Logical_Operator_out11097_out1;

  out858 <= Logical_Operator_out11098_out1;

  out859 <= Logical_Operator_out11099_out1;

  out860 <= Logical_Operator_out11100_out1;

  out861 <= Logical_Operator_out11101_out1;

  out862 <= Logical_Operator_out11102_out1;

  out863 <= Logical_Operator_out11103_out1;

  out864 <= Logical_Operator_out11104_out1;

  out865 <= Logical_Operator_out11105_out1;

  out866 <= Logical_Operator_out11106_out1;

  out867 <= Logical_Operator_out11107_out1;

  out868 <= Logical_Operator_out11108_out1;

  out869 <= Logical_Operator_out11109_out1;

  out870 <= Logical_Operator_out11110_out1;

  out871 <= Logical_Operator_out11111_out1;

  out872 <= Logical_Operator_out11112_out1;

  out873 <= Logical_Operator_out11113_out1;

  out874 <= Logical_Operator_out11114_out1;

  out875 <= Logical_Operator_out11115_out1;

  out876 <= Logical_Operator_out11116_out1;

  out877 <= Logical_Operator_out11117_out1;

  out878 <= Logical_Operator_out11118_out1;

  out879 <= Logical_Operator_out11119_out1;

  out880 <= Logical_Operator_out11120_out1;

  out881 <= Logical_Operator_out11121_out1;

  out882 <= Logical_Operator_out11122_out1;

  out883 <= Logical_Operator_out11123_out1;

  out884 <= Logical_Operator_out11124_out1;

  out885 <= Logical_Operator_out11125_out1;

  out886 <= Logical_Operator_out11126_out1;

  out887 <= Logical_Operator_out11127_out1;

  out888 <= Logical_Operator_out11128_out1;

  out889 <= Logical_Operator_out11129_out1;

  out890 <= Logical_Operator_out11130_out1;

  out891 <= Logical_Operator_out11131_out1;

  out892 <= Logical_Operator_out11132_out1;

  out893 <= Logical_Operator_out11133_out1;

  out894 <= Logical_Operator_out11134_out1;

  out895 <= Logical_Operator_out11135_out1;

  out896 <= Logical_Operator_out11136_out1;

  out897 <= Logical_Operator_out11137_out1;

  out898 <= Logical_Operator_out11138_out1;

  out899 <= Logical_Operator_out11139_out1;

  out900 <= Logical_Operator_out11140_out1;

  out901 <= Logical_Operator_out11141_out1;

  out902 <= Logical_Operator_out11142_out1;

  out903 <= Logical_Operator_out11143_out1;

  out904 <= Logical_Operator_out11144_out1;

  out905 <= Logical_Operator_out11145_out1;

  out906 <= Logical_Operator_out11146_out1;

  out907 <= Logical_Operator_out11147_out1;

  out908 <= Logical_Operator_out11148_out1;

  out909 <= Logical_Operator_out11149_out1;

  out910 <= Logical_Operator_out11150_out1;

  out911 <= Logical_Operator_out11151_out1;

  out912 <= Logical_Operator_out11152_out1;

  out913 <= Logical_Operator_out11153_out1;

  out914 <= Logical_Operator_out11154_out1;

  out915 <= Logical_Operator_out11155_out1;

  out916 <= Logical_Operator_out11156_out1;

  out917 <= Logical_Operator_out11157_out1;

  out918 <= Logical_Operator_out11158_out1;

  out919 <= Logical_Operator_out11159_out1;

  out920 <= Logical_Operator_out11160_out1;

  out921 <= Logical_Operator_out11161_out1;

  out922 <= Logical_Operator_out11162_out1;

  out923 <= Logical_Operator_out11163_out1;

  out924 <= Logical_Operator_out11164_out1;

  out925 <= Logical_Operator_out11165_out1;

  out926 <= Logical_Operator_out11166_out1;

  out927 <= Logical_Operator_out11167_out1;

  out928 <= Logical_Operator_out11168_out1;

  out929 <= Logical_Operator_out11169_out1;

  out930 <= Logical_Operator_out11170_out1;

  out931 <= Logical_Operator_out11171_out1;

  out932 <= Logical_Operator_out11172_out1;

  out933 <= Logical_Operator_out11173_out1;

  out934 <= Logical_Operator_out11174_out1;

  out935 <= Logical_Operator_out11175_out1;

  out936 <= Logical_Operator_out11176_out1;

  out937 <= Logical_Operator_out11177_out1;

  out938 <= Logical_Operator_out11178_out1;

  out939 <= Logical_Operator_out11179_out1;

  out940 <= Logical_Operator_out11180_out1;

  out941 <= Logical_Operator_out11181_out1;

  out942 <= Logical_Operator_out11182_out1;

  out943 <= Logical_Operator_out11183_out1;

  out944 <= Logical_Operator_out11184_out1;

  out945 <= Logical_Operator_out11185_out1;

  out946 <= Logical_Operator_out11186_out1;

  out947 <= Logical_Operator_out11187_out1;

  out948 <= Logical_Operator_out11188_out1;

  out949 <= Logical_Operator_out11189_out1;

  out950 <= Logical_Operator_out11190_out1;

  out951 <= Logical_Operator_out11191_out1;

  out952 <= Logical_Operator_out11192_out1;

  out953 <= Logical_Operator_out11193_out1;

  out954 <= Logical_Operator_out11194_out1;

  out955 <= Logical_Operator_out11195_out1;

  out956 <= Logical_Operator_out11196_out1;

  out957 <= Logical_Operator_out11197_out1;

  out958 <= Logical_Operator_out11198_out1;

  out959 <= Logical_Operator_out11199_out1;

  out960 <= Logical_Operator_out11200_out1;

  out961 <= Logical_Operator_out11201_out1;

  out962 <= Logical_Operator_out11202_out1;

  out963 <= Logical_Operator_out11203_out1;

  out964 <= Logical_Operator_out11204_out1;

  out965 <= Logical_Operator_out11205_out1;

  out966 <= Logical_Operator_out11206_out1;

  out967 <= Logical_Operator_out11207_out1;

  out968 <= Logical_Operator_out11208_out1;

  out969 <= Logical_Operator_out11209_out1;

  out970 <= Logical_Operator_out11210_out1;

  out971 <= Logical_Operator_out11211_out1;

  out972 <= Logical_Operator_out11212_out1;

  out973 <= Logical_Operator_out11213_out1;

  out974 <= Logical_Operator_out11214_out1;

  out975 <= Logical_Operator_out11215_out1;

  out976 <= Logical_Operator_out11216_out1;

  out977 <= Logical_Operator_out11217_out1;

  out978 <= Logical_Operator_out11218_out1;

  out979 <= Logical_Operator_out11219_out1;

  out980 <= Logical_Operator_out11220_out1;

  out981 <= Logical_Operator_out11221_out1;

  out982 <= Logical_Operator_out11222_out1;

  out983 <= Logical_Operator_out11223_out1;

  out984 <= Logical_Operator_out11224_out1;

  out985 <= Logical_Operator_out11225_out1;

  out986 <= Logical_Operator_out11226_out1;

  out987 <= Logical_Operator_out11227_out1;

  out988 <= Logical_Operator_out11228_out1;

  out989 <= Logical_Operator_out11229_out1;

  out990 <= Logical_Operator_out11230_out1;

  out991 <= Logical_Operator_out11231_out1;

  out992 <= Logical_Operator_out11232_out1;

  out993 <= Logical_Operator_out11233_out1;

  out994 <= Logical_Operator_out11234_out1;

  out995 <= Logical_Operator_out11235_out1;

  out996 <= Logical_Operator_out11236_out1;

  out997 <= Logical_Operator_out11237_out1;

  out998 <= Logical_Operator_out11238_out1;

  out999 <= Logical_Operator_out11239_out1;

  out1000 <= Logical_Operator_out11240_out1;

  out1001 <= Logical_Operator_out11241_out1;

  out1002 <= Logical_Operator_out11242_out1;

  out1003 <= Logical_Operator_out11243_out1;

  out1004 <= Logical_Operator_out11244_out1;

  out1005 <= Logical_Operator_out11245_out1;

  out1006 <= Logical_Operator_out11246_out1;

  out1007 <= Logical_Operator_out11247_out1;

  out1008 <= Logical_Operator_out11248_out1;

  out1009 <= Logical_Operator_out11249_out1;

  out1010 <= Logical_Operator_out11250_out1;

  out1011 <= Logical_Operator_out11251_out1;

  out1012 <= Logical_Operator_out11252_out1;

  out1013 <= Logical_Operator_out11253_out1;

  out1014 <= Logical_Operator_out11254_out1;

  out1015 <= Logical_Operator_out11255_out1;

  out1016 <= Logical_Operator_out11256_out1;

  out1017 <= Logical_Operator_out11257_out1;

  out1018 <= Logical_Operator_out11258_out1;

  out1019 <= Logical_Operator_out11259_out1;

  out1020 <= Logical_Operator_out11260_out1;

  out1021 <= Logical_Operator_out11261_out1;

  out1022 <= Logical_Operator_out11262_out1;

  out1023 <= Logical_Operator_out11263_out1;

  out1024 <= Logical_Operator_out11264_out1;

  out1025 <= Logical_Operator_out9729_out1;

  out1026 <= Logical_Operator_out9730_out1;

  out1027 <= Logical_Operator_out9731_out1;

  out1028 <= Logical_Operator_out9732_out1;

  out1029 <= Logical_Operator_out9733_out1;

  out1030 <= Logical_Operator_out9734_out1;

  out1031 <= Logical_Operator_out9735_out1;

  out1032 <= Logical_Operator_out9736_out1;

  out1033 <= Logical_Operator_out9737_out1;

  out1034 <= Logical_Operator_out9738_out1;

  out1035 <= Logical_Operator_out9739_out1;

  out1036 <= Logical_Operator_out9740_out1;

  out1037 <= Logical_Operator_out9741_out1;

  out1038 <= Logical_Operator_out9742_out1;

  out1039 <= Logical_Operator_out9743_out1;

  out1040 <= Logical_Operator_out9744_out1;

  out1041 <= Logical_Operator_out9745_out1;

  out1042 <= Logical_Operator_out9746_out1;

  out1043 <= Logical_Operator_out9747_out1;

  out1044 <= Logical_Operator_out9748_out1;

  out1045 <= Logical_Operator_out9749_out1;

  out1046 <= Logical_Operator_out9750_out1;

  out1047 <= Logical_Operator_out9751_out1;

  out1048 <= Logical_Operator_out9752_out1;

  out1049 <= Logical_Operator_out9753_out1;

  out1050 <= Logical_Operator_out9754_out1;

  out1051 <= Logical_Operator_out9755_out1;

  out1052 <= Logical_Operator_out9756_out1;

  out1053 <= Logical_Operator_out9757_out1;

  out1054 <= Logical_Operator_out9758_out1;

  out1055 <= Logical_Operator_out9759_out1;

  out1056 <= Logical_Operator_out9760_out1;

  out1057 <= Logical_Operator_out9761_out1;

  out1058 <= Logical_Operator_out9762_out1;

  out1059 <= Logical_Operator_out9763_out1;

  out1060 <= Logical_Operator_out9764_out1;

  out1061 <= Logical_Operator_out9765_out1;

  out1062 <= Logical_Operator_out9766_out1;

  out1063 <= Logical_Operator_out9767_out1;

  out1064 <= Logical_Operator_out9768_out1;

  out1065 <= Logical_Operator_out9769_out1;

  out1066 <= Logical_Operator_out9770_out1;

  out1067 <= Logical_Operator_out9771_out1;

  out1068 <= Logical_Operator_out9772_out1;

  out1069 <= Logical_Operator_out9773_out1;

  out1070 <= Logical_Operator_out9774_out1;

  out1071 <= Logical_Operator_out9775_out1;

  out1072 <= Logical_Operator_out9776_out1;

  out1073 <= Logical_Operator_out9777_out1;

  out1074 <= Logical_Operator_out9778_out1;

  out1075 <= Logical_Operator_out9779_out1;

  out1076 <= Logical_Operator_out9780_out1;

  out1077 <= Logical_Operator_out9781_out1;

  out1078 <= Logical_Operator_out9782_out1;

  out1079 <= Logical_Operator_out9783_out1;

  out1080 <= Logical_Operator_out9784_out1;

  out1081 <= Logical_Operator_out9785_out1;

  out1082 <= Logical_Operator_out9786_out1;

  out1083 <= Logical_Operator_out9787_out1;

  out1084 <= Logical_Operator_out9788_out1;

  out1085 <= Logical_Operator_out9789_out1;

  out1086 <= Logical_Operator_out9790_out1;

  out1087 <= Logical_Operator_out9791_out1;

  out1088 <= Logical_Operator_out9792_out1;

  out1089 <= Logical_Operator_out9793_out1;

  out1090 <= Logical_Operator_out9794_out1;

  out1091 <= Logical_Operator_out9795_out1;

  out1092 <= Logical_Operator_out9796_out1;

  out1093 <= Logical_Operator_out9797_out1;

  out1094 <= Logical_Operator_out9798_out1;

  out1095 <= Logical_Operator_out9799_out1;

  out1096 <= Logical_Operator_out9800_out1;

  out1097 <= Logical_Operator_out9801_out1;

  out1098 <= Logical_Operator_out9802_out1;

  out1099 <= Logical_Operator_out9803_out1;

  out1100 <= Logical_Operator_out9804_out1;

  out1101 <= Logical_Operator_out9805_out1;

  out1102 <= Logical_Operator_out9806_out1;

  out1103 <= Logical_Operator_out9807_out1;

  out1104 <= Logical_Operator_out9808_out1;

  out1105 <= Logical_Operator_out9809_out1;

  out1106 <= Logical_Operator_out9810_out1;

  out1107 <= Logical_Operator_out9811_out1;

  out1108 <= Logical_Operator_out9812_out1;

  out1109 <= Logical_Operator_out9813_out1;

  out1110 <= Logical_Operator_out9814_out1;

  out1111 <= Logical_Operator_out9815_out1;

  out1112 <= Logical_Operator_out9816_out1;

  out1113 <= Logical_Operator_out9817_out1;

  out1114 <= Logical_Operator_out9818_out1;

  out1115 <= Logical_Operator_out9819_out1;

  out1116 <= Logical_Operator_out9820_out1;

  out1117 <= Logical_Operator_out9821_out1;

  out1118 <= Logical_Operator_out9822_out1;

  out1119 <= Logical_Operator_out9823_out1;

  out1120 <= Logical_Operator_out9824_out1;

  out1121 <= Logical_Operator_out9825_out1;

  out1122 <= Logical_Operator_out9826_out1;

  out1123 <= Logical_Operator_out9827_out1;

  out1124 <= Logical_Operator_out9828_out1;

  out1125 <= Logical_Operator_out9829_out1;

  out1126 <= Logical_Operator_out9830_out1;

  out1127 <= Logical_Operator_out9831_out1;

  out1128 <= Logical_Operator_out9832_out1;

  out1129 <= Logical_Operator_out9833_out1;

  out1130 <= Logical_Operator_out9834_out1;

  out1131 <= Logical_Operator_out9835_out1;

  out1132 <= Logical_Operator_out9836_out1;

  out1133 <= Logical_Operator_out9837_out1;

  out1134 <= Logical_Operator_out9838_out1;

  out1135 <= Logical_Operator_out9839_out1;

  out1136 <= Logical_Operator_out9840_out1;

  out1137 <= Logical_Operator_out9841_out1;

  out1138 <= Logical_Operator_out9842_out1;

  out1139 <= Logical_Operator_out9843_out1;

  out1140 <= Logical_Operator_out9844_out1;

  out1141 <= Logical_Operator_out9845_out1;

  out1142 <= Logical_Operator_out9846_out1;

  out1143 <= Logical_Operator_out9847_out1;

  out1144 <= Logical_Operator_out9848_out1;

  out1145 <= Logical_Operator_out9849_out1;

  out1146 <= Logical_Operator_out9850_out1;

  out1147 <= Logical_Operator_out9851_out1;

  out1148 <= Logical_Operator_out9852_out1;

  out1149 <= Logical_Operator_out9853_out1;

  out1150 <= Logical_Operator_out9854_out1;

  out1151 <= Logical_Operator_out9855_out1;

  out1152 <= Logical_Operator_out9856_out1;

  out1153 <= Logical_Operator_out9857_out1;

  out1154 <= Logical_Operator_out9858_out1;

  out1155 <= Logical_Operator_out9859_out1;

  out1156 <= Logical_Operator_out9860_out1;

  out1157 <= Logical_Operator_out9861_out1;

  out1158 <= Logical_Operator_out9862_out1;

  out1159 <= Logical_Operator_out9863_out1;

  out1160 <= Logical_Operator_out9864_out1;

  out1161 <= Logical_Operator_out9865_out1;

  out1162 <= Logical_Operator_out9866_out1;

  out1163 <= Logical_Operator_out9867_out1;

  out1164 <= Logical_Operator_out9868_out1;

  out1165 <= Logical_Operator_out9869_out1;

  out1166 <= Logical_Operator_out9870_out1;

  out1167 <= Logical_Operator_out9871_out1;

  out1168 <= Logical_Operator_out9872_out1;

  out1169 <= Logical_Operator_out9873_out1;

  out1170 <= Logical_Operator_out9874_out1;

  out1171 <= Logical_Operator_out9875_out1;

  out1172 <= Logical_Operator_out9876_out1;

  out1173 <= Logical_Operator_out9877_out1;

  out1174 <= Logical_Operator_out9878_out1;

  out1175 <= Logical_Operator_out9879_out1;

  out1176 <= Logical_Operator_out9880_out1;

  out1177 <= Logical_Operator_out9881_out1;

  out1178 <= Logical_Operator_out9882_out1;

  out1179 <= Logical_Operator_out9883_out1;

  out1180 <= Logical_Operator_out9884_out1;

  out1181 <= Logical_Operator_out9885_out1;

  out1182 <= Logical_Operator_out9886_out1;

  out1183 <= Logical_Operator_out9887_out1;

  out1184 <= Logical_Operator_out9888_out1;

  out1185 <= Logical_Operator_out9889_out1;

  out1186 <= Logical_Operator_out9890_out1;

  out1187 <= Logical_Operator_out9891_out1;

  out1188 <= Logical_Operator_out9892_out1;

  out1189 <= Logical_Operator_out9893_out1;

  out1190 <= Logical_Operator_out9894_out1;

  out1191 <= Logical_Operator_out9895_out1;

  out1192 <= Logical_Operator_out9896_out1;

  out1193 <= Logical_Operator_out9897_out1;

  out1194 <= Logical_Operator_out9898_out1;

  out1195 <= Logical_Operator_out9899_out1;

  out1196 <= Logical_Operator_out9900_out1;

  out1197 <= Logical_Operator_out9901_out1;

  out1198 <= Logical_Operator_out9902_out1;

  out1199 <= Logical_Operator_out9903_out1;

  out1200 <= Logical_Operator_out9904_out1;

  out1201 <= Logical_Operator_out9905_out1;

  out1202 <= Logical_Operator_out9906_out1;

  out1203 <= Logical_Operator_out9907_out1;

  out1204 <= Logical_Operator_out9908_out1;

  out1205 <= Logical_Operator_out9909_out1;

  out1206 <= Logical_Operator_out9910_out1;

  out1207 <= Logical_Operator_out9911_out1;

  out1208 <= Logical_Operator_out9912_out1;

  out1209 <= Logical_Operator_out9913_out1;

  out1210 <= Logical_Operator_out9914_out1;

  out1211 <= Logical_Operator_out9915_out1;

  out1212 <= Logical_Operator_out9916_out1;

  out1213 <= Logical_Operator_out9917_out1;

  out1214 <= Logical_Operator_out9918_out1;

  out1215 <= Logical_Operator_out9919_out1;

  out1216 <= Logical_Operator_out9920_out1;

  out1217 <= Logical_Operator_out9921_out1;

  out1218 <= Logical_Operator_out9922_out1;

  out1219 <= Logical_Operator_out9923_out1;

  out1220 <= Logical_Operator_out9924_out1;

  out1221 <= Logical_Operator_out9925_out1;

  out1222 <= Logical_Operator_out9926_out1;

  out1223 <= Logical_Operator_out9927_out1;

  out1224 <= Logical_Operator_out9928_out1;

  out1225 <= Logical_Operator_out9929_out1;

  out1226 <= Logical_Operator_out9930_out1;

  out1227 <= Logical_Operator_out9931_out1;

  out1228 <= Logical_Operator_out9932_out1;

  out1229 <= Logical_Operator_out9933_out1;

  out1230 <= Logical_Operator_out9934_out1;

  out1231 <= Logical_Operator_out9935_out1;

  out1232 <= Logical_Operator_out9936_out1;

  out1233 <= Logical_Operator_out9937_out1;

  out1234 <= Logical_Operator_out9938_out1;

  out1235 <= Logical_Operator_out9939_out1;

  out1236 <= Logical_Operator_out9940_out1;

  out1237 <= Logical_Operator_out9941_out1;

  out1238 <= Logical_Operator_out9942_out1;

  out1239 <= Logical_Operator_out9943_out1;

  out1240 <= Logical_Operator_out9944_out1;

  out1241 <= Logical_Operator_out9945_out1;

  out1242 <= Logical_Operator_out9946_out1;

  out1243 <= Logical_Operator_out9947_out1;

  out1244 <= Logical_Operator_out9948_out1;

  out1245 <= Logical_Operator_out9949_out1;

  out1246 <= Logical_Operator_out9950_out1;

  out1247 <= Logical_Operator_out9951_out1;

  out1248 <= Logical_Operator_out9952_out1;

  out1249 <= Logical_Operator_out9953_out1;

  out1250 <= Logical_Operator_out9954_out1;

  out1251 <= Logical_Operator_out9955_out1;

  out1252 <= Logical_Operator_out9956_out1;

  out1253 <= Logical_Operator_out9957_out1;

  out1254 <= Logical_Operator_out9958_out1;

  out1255 <= Logical_Operator_out9959_out1;

  out1256 <= Logical_Operator_out9960_out1;

  out1257 <= Logical_Operator_out9961_out1;

  out1258 <= Logical_Operator_out9962_out1;

  out1259 <= Logical_Operator_out9963_out1;

  out1260 <= Logical_Operator_out9964_out1;

  out1261 <= Logical_Operator_out9965_out1;

  out1262 <= Logical_Operator_out9966_out1;

  out1263 <= Logical_Operator_out9967_out1;

  out1264 <= Logical_Operator_out9968_out1;

  out1265 <= Logical_Operator_out9969_out1;

  out1266 <= Logical_Operator_out9970_out1;

  out1267 <= Logical_Operator_out9971_out1;

  out1268 <= Logical_Operator_out9972_out1;

  out1269 <= Logical_Operator_out9973_out1;

  out1270 <= Logical_Operator_out9974_out1;

  out1271 <= Logical_Operator_out9975_out1;

  out1272 <= Logical_Operator_out9976_out1;

  out1273 <= Logical_Operator_out9977_out1;

  out1274 <= Logical_Operator_out9978_out1;

  out1275 <= Logical_Operator_out9979_out1;

  out1276 <= Logical_Operator_out9980_out1;

  out1277 <= Logical_Operator_out9981_out1;

  out1278 <= Logical_Operator_out9982_out1;

  out1279 <= Logical_Operator_out9983_out1;

  out1280 <= Logical_Operator_out9984_out1;

  out1281 <= Logical_Operator_out9985_out1;

  out1282 <= Logical_Operator_out9986_out1;

  out1283 <= Logical_Operator_out9987_out1;

  out1284 <= Logical_Operator_out9988_out1;

  out1285 <= Logical_Operator_out9989_out1;

  out1286 <= Logical_Operator_out9990_out1;

  out1287 <= Logical_Operator_out9991_out1;

  out1288 <= Logical_Operator_out9992_out1;

  out1289 <= Logical_Operator_out9993_out1;

  out1290 <= Logical_Operator_out9994_out1;

  out1291 <= Logical_Operator_out9995_out1;

  out1292 <= Logical_Operator_out9996_out1;

  out1293 <= Logical_Operator_out9997_out1;

  out1294 <= Logical_Operator_out9998_out1;

  out1295 <= Logical_Operator_out9999_out1;

  out1296 <= Logical_Operator_out10000_out1;

  out1297 <= Logical_Operator_out10001_out1;

  out1298 <= Logical_Operator_out10002_out1;

  out1299 <= Logical_Operator_out10003_out1;

  out1300 <= Logical_Operator_out10004_out1;

  out1301 <= Logical_Operator_out10005_out1;

  out1302 <= Logical_Operator_out10006_out1;

  out1303 <= Logical_Operator_out10007_out1;

  out1304 <= Logical_Operator_out10008_out1;

  out1305 <= Logical_Operator_out10009_out1;

  out1306 <= Logical_Operator_out10010_out1;

  out1307 <= Logical_Operator_out10011_out1;

  out1308 <= Logical_Operator_out10012_out1;

  out1309 <= Logical_Operator_out10013_out1;

  out1310 <= Logical_Operator_out10014_out1;

  out1311 <= Logical_Operator_out10015_out1;

  out1312 <= Logical_Operator_out10016_out1;

  out1313 <= Logical_Operator_out10017_out1;

  out1314 <= Logical_Operator_out10018_out1;

  out1315 <= Logical_Operator_out10019_out1;

  out1316 <= Logical_Operator_out10020_out1;

  out1317 <= Logical_Operator_out10021_out1;

  out1318 <= Logical_Operator_out10022_out1;

  out1319 <= Logical_Operator_out10023_out1;

  out1320 <= Logical_Operator_out10024_out1;

  out1321 <= Logical_Operator_out10025_out1;

  out1322 <= Logical_Operator_out10026_out1;

  out1323 <= Logical_Operator_out10027_out1;

  out1324 <= Logical_Operator_out10028_out1;

  out1325 <= Logical_Operator_out10029_out1;

  out1326 <= Logical_Operator_out10030_out1;

  out1327 <= Logical_Operator_out10031_out1;

  out1328 <= Logical_Operator_out10032_out1;

  out1329 <= Logical_Operator_out10033_out1;

  out1330 <= Logical_Operator_out10034_out1;

  out1331 <= Logical_Operator_out10035_out1;

  out1332 <= Logical_Operator_out10036_out1;

  out1333 <= Logical_Operator_out10037_out1;

  out1334 <= Logical_Operator_out10038_out1;

  out1335 <= Logical_Operator_out10039_out1;

  out1336 <= Logical_Operator_out10040_out1;

  out1337 <= Logical_Operator_out10041_out1;

  out1338 <= Logical_Operator_out10042_out1;

  out1339 <= Logical_Operator_out10043_out1;

  out1340 <= Logical_Operator_out10044_out1;

  out1341 <= Logical_Operator_out10045_out1;

  out1342 <= Logical_Operator_out10046_out1;

  out1343 <= Logical_Operator_out10047_out1;

  out1344 <= Logical_Operator_out10048_out1;

  out1345 <= Logical_Operator_out10049_out1;

  out1346 <= Logical_Operator_out10050_out1;

  out1347 <= Logical_Operator_out10051_out1;

  out1348 <= Logical_Operator_out10052_out1;

  out1349 <= Logical_Operator_out10053_out1;

  out1350 <= Logical_Operator_out10054_out1;

  out1351 <= Logical_Operator_out10055_out1;

  out1352 <= Logical_Operator_out10056_out1;

  out1353 <= Logical_Operator_out10057_out1;

  out1354 <= Logical_Operator_out10058_out1;

  out1355 <= Logical_Operator_out10059_out1;

  out1356 <= Logical_Operator_out10060_out1;

  out1357 <= Logical_Operator_out10061_out1;

  out1358 <= Logical_Operator_out10062_out1;

  out1359 <= Logical_Operator_out10063_out1;

  out1360 <= Logical_Operator_out10064_out1;

  out1361 <= Logical_Operator_out10065_out1;

  out1362 <= Logical_Operator_out10066_out1;

  out1363 <= Logical_Operator_out10067_out1;

  out1364 <= Logical_Operator_out10068_out1;

  out1365 <= Logical_Operator_out10069_out1;

  out1366 <= Logical_Operator_out10070_out1;

  out1367 <= Logical_Operator_out10071_out1;

  out1368 <= Logical_Operator_out10072_out1;

  out1369 <= Logical_Operator_out10073_out1;

  out1370 <= Logical_Operator_out10074_out1;

  out1371 <= Logical_Operator_out10075_out1;

  out1372 <= Logical_Operator_out10076_out1;

  out1373 <= Logical_Operator_out10077_out1;

  out1374 <= Logical_Operator_out10078_out1;

  out1375 <= Logical_Operator_out10079_out1;

  out1376 <= Logical_Operator_out10080_out1;

  out1377 <= Logical_Operator_out10081_out1;

  out1378 <= Logical_Operator_out10082_out1;

  out1379 <= Logical_Operator_out10083_out1;

  out1380 <= Logical_Operator_out10084_out1;

  out1381 <= Logical_Operator_out10085_out1;

  out1382 <= Logical_Operator_out10086_out1;

  out1383 <= Logical_Operator_out10087_out1;

  out1384 <= Logical_Operator_out10088_out1;

  out1385 <= Logical_Operator_out10089_out1;

  out1386 <= Logical_Operator_out10090_out1;

  out1387 <= Logical_Operator_out10091_out1;

  out1388 <= Logical_Operator_out10092_out1;

  out1389 <= Logical_Operator_out10093_out1;

  out1390 <= Logical_Operator_out10094_out1;

  out1391 <= Logical_Operator_out10095_out1;

  out1392 <= Logical_Operator_out10096_out1;

  out1393 <= Logical_Operator_out10097_out1;

  out1394 <= Logical_Operator_out10098_out1;

  out1395 <= Logical_Operator_out10099_out1;

  out1396 <= Logical_Operator_out10100_out1;

  out1397 <= Logical_Operator_out10101_out1;

  out1398 <= Logical_Operator_out10102_out1;

  out1399 <= Logical_Operator_out10103_out1;

  out1400 <= Logical_Operator_out10104_out1;

  out1401 <= Logical_Operator_out10105_out1;

  out1402 <= Logical_Operator_out10106_out1;

  out1403 <= Logical_Operator_out10107_out1;

  out1404 <= Logical_Operator_out10108_out1;

  out1405 <= Logical_Operator_out10109_out1;

  out1406 <= Logical_Operator_out10110_out1;

  out1407 <= Logical_Operator_out10111_out1;

  out1408 <= Logical_Operator_out10112_out1;

  out1409 <= Logical_Operator_out10113_out1;

  out1410 <= Logical_Operator_out10114_out1;

  out1411 <= Logical_Operator_out10115_out1;

  out1412 <= Logical_Operator_out10116_out1;

  out1413 <= Logical_Operator_out10117_out1;

  out1414 <= Logical_Operator_out10118_out1;

  out1415 <= Logical_Operator_out10119_out1;

  out1416 <= Logical_Operator_out10120_out1;

  out1417 <= Logical_Operator_out10121_out1;

  out1418 <= Logical_Operator_out10122_out1;

  out1419 <= Logical_Operator_out10123_out1;

  out1420 <= Logical_Operator_out10124_out1;

  out1421 <= Logical_Operator_out10125_out1;

  out1422 <= Logical_Operator_out10126_out1;

  out1423 <= Logical_Operator_out10127_out1;

  out1424 <= Logical_Operator_out10128_out1;

  out1425 <= Logical_Operator_out10129_out1;

  out1426 <= Logical_Operator_out10130_out1;

  out1427 <= Logical_Operator_out10131_out1;

  out1428 <= Logical_Operator_out10132_out1;

  out1429 <= Logical_Operator_out10133_out1;

  out1430 <= Logical_Operator_out10134_out1;

  out1431 <= Logical_Operator_out10135_out1;

  out1432 <= Logical_Operator_out10136_out1;

  out1433 <= Logical_Operator_out10137_out1;

  out1434 <= Logical_Operator_out10138_out1;

  out1435 <= Logical_Operator_out10139_out1;

  out1436 <= Logical_Operator_out10140_out1;

  out1437 <= Logical_Operator_out10141_out1;

  out1438 <= Logical_Operator_out10142_out1;

  out1439 <= Logical_Operator_out10143_out1;

  out1440 <= Logical_Operator_out10144_out1;

  out1441 <= Logical_Operator_out10145_out1;

  out1442 <= Logical_Operator_out10146_out1;

  out1443 <= Logical_Operator_out10147_out1;

  out1444 <= Logical_Operator_out10148_out1;

  out1445 <= Logical_Operator_out10149_out1;

  out1446 <= Logical_Operator_out10150_out1;

  out1447 <= Logical_Operator_out10151_out1;

  out1448 <= Logical_Operator_out10152_out1;

  out1449 <= Logical_Operator_out10153_out1;

  out1450 <= Logical_Operator_out10154_out1;

  out1451 <= Logical_Operator_out10155_out1;

  out1452 <= Logical_Operator_out10156_out1;

  out1453 <= Logical_Operator_out10157_out1;

  out1454 <= Logical_Operator_out10158_out1;

  out1455 <= Logical_Operator_out10159_out1;

  out1456 <= Logical_Operator_out10160_out1;

  out1457 <= Logical_Operator_out10161_out1;

  out1458 <= Logical_Operator_out10162_out1;

  out1459 <= Logical_Operator_out10163_out1;

  out1460 <= Logical_Operator_out10164_out1;

  out1461 <= Logical_Operator_out10165_out1;

  out1462 <= Logical_Operator_out10166_out1;

  out1463 <= Logical_Operator_out10167_out1;

  out1464 <= Logical_Operator_out10168_out1;

  out1465 <= Logical_Operator_out10169_out1;

  out1466 <= Logical_Operator_out10170_out1;

  out1467 <= Logical_Operator_out10171_out1;

  out1468 <= Logical_Operator_out10172_out1;

  out1469 <= Logical_Operator_out10173_out1;

  out1470 <= Logical_Operator_out10174_out1;

  out1471 <= Logical_Operator_out10175_out1;

  out1472 <= Logical_Operator_out10176_out1;

  out1473 <= Logical_Operator_out10177_out1;

  out1474 <= Logical_Operator_out10178_out1;

  out1475 <= Logical_Operator_out10179_out1;

  out1476 <= Logical_Operator_out10180_out1;

  out1477 <= Logical_Operator_out10181_out1;

  out1478 <= Logical_Operator_out10182_out1;

  out1479 <= Logical_Operator_out10183_out1;

  out1480 <= Logical_Operator_out10184_out1;

  out1481 <= Logical_Operator_out10185_out1;

  out1482 <= Logical_Operator_out10186_out1;

  out1483 <= Logical_Operator_out10187_out1;

  out1484 <= Logical_Operator_out10188_out1;

  out1485 <= Logical_Operator_out10189_out1;

  out1486 <= Logical_Operator_out10190_out1;

  out1487 <= Logical_Operator_out10191_out1;

  out1488 <= Logical_Operator_out10192_out1;

  out1489 <= Logical_Operator_out10193_out1;

  out1490 <= Logical_Operator_out10194_out1;

  out1491 <= Logical_Operator_out10195_out1;

  out1492 <= Logical_Operator_out10196_out1;

  out1493 <= Logical_Operator_out10197_out1;

  out1494 <= Logical_Operator_out10198_out1;

  out1495 <= Logical_Operator_out10199_out1;

  out1496 <= Logical_Operator_out10200_out1;

  out1497 <= Logical_Operator_out10201_out1;

  out1498 <= Logical_Operator_out10202_out1;

  out1499 <= Logical_Operator_out10203_out1;

  out1500 <= Logical_Operator_out10204_out1;

  out1501 <= Logical_Operator_out10205_out1;

  out1502 <= Logical_Operator_out10206_out1;

  out1503 <= Logical_Operator_out10207_out1;

  out1504 <= Logical_Operator_out10208_out1;

  out1505 <= Logical_Operator_out10209_out1;

  out1506 <= Logical_Operator_out10210_out1;

  out1507 <= Logical_Operator_out10211_out1;

  out1508 <= Logical_Operator_out10212_out1;

  out1509 <= Logical_Operator_out10213_out1;

  out1510 <= Logical_Operator_out10214_out1;

  out1511 <= Logical_Operator_out10215_out1;

  out1512 <= Logical_Operator_out10216_out1;

  out1513 <= Logical_Operator_out10217_out1;

  out1514 <= Logical_Operator_out10218_out1;

  out1515 <= Logical_Operator_out10219_out1;

  out1516 <= Logical_Operator_out10220_out1;

  out1517 <= Logical_Operator_out10221_out1;

  out1518 <= Logical_Operator_out10222_out1;

  out1519 <= Logical_Operator_out10223_out1;

  out1520 <= Logical_Operator_out10224_out1;

  out1521 <= Logical_Operator_out10225_out1;

  out1522 <= Logical_Operator_out10226_out1;

  out1523 <= Logical_Operator_out10227_out1;

  out1524 <= Logical_Operator_out10228_out1;

  out1525 <= Logical_Operator_out10229_out1;

  out1526 <= Logical_Operator_out10230_out1;

  out1527 <= Logical_Operator_out10231_out1;

  out1528 <= Logical_Operator_out10232_out1;

  out1529 <= Logical_Operator_out10233_out1;

  out1530 <= Logical_Operator_out10234_out1;

  out1531 <= Logical_Operator_out10235_out1;

  out1532 <= Logical_Operator_out10236_out1;

  out1533 <= Logical_Operator_out10237_out1;

  out1534 <= Logical_Operator_out10238_out1;

  out1535 <= Logical_Operator_out10239_out1;

  out1536 <= Logical_Operator_out10240_out1;

  out1537 <= Logical_Operator_out8961_out1;

  out1538 <= Logical_Operator_out8962_out1;

  out1539 <= Logical_Operator_out8963_out1;

  out1540 <= Logical_Operator_out8964_out1;

  out1541 <= Logical_Operator_out8965_out1;

  out1542 <= Logical_Operator_out8966_out1;

  out1543 <= Logical_Operator_out8967_out1;

  out1544 <= Logical_Operator_out8968_out1;

  out1545 <= Logical_Operator_out8969_out1;

  out1546 <= Logical_Operator_out8970_out1;

  out1547 <= Logical_Operator_out8971_out1;

  out1548 <= Logical_Operator_out8972_out1;

  out1549 <= Logical_Operator_out8973_out1;

  out1550 <= Logical_Operator_out8974_out1;

  out1551 <= Logical_Operator_out8975_out1;

  out1552 <= Logical_Operator_out8976_out1;

  out1553 <= Logical_Operator_out8977_out1;

  out1554 <= Logical_Operator_out8978_out1;

  out1555 <= Logical_Operator_out8979_out1;

  out1556 <= Logical_Operator_out8980_out1;

  out1557 <= Logical_Operator_out8981_out1;

  out1558 <= Logical_Operator_out8982_out1;

  out1559 <= Logical_Operator_out8983_out1;

  out1560 <= Logical_Operator_out8984_out1;

  out1561 <= Logical_Operator_out8985_out1;

  out1562 <= Logical_Operator_out8986_out1;

  out1563 <= Logical_Operator_out8987_out1;

  out1564 <= Logical_Operator_out8988_out1;

  out1565 <= Logical_Operator_out8989_out1;

  out1566 <= Logical_Operator_out8990_out1;

  out1567 <= Logical_Operator_out8991_out1;

  out1568 <= Logical_Operator_out8992_out1;

  out1569 <= Logical_Operator_out8993_out1;

  out1570 <= Logical_Operator_out8994_out1;

  out1571 <= Logical_Operator_out8995_out1;

  out1572 <= Logical_Operator_out8996_out1;

  out1573 <= Logical_Operator_out8997_out1;

  out1574 <= Logical_Operator_out8998_out1;

  out1575 <= Logical_Operator_out8999_out1;

  out1576 <= Logical_Operator_out9000_out1;

  out1577 <= Logical_Operator_out9001_out1;

  out1578 <= Logical_Operator_out9002_out1;

  out1579 <= Logical_Operator_out9003_out1;

  out1580 <= Logical_Operator_out9004_out1;

  out1581 <= Logical_Operator_out9005_out1;

  out1582 <= Logical_Operator_out9006_out1;

  out1583 <= Logical_Operator_out9007_out1;

  out1584 <= Logical_Operator_out9008_out1;

  out1585 <= Logical_Operator_out9009_out1;

  out1586 <= Logical_Operator_out9010_out1;

  out1587 <= Logical_Operator_out9011_out1;

  out1588 <= Logical_Operator_out9012_out1;

  out1589 <= Logical_Operator_out9013_out1;

  out1590 <= Logical_Operator_out9014_out1;

  out1591 <= Logical_Operator_out9015_out1;

  out1592 <= Logical_Operator_out9016_out1;

  out1593 <= Logical_Operator_out9017_out1;

  out1594 <= Logical_Operator_out9018_out1;

  out1595 <= Logical_Operator_out9019_out1;

  out1596 <= Logical_Operator_out9020_out1;

  out1597 <= Logical_Operator_out9021_out1;

  out1598 <= Logical_Operator_out9022_out1;

  out1599 <= Logical_Operator_out9023_out1;

  out1600 <= Logical_Operator_out9024_out1;

  out1601 <= Logical_Operator_out9025_out1;

  out1602 <= Logical_Operator_out9026_out1;

  out1603 <= Logical_Operator_out9027_out1;

  out1604 <= Logical_Operator_out9028_out1;

  out1605 <= Logical_Operator_out9029_out1;

  out1606 <= Logical_Operator_out9030_out1;

  out1607 <= Logical_Operator_out9031_out1;

  out1608 <= Logical_Operator_out9032_out1;

  out1609 <= Logical_Operator_out9033_out1;

  out1610 <= Logical_Operator_out9034_out1;

  out1611 <= Logical_Operator_out9035_out1;

  out1612 <= Logical_Operator_out9036_out1;

  out1613 <= Logical_Operator_out9037_out1;

  out1614 <= Logical_Operator_out9038_out1;

  out1615 <= Logical_Operator_out9039_out1;

  out1616 <= Logical_Operator_out9040_out1;

  out1617 <= Logical_Operator_out9041_out1;

  out1618 <= Logical_Operator_out9042_out1;

  out1619 <= Logical_Operator_out9043_out1;

  out1620 <= Logical_Operator_out9044_out1;

  out1621 <= Logical_Operator_out9045_out1;

  out1622 <= Logical_Operator_out9046_out1;

  out1623 <= Logical_Operator_out9047_out1;

  out1624 <= Logical_Operator_out9048_out1;

  out1625 <= Logical_Operator_out9049_out1;

  out1626 <= Logical_Operator_out9050_out1;

  out1627 <= Logical_Operator_out9051_out1;

  out1628 <= Logical_Operator_out9052_out1;

  out1629 <= Logical_Operator_out9053_out1;

  out1630 <= Logical_Operator_out9054_out1;

  out1631 <= Logical_Operator_out9055_out1;

  out1632 <= Logical_Operator_out9056_out1;

  out1633 <= Logical_Operator_out9057_out1;

  out1634 <= Logical_Operator_out9058_out1;

  out1635 <= Logical_Operator_out9059_out1;

  out1636 <= Logical_Operator_out9060_out1;

  out1637 <= Logical_Operator_out9061_out1;

  out1638 <= Logical_Operator_out9062_out1;

  out1639 <= Logical_Operator_out9063_out1;

  out1640 <= Logical_Operator_out9064_out1;

  out1641 <= Logical_Operator_out9065_out1;

  out1642 <= Logical_Operator_out9066_out1;

  out1643 <= Logical_Operator_out9067_out1;

  out1644 <= Logical_Operator_out9068_out1;

  out1645 <= Logical_Operator_out9069_out1;

  out1646 <= Logical_Operator_out9070_out1;

  out1647 <= Logical_Operator_out9071_out1;

  out1648 <= Logical_Operator_out9072_out1;

  out1649 <= Logical_Operator_out9073_out1;

  out1650 <= Logical_Operator_out9074_out1;

  out1651 <= Logical_Operator_out9075_out1;

  out1652 <= Logical_Operator_out9076_out1;

  out1653 <= Logical_Operator_out9077_out1;

  out1654 <= Logical_Operator_out9078_out1;

  out1655 <= Logical_Operator_out9079_out1;

  out1656 <= Logical_Operator_out9080_out1;

  out1657 <= Logical_Operator_out9081_out1;

  out1658 <= Logical_Operator_out9082_out1;

  out1659 <= Logical_Operator_out9083_out1;

  out1660 <= Logical_Operator_out9084_out1;

  out1661 <= Logical_Operator_out9085_out1;

  out1662 <= Logical_Operator_out9086_out1;

  out1663 <= Logical_Operator_out9087_out1;

  out1664 <= Logical_Operator_out9088_out1;

  out1665 <= Logical_Operator_out9089_out1;

  out1666 <= Logical_Operator_out9090_out1;

  out1667 <= Logical_Operator_out9091_out1;

  out1668 <= Logical_Operator_out9092_out1;

  out1669 <= Logical_Operator_out9093_out1;

  out1670 <= Logical_Operator_out9094_out1;

  out1671 <= Logical_Operator_out9095_out1;

  out1672 <= Logical_Operator_out9096_out1;

  out1673 <= Logical_Operator_out9097_out1;

  out1674 <= Logical_Operator_out9098_out1;

  out1675 <= Logical_Operator_out9099_out1;

  out1676 <= Logical_Operator_out9100_out1;

  out1677 <= Logical_Operator_out9101_out1;

  out1678 <= Logical_Operator_out9102_out1;

  out1679 <= Logical_Operator_out9103_out1;

  out1680 <= Logical_Operator_out9104_out1;

  out1681 <= Logical_Operator_out9105_out1;

  out1682 <= Logical_Operator_out9106_out1;

  out1683 <= Logical_Operator_out9107_out1;

  out1684 <= Logical_Operator_out9108_out1;

  out1685 <= Logical_Operator_out9109_out1;

  out1686 <= Logical_Operator_out9110_out1;

  out1687 <= Logical_Operator_out9111_out1;

  out1688 <= Logical_Operator_out9112_out1;

  out1689 <= Logical_Operator_out9113_out1;

  out1690 <= Logical_Operator_out9114_out1;

  out1691 <= Logical_Operator_out9115_out1;

  out1692 <= Logical_Operator_out9116_out1;

  out1693 <= Logical_Operator_out9117_out1;

  out1694 <= Logical_Operator_out9118_out1;

  out1695 <= Logical_Operator_out9119_out1;

  out1696 <= Logical_Operator_out9120_out1;

  out1697 <= Logical_Operator_out9121_out1;

  out1698 <= Logical_Operator_out9122_out1;

  out1699 <= Logical_Operator_out9123_out1;

  out1700 <= Logical_Operator_out9124_out1;

  out1701 <= Logical_Operator_out9125_out1;

  out1702 <= Logical_Operator_out9126_out1;

  out1703 <= Logical_Operator_out9127_out1;

  out1704 <= Logical_Operator_out9128_out1;

  out1705 <= Logical_Operator_out9129_out1;

  out1706 <= Logical_Operator_out9130_out1;

  out1707 <= Logical_Operator_out9131_out1;

  out1708 <= Logical_Operator_out9132_out1;

  out1709 <= Logical_Operator_out9133_out1;

  out1710 <= Logical_Operator_out9134_out1;

  out1711 <= Logical_Operator_out9135_out1;

  out1712 <= Logical_Operator_out9136_out1;

  out1713 <= Logical_Operator_out9137_out1;

  out1714 <= Logical_Operator_out9138_out1;

  out1715 <= Logical_Operator_out9139_out1;

  out1716 <= Logical_Operator_out9140_out1;

  out1717 <= Logical_Operator_out9141_out1;

  out1718 <= Logical_Operator_out9142_out1;

  out1719 <= Logical_Operator_out9143_out1;

  out1720 <= Logical_Operator_out9144_out1;

  out1721 <= Logical_Operator_out9145_out1;

  out1722 <= Logical_Operator_out9146_out1;

  out1723 <= Logical_Operator_out9147_out1;

  out1724 <= Logical_Operator_out9148_out1;

  out1725 <= Logical_Operator_out9149_out1;

  out1726 <= Logical_Operator_out9150_out1;

  out1727 <= Logical_Operator_out9151_out1;

  out1728 <= Logical_Operator_out9152_out1;

  out1729 <= Logical_Operator_out9153_out1;

  out1730 <= Logical_Operator_out9154_out1;

  out1731 <= Logical_Operator_out9155_out1;

  out1732 <= Logical_Operator_out9156_out1;

  out1733 <= Logical_Operator_out9157_out1;

  out1734 <= Logical_Operator_out9158_out1;

  out1735 <= Logical_Operator_out9159_out1;

  out1736 <= Logical_Operator_out9160_out1;

  out1737 <= Logical_Operator_out9161_out1;

  out1738 <= Logical_Operator_out9162_out1;

  out1739 <= Logical_Operator_out9163_out1;

  out1740 <= Logical_Operator_out9164_out1;

  out1741 <= Logical_Operator_out9165_out1;

  out1742 <= Logical_Operator_out9166_out1;

  out1743 <= Logical_Operator_out9167_out1;

  out1744 <= Logical_Operator_out9168_out1;

  out1745 <= Logical_Operator_out9169_out1;

  out1746 <= Logical_Operator_out9170_out1;

  out1747 <= Logical_Operator_out9171_out1;

  out1748 <= Logical_Operator_out9172_out1;

  out1749 <= Logical_Operator_out9173_out1;

  out1750 <= Logical_Operator_out9174_out1;

  out1751 <= Logical_Operator_out9175_out1;

  out1752 <= Logical_Operator_out9176_out1;

  out1753 <= Logical_Operator_out9177_out1;

  out1754 <= Logical_Operator_out9178_out1;

  out1755 <= Logical_Operator_out9179_out1;

  out1756 <= Logical_Operator_out9180_out1;

  out1757 <= Logical_Operator_out9181_out1;

  out1758 <= Logical_Operator_out9182_out1;

  out1759 <= Logical_Operator_out9183_out1;

  out1760 <= Logical_Operator_out9184_out1;

  out1761 <= Logical_Operator_out9185_out1;

  out1762 <= Logical_Operator_out9186_out1;

  out1763 <= Logical_Operator_out9187_out1;

  out1764 <= Logical_Operator_out9188_out1;

  out1765 <= Logical_Operator_out9189_out1;

  out1766 <= Logical_Operator_out9190_out1;

  out1767 <= Logical_Operator_out9191_out1;

  out1768 <= Logical_Operator_out9192_out1;

  out1769 <= Logical_Operator_out9193_out1;

  out1770 <= Logical_Operator_out9194_out1;

  out1771 <= Logical_Operator_out9195_out1;

  out1772 <= Logical_Operator_out9196_out1;

  out1773 <= Logical_Operator_out9197_out1;

  out1774 <= Logical_Operator_out9198_out1;

  out1775 <= Logical_Operator_out9199_out1;

  out1776 <= Logical_Operator_out9200_out1;

  out1777 <= Logical_Operator_out9201_out1;

  out1778 <= Logical_Operator_out9202_out1;

  out1779 <= Logical_Operator_out9203_out1;

  out1780 <= Logical_Operator_out9204_out1;

  out1781 <= Logical_Operator_out9205_out1;

  out1782 <= Logical_Operator_out9206_out1;

  out1783 <= Logical_Operator_out9207_out1;

  out1784 <= Logical_Operator_out9208_out1;

  out1785 <= Logical_Operator_out9209_out1;

  out1786 <= Logical_Operator_out9210_out1;

  out1787 <= Logical_Operator_out9211_out1;

  out1788 <= Logical_Operator_out9212_out1;

  out1789 <= Logical_Operator_out9213_out1;

  out1790 <= Logical_Operator_out9214_out1;

  out1791 <= Logical_Operator_out9215_out1;

  out1792 <= Logical_Operator_out9216_out1;

  out1793 <= Logical_Operator_out8065_out1;

  out1794 <= Logical_Operator_out8066_out1;

  out1795 <= Logical_Operator_out8067_out1;

  out1796 <= Logical_Operator_out8068_out1;

  out1797 <= Logical_Operator_out8069_out1;

  out1798 <= Logical_Operator_out8070_out1;

  out1799 <= Logical_Operator_out8071_out1;

  out1800 <= Logical_Operator_out8072_out1;

  out1801 <= Logical_Operator_out8073_out1;

  out1802 <= Logical_Operator_out8074_out1;

  out1803 <= Logical_Operator_out8075_out1;

  out1804 <= Logical_Operator_out8076_out1;

  out1805 <= Logical_Operator_out8077_out1;

  out1806 <= Logical_Operator_out8078_out1;

  out1807 <= Logical_Operator_out8079_out1;

  out1808 <= Logical_Operator_out8080_out1;

  out1809 <= Logical_Operator_out8081_out1;

  out1810 <= Logical_Operator_out8082_out1;

  out1811 <= Logical_Operator_out8083_out1;

  out1812 <= Logical_Operator_out8084_out1;

  out1813 <= Logical_Operator_out8085_out1;

  out1814 <= Logical_Operator_out8086_out1;

  out1815 <= Logical_Operator_out8087_out1;

  out1816 <= Logical_Operator_out8088_out1;

  out1817 <= Logical_Operator_out8089_out1;

  out1818 <= Logical_Operator_out8090_out1;

  out1819 <= Logical_Operator_out8091_out1;

  out1820 <= Logical_Operator_out8092_out1;

  out1821 <= Logical_Operator_out8093_out1;

  out1822 <= Logical_Operator_out8094_out1;

  out1823 <= Logical_Operator_out8095_out1;

  out1824 <= Logical_Operator_out8096_out1;

  out1825 <= Logical_Operator_out8097_out1;

  out1826 <= Logical_Operator_out8098_out1;

  out1827 <= Logical_Operator_out8099_out1;

  out1828 <= Logical_Operator_out8100_out1;

  out1829 <= Logical_Operator_out8101_out1;

  out1830 <= Logical_Operator_out8102_out1;

  out1831 <= Logical_Operator_out8103_out1;

  out1832 <= Logical_Operator_out8104_out1;

  out1833 <= Logical_Operator_out8105_out1;

  out1834 <= Logical_Operator_out8106_out1;

  out1835 <= Logical_Operator_out8107_out1;

  out1836 <= Logical_Operator_out8108_out1;

  out1837 <= Logical_Operator_out8109_out1;

  out1838 <= Logical_Operator_out8110_out1;

  out1839 <= Logical_Operator_out8111_out1;

  out1840 <= Logical_Operator_out8112_out1;

  out1841 <= Logical_Operator_out8113_out1;

  out1842 <= Logical_Operator_out8114_out1;

  out1843 <= Logical_Operator_out8115_out1;

  out1844 <= Logical_Operator_out8116_out1;

  out1845 <= Logical_Operator_out8117_out1;

  out1846 <= Logical_Operator_out8118_out1;

  out1847 <= Logical_Operator_out8119_out1;

  out1848 <= Logical_Operator_out8120_out1;

  out1849 <= Logical_Operator_out8121_out1;

  out1850 <= Logical_Operator_out8122_out1;

  out1851 <= Logical_Operator_out8123_out1;

  out1852 <= Logical_Operator_out8124_out1;

  out1853 <= Logical_Operator_out8125_out1;

  out1854 <= Logical_Operator_out8126_out1;

  out1855 <= Logical_Operator_out8127_out1;

  out1856 <= Logical_Operator_out8128_out1;

  out1857 <= Logical_Operator_out8129_out1;

  out1858 <= Logical_Operator_out8130_out1;

  out1859 <= Logical_Operator_out8131_out1;

  out1860 <= Logical_Operator_out8132_out1;

  out1861 <= Logical_Operator_out8133_out1;

  out1862 <= Logical_Operator_out8134_out1;

  out1863 <= Logical_Operator_out8135_out1;

  out1864 <= Logical_Operator_out8136_out1;

  out1865 <= Logical_Operator_out8137_out1;

  out1866 <= Logical_Operator_out8138_out1;

  out1867 <= Logical_Operator_out8139_out1;

  out1868 <= Logical_Operator_out8140_out1;

  out1869 <= Logical_Operator_out8141_out1;

  out1870 <= Logical_Operator_out8142_out1;

  out1871 <= Logical_Operator_out8143_out1;

  out1872 <= Logical_Operator_out8144_out1;

  out1873 <= Logical_Operator_out8145_out1;

  out1874 <= Logical_Operator_out8146_out1;

  out1875 <= Logical_Operator_out8147_out1;

  out1876 <= Logical_Operator_out8148_out1;

  out1877 <= Logical_Operator_out8149_out1;

  out1878 <= Logical_Operator_out8150_out1;

  out1879 <= Logical_Operator_out8151_out1;

  out1880 <= Logical_Operator_out8152_out1;

  out1881 <= Logical_Operator_out8153_out1;

  out1882 <= Logical_Operator_out8154_out1;

  out1883 <= Logical_Operator_out8155_out1;

  out1884 <= Logical_Operator_out8156_out1;

  out1885 <= Logical_Operator_out8157_out1;

  out1886 <= Logical_Operator_out8158_out1;

  out1887 <= Logical_Operator_out8159_out1;

  out1888 <= Logical_Operator_out8160_out1;

  out1889 <= Logical_Operator_out8161_out1;

  out1890 <= Logical_Operator_out8162_out1;

  out1891 <= Logical_Operator_out8163_out1;

  out1892 <= Logical_Operator_out8164_out1;

  out1893 <= Logical_Operator_out8165_out1;

  out1894 <= Logical_Operator_out8166_out1;

  out1895 <= Logical_Operator_out8167_out1;

  out1896 <= Logical_Operator_out8168_out1;

  out1897 <= Logical_Operator_out8169_out1;

  out1898 <= Logical_Operator_out8170_out1;

  out1899 <= Logical_Operator_out8171_out1;

  out1900 <= Logical_Operator_out8172_out1;

  out1901 <= Logical_Operator_out8173_out1;

  out1902 <= Logical_Operator_out8174_out1;

  out1903 <= Logical_Operator_out8175_out1;

  out1904 <= Logical_Operator_out8176_out1;

  out1905 <= Logical_Operator_out8177_out1;

  out1906 <= Logical_Operator_out8178_out1;

  out1907 <= Logical_Operator_out8179_out1;

  out1908 <= Logical_Operator_out8180_out1;

  out1909 <= Logical_Operator_out8181_out1;

  out1910 <= Logical_Operator_out8182_out1;

  out1911 <= Logical_Operator_out8183_out1;

  out1912 <= Logical_Operator_out8184_out1;

  out1913 <= Logical_Operator_out8185_out1;

  out1914 <= Logical_Operator_out8186_out1;

  out1915 <= Logical_Operator_out8187_out1;

  out1916 <= Logical_Operator_out8188_out1;

  out1917 <= Logical_Operator_out8189_out1;

  out1918 <= Logical_Operator_out8190_out1;

  out1919 <= Logical_Operator_out8191_out1;

  out1920 <= Logical_Operator_out8192_out1;

  out1921 <= Logical_Operator_out7105_out1;

  out1922 <= Logical_Operator_out7106_out1;

  out1923 <= Logical_Operator_out7107_out1;

  out1924 <= Logical_Operator_out7108_out1;

  out1925 <= Logical_Operator_out7109_out1;

  out1926 <= Logical_Operator_out7110_out1;

  out1927 <= Logical_Operator_out7111_out1;

  out1928 <= Logical_Operator_out7112_out1;

  out1929 <= Logical_Operator_out7113_out1;

  out1930 <= Logical_Operator_out7114_out1;

  out1931 <= Logical_Operator_out7115_out1;

  out1932 <= Logical_Operator_out7116_out1;

  out1933 <= Logical_Operator_out7117_out1;

  out1934 <= Logical_Operator_out7118_out1;

  out1935 <= Logical_Operator_out7119_out1;

  out1936 <= Logical_Operator_out7120_out1;

  out1937 <= Logical_Operator_out7121_out1;

  out1938 <= Logical_Operator_out7122_out1;

  out1939 <= Logical_Operator_out7123_out1;

  out1940 <= Logical_Operator_out7124_out1;

  out1941 <= Logical_Operator_out7125_out1;

  out1942 <= Logical_Operator_out7126_out1;

  out1943 <= Logical_Operator_out7127_out1;

  out1944 <= Logical_Operator_out7128_out1;

  out1945 <= Logical_Operator_out7129_out1;

  out1946 <= Logical_Operator_out7130_out1;

  out1947 <= Logical_Operator_out7131_out1;

  out1948 <= Logical_Operator_out7132_out1;

  out1949 <= Logical_Operator_out7133_out1;

  out1950 <= Logical_Operator_out7134_out1;

  out1951 <= Logical_Operator_out7135_out1;

  out1952 <= Logical_Operator_out7136_out1;

  out1953 <= Logical_Operator_out7137_out1;

  out1954 <= Logical_Operator_out7138_out1;

  out1955 <= Logical_Operator_out7139_out1;

  out1956 <= Logical_Operator_out7140_out1;

  out1957 <= Logical_Operator_out7141_out1;

  out1958 <= Logical_Operator_out7142_out1;

  out1959 <= Logical_Operator_out7143_out1;

  out1960 <= Logical_Operator_out7144_out1;

  out1961 <= Logical_Operator_out7145_out1;

  out1962 <= Logical_Operator_out7146_out1;

  out1963 <= Logical_Operator_out7147_out1;

  out1964 <= Logical_Operator_out7148_out1;

  out1965 <= Logical_Operator_out7149_out1;

  out1966 <= Logical_Operator_out7150_out1;

  out1967 <= Logical_Operator_out7151_out1;

  out1968 <= Logical_Operator_out7152_out1;

  out1969 <= Logical_Operator_out7153_out1;

  out1970 <= Logical_Operator_out7154_out1;

  out1971 <= Logical_Operator_out7155_out1;

  out1972 <= Logical_Operator_out7156_out1;

  out1973 <= Logical_Operator_out7157_out1;

  out1974 <= Logical_Operator_out7158_out1;

  out1975 <= Logical_Operator_out7159_out1;

  out1976 <= Logical_Operator_out7160_out1;

  out1977 <= Logical_Operator_out7161_out1;

  out1978 <= Logical_Operator_out7162_out1;

  out1979 <= Logical_Operator_out7163_out1;

  out1980 <= Logical_Operator_out7164_out1;

  out1981 <= Logical_Operator_out7165_out1;

  out1982 <= Logical_Operator_out7166_out1;

  out1983 <= Logical_Operator_out7167_out1;

  out1984 <= Logical_Operator_out7168_out1;

  out1985 <= Logical_Operator_out6113_out1;

  out1986 <= Logical_Operator_out6114_out1;

  out1987 <= Logical_Operator_out6115_out1;

  out1988 <= Logical_Operator_out6116_out1;

  out1989 <= Logical_Operator_out6117_out1;

  out1990 <= Logical_Operator_out6118_out1;

  out1991 <= Logical_Operator_out6119_out1;

  out1992 <= Logical_Operator_out6120_out1;

  out1993 <= Logical_Operator_out6121_out1;

  out1994 <= Logical_Operator_out6122_out1;

  out1995 <= Logical_Operator_out6123_out1;

  out1996 <= Logical_Operator_out6124_out1;

  out1997 <= Logical_Operator_out6125_out1;

  out1998 <= Logical_Operator_out6126_out1;

  out1999 <= Logical_Operator_out6127_out1;

  out2000 <= Logical_Operator_out6128_out1;

  out2001 <= Logical_Operator_out6129_out1;

  out2002 <= Logical_Operator_out6130_out1;

  out2003 <= Logical_Operator_out6131_out1;

  out2004 <= Logical_Operator_out6132_out1;

  out2005 <= Logical_Operator_out6133_out1;

  out2006 <= Logical_Operator_out6134_out1;

  out2007 <= Logical_Operator_out6135_out1;

  out2008 <= Logical_Operator_out6136_out1;

  out2009 <= Logical_Operator_out6137_out1;

  out2010 <= Logical_Operator_out6138_out1;

  out2011 <= Logical_Operator_out6139_out1;

  out2012 <= Logical_Operator_out6140_out1;

  out2013 <= Logical_Operator_out6141_out1;

  out2014 <= Logical_Operator_out6142_out1;

  out2015 <= Logical_Operator_out6143_out1;

  out2016 <= Logical_Operator_out6144_out1;

  out2017 <= Logical_Operator_out5105_out1;

  out2018 <= Logical_Operator_out5106_out1;

  out2019 <= Logical_Operator_out5107_out1;

  out2020 <= Logical_Operator_out5108_out1;

  out2021 <= Logical_Operator_out5109_out1;

  out2022 <= Logical_Operator_out5110_out1;

  out2023 <= Logical_Operator_out5111_out1;

  out2024 <= Logical_Operator_out5112_out1;

  out2025 <= Logical_Operator_out5113_out1;

  out2026 <= Logical_Operator_out5114_out1;

  out2027 <= Logical_Operator_out5115_out1;

  out2028 <= Logical_Operator_out5116_out1;

  out2029 <= Logical_Operator_out5117_out1;

  out2030 <= Logical_Operator_out5118_out1;

  out2031 <= Logical_Operator_out5119_out1;

  out2032 <= Logical_Operator_out5120_out1;

  out2033 <= Logical_Operator_out4089_out1;

  out2034 <= Logical_Operator_out4090_out1;

  out2035 <= Logical_Operator_out4091_out1;

  out2036 <= Logical_Operator_out4092_out1;

  out2037 <= Logical_Operator_out4093_out1;

  out2038 <= Logical_Operator_out4094_out1;

  out2039 <= Logical_Operator_out4095_out1;

  out2040 <= Logical_Operator_out4096_out1;

  out2041 <= Logical_Operator_out3069_out1;

  out2042 <= Logical_Operator_out3070_out1;

  out2043 <= Logical_Operator_out3071_out1;

  out2044 <= Logical_Operator_out3072_out1;

  out2045 <= Logical_Operator_out2047_out1;

  out2046 <= Logical_Operator_out2048_out1;

  out2047 <= Logical_Operator_out1024_out1;

  out2048 <= in2048;

END rtl;
